// Generated using findDep.cpp 
module query10_query45_1344n (v_1, v_2, v_3, v_4, v_5, v_6, v_7, v_8, v_9, v_10, v_11, v_12, v_13, v_14, v_15, v_16, v_17, v_18, v_20, v_21, v_22, v_23, v_24, v_25, v_26, v_27, v_28, v_29, v_30, v_31, v_32, v_33, v_34, v_35, v_36, v_37, v_38, v_39, v_40, v_41, v_42, v_43, v_44, v_45, v_46, v_47, v_48, v_49, v_50, v_51, v_52, v_53, v_54, v_55, v_56, v_57, v_58, v_59, v_60, v_61, v_62, v_63, v_64, v_65, v_66, v_67, v_68, v_69, v_70, v_71, v_72, v_73, v_74, v_75, v_76, v_77, v_78, v_79, v_80, v_81, v_82, v_83, v_84, v_85, v_86, v_87, v_88, v_89, v_90, v_91, v_92, v_93, v_94, v_95, v_96, v_97, v_98, v_99, v_100, v_101, v_102, v_103, v_104, v_105, v_106, v_107, v_108, v_109, v_110, v_111, v_112, v_113, v_114, v_115, v_116, v_117, v_118, v_119, v_120, v_121, v_122, v_123, v_124, v_125, v_126, v_127, v_128, v_129, v_130, v_131, v_132, v_133, v_134, v_135, v_136, v_137, v_138, v_142, v_143, v_144, v_145, v_146, v_147, v_148, v_149, v_150, v_151, v_155, v_159, v_160, v_161, v_162, v_163, v_164, v_165, v_166, v_167, v_168, v_169, v_170, v_171, v_172, v_179, v_180, v_181, v_182, v_183, v_184, v_19, v_139, v_140, v_141, v_152, v_153, v_154, v_156, v_157, v_158, v_173, v_174, v_175, v_176, v_177, v_178, v_185, v_186, v_187, v_188, v_189, v_190, v_191, v_192, v_193, v_194, v_195, v_196, v_197, v_198, v_199, v_200, v_201, v_202, v_203, v_204, v_205, v_206, v_207, v_208, v_209, v_210, v_211, v_212, v_213, v_214, v_215, v_216, v_217, v_218, v_219, v_220, v_221, v_222, v_223, v_224, v_225, v_226, v_227, v_228, v_229, v_230, v_231, v_232, v_233, v_234, v_235, v_236, v_237, v_238, v_239, v_240, v_241, v_242, v_243, v_244, v_245, v_246, v_247, v_248, v_249, v_250, v_251, v_252, v_253, v_254, v_255, v_256, v_257, v_258, v_259, v_260, v_261, v_262, v_263, v_264, v_265, v_266, v_267, v_268, v_269, v_270, v_271, v_272, v_273, v_274, v_275, v_276, v_277, v_278, v_279, v_280, v_281, v_282, v_283, v_284, v_285, v_286, v_287, v_288, v_289, v_290, v_291, v_292, v_293, v_294, v_295, v_296, v_297, v_298, v_299, v_300, v_301, v_302, v_303, v_304, v_305, v_306, v_307, v_308, v_309, v_310, v_311, v_312, v_313, v_314, v_315, v_316, v_317, v_318, v_319, v_320, v_321, v_322, v_323, v_324, v_325, v_326, v_327, v_328, v_329, v_330, v_331, v_332, v_333, v_334, v_335, v_336, v_337, v_338, v_339, v_340, v_341, v_342, v_343, v_344, v_345, v_346, v_347, v_348, v_349, v_350, v_351, v_352, v_353, v_354, v_355, v_356, v_357, v_358, v_359, v_360, v_361, v_362, v_363, v_364, v_365, v_366, v_367, v_368, v_369, v_370, v_371, v_372, v_373, v_374, v_375, v_376, v_377, v_378, v_379, v_380, v_381, v_382, v_383, v_384, v_385, v_386, v_387, v_388, v_389, v_390, v_391, v_392, v_393, v_394, v_395, v_396, v_397, v_398, v_399, v_400, v_401, v_402, v_403, v_404, v_405, v_406, v_407, v_408, v_409, v_410, v_411, v_412, v_413, v_414, v_415, v_416, v_417, v_418, v_419, v_420, v_421, v_422, v_423, v_424, v_425, v_426, v_427, v_428, v_429, v_430, v_431, v_432, v_433, v_434, v_435, v_436, v_437, v_438, v_439, v_440, v_441, v_442, v_443, v_444, v_445, v_446, v_447, v_448, v_449, v_450, v_451, v_452, v_453, v_454, v_455, v_456, v_457, v_458, v_459, v_460, v_461, v_462, v_463, v_464, v_465, v_466, v_467, v_468, v_469, v_470, v_471, v_472, v_473, v_474, v_475, v_476, v_477, v_478, v_479, v_480, v_481, v_482, v_483, v_484, v_485, v_486, v_487, v_488, v_489, v_490, v_491, v_492, v_493, v_494, v_495, v_496, v_497, v_498, v_499, v_500, v_501, v_502, v_503, v_504, v_505, v_506, v_507, v_508, v_509, v_510, v_511, v_512, v_513, v_514, v_515, v_516, v_517, v_518, v_519, v_520, v_521, v_522, v_523, v_524, v_525, v_526, v_527, v_528, v_529, v_530, v_531, v_532, v_533, v_534, v_535, v_536, v_537, v_538, v_539, v_540, v_541, v_542, v_543, v_544, v_545, v_546, v_547, v_548, v_549, v_550, v_551, v_552, v_553, v_554, v_555, v_556, v_557, v_558, v_559, v_560, v_561, v_562, v_563, v_564, v_565, v_566, v_567, v_568, v_569, v_570, v_571, v_572, v_573, v_574, v_575, v_576, v_577, v_578, v_579, v_580, v_581, v_582, v_583, v_584, v_585, v_586, v_587, v_588, v_589, v_590, v_591, v_592, v_593, v_594, v_595, v_596, v_597, v_598, v_599, v_600, v_601, v_602, v_603, v_604, v_605, v_606, v_607, v_608, v_609, v_610, v_611, v_612, v_613, v_614, v_615, v_616, v_617, v_618, v_619, v_620, v_621, v_622, v_623, v_624, v_625, v_626, v_627, v_628, v_629, v_630, v_631, v_632, v_633, v_634, v_635, v_636, v_637, v_638, v_639, v_640, v_641, v_642, v_643, v_644, v_645, v_646, v_647, v_648, v_649, v_650, v_651, v_652, v_653, v_654, v_655, v_656, v_657, v_658, v_659, v_660, v_661, v_662, v_663, v_664, v_665, v_666, v_667, v_668, v_669, v_670, v_671, v_672, v_673, v_674, v_675, v_676, v_677, v_678, v_679, v_680, v_681, v_682, v_683, v_684, v_685, v_686, v_687, v_688, v_689, v_690, v_691, v_692, v_693, v_694, v_695, v_696, v_697, v_698, v_699, v_700, v_701, v_702, v_703, v_704, v_705, v_706, v_707, v_708, v_709, v_710, v_711, v_712, v_713, v_714, v_715, v_716, v_717, v_718, v_719, v_720, v_721, v_722, v_723, v_724, v_725, v_726, v_727, v_728, v_729, v_730, v_731, v_732, v_733, v_734, v_735, v_736, v_737, v_738, v_739, v_740, v_741, v_742, v_743, v_744, v_745, v_746, v_747, v_748, v_749, v_750, v_751, v_752, v_753, v_754, v_755, v_756, v_757, v_758, v_759, v_760, v_761, v_762, v_763, v_764, v_765, v_766, v_767, v_768, v_769, v_770, v_771, v_772, v_773, v_774, v_775, v_776, v_777, v_778, v_779, v_780, v_781, v_782, v_783, v_784, v_785, v_786, v_787, v_788, v_789, v_790, v_791, v_792, v_793, v_794, v_795, v_796, v_797, v_798, v_799, v_800, v_801, v_802, v_803, v_804, v_805, v_806, v_807, v_808, v_809, v_810, v_811, v_812, v_813, v_814, v_815, v_816, v_817, v_818, v_819, v_820, v_821, v_822, v_823, v_824, v_825, v_826, v_827, v_828, v_829, v_830, v_831, v_832, v_833, v_834, v_835, v_836, v_837, v_838, v_839, v_840, v_841, v_842, v_843, v_844, v_845, v_846, v_847, v_848, v_849, v_850, v_851, v_852, v_853, v_854, v_855, v_856, v_857, v_858, v_859, v_860, v_861, v_862, v_863, v_864, v_865, v_866, v_867, v_868, v_869, v_870, v_871, v_872, v_873, v_874, v_875, v_876, v_877, v_878, v_879, v_880, v_881, v_882, v_883, v_884, v_885, v_886, v_887, v_888, v_889, v_890, v_891, v_892, v_893, v_894, v_895, v_896, v_897, v_898, v_899, v_900, v_901, v_902, v_903, v_904, v_905, v_906, v_907, v_908, v_909, v_910, v_911, v_912, v_913, v_914, v_915, v_916, v_917, v_918, v_919, v_920, v_921, v_922, v_923, v_924, v_925, v_926, v_927, v_928, v_929, v_930, v_931, v_932, v_933, v_934, v_935, v_936, v_937, v_938, v_939, v_940, v_941, v_942, v_943, v_944, v_945, v_946, v_947, v_948, v_949, v_950, v_951, v_952, v_953, v_954, v_955, v_956, v_957, v_958, v_959, v_960, v_961, v_962, v_963, v_964, v_965, v_966, v_967, v_968, v_969, v_970, v_971, v_972, v_973, v_974, v_975, v_976, v_977, v_978, v_979, v_980, v_981, v_982, v_983, v_984, v_985, v_986, v_987, v_988, v_989, v_990, v_991, v_992, v_993, v_994, v_995, v_996, v_997, v_998, v_999, v_1000, v_1001, v_1002, v_1003, v_1004, v_1005, v_1006, v_1007, v_1008, v_1009, v_1010, v_1011, v_1012, v_1013, v_1014, v_1015, v_1016, v_1017, v_1018, v_1019, v_1020, v_1021, v_1022, v_1023, v_1024, v_1025, v_1026, v_1027, v_1028, v_1029, v_1030, v_1031, v_1032, v_1033, v_1034, v_1035, v_1036, v_1037, v_1038, v_1039, v_1040, v_1041, v_1042, v_1043, v_1044, v_1045, v_1046, v_1047, v_1048, v_1049, v_1050, v_1051, v_1052, v_1053, v_1054, v_1055, v_1056, v_1057, v_1058, v_1059, v_1060, v_1061, v_1062, v_1063, v_1064, v_1065, v_1066, v_1067, v_1068, v_1069, v_1070, v_1071, v_1072, v_1073, v_1074, v_1075, v_1076, v_1077, v_1078, v_1079, v_1080, v_1081, v_1082, v_1083, v_1084, v_1085, v_1086, v_1087, v_1088, v_1089, v_1090, v_1091, v_1092, v_1093, v_1094, v_1095, v_1096, v_1097, v_1098, v_1099, v_1100, v_1101, v_1102, v_1103, v_1104, v_1105, v_1106, v_1107, v_1108, v_1109, v_1110, v_1111, v_1112, v_1113, v_1114, v_1115, v_1116, v_1117, v_1118, v_1119, v_1120, v_1121, v_1122, v_1123, v_1124, v_1125, v_1126, v_1127, v_1128, v_1129, v_1130, v_1131, v_1132, v_1133, v_1134, v_1135, v_1136, v_1137, v_1138, v_1139, v_1140, v_1141, v_1142, v_1143, v_1144, v_1145, v_1146, v_1147, v_1148, v_1149, v_1150, v_1151, v_1152, v_1153, v_1154, v_1155, v_1156, v_1157, v_1158, v_1159, v_1160, v_1161, v_1162, v_1163, v_1164, v_1165, v_1166, v_1167, v_1168, v_1169, v_1170, v_1171, v_1172, v_1173, v_1174, v_1175, v_1176, v_1177, v_1178, v_1179, v_1180, v_1181, v_1182, v_1183, v_1184, v_1185, v_1186, v_1187, v_1188, v_1189, v_1190, v_1191, v_1192, v_1193, v_1194, v_1195, v_1196, v_1197, v_1198, v_1199, v_1200, v_1201, v_1202, v_1203, v_1204, v_1205, v_1206, v_1207, v_1208, v_1209, v_1210, v_1211, v_1212, v_1213, v_1214, v_1215, v_1216, v_1217, v_1218, v_1219, v_1220, v_1221, v_1222, v_1223, v_1224, v_1225, v_1226, v_1227, v_1228, v_1229, v_1230, v_1231, v_1232, v_1233, v_1234, v_1235, v_1236, v_1237, v_1238, v_1239, v_1240, v_1241, v_1242, v_1243, v_1244, v_1245, v_1246, v_1247, v_1248, v_1249, v_1250, v_1251, v_1252, v_1253, v_1254, v_1255, v_1256, v_1257, v_1258, v_1259, v_1260, v_1261, v_1262, v_1263, v_1264, v_1265, v_1266, v_1267, v_1268, v_1269, v_1270, v_1271, v_1272, v_1273, v_1274, v_1275, v_1276, v_1277, v_1278, v_1279, v_1280, v_1281, v_1282, v_1283, v_1284, v_1285, v_1286, v_1287, v_1288, v_1289, v_1290, v_1291, v_1292, v_1293, v_1294, v_1295, v_1296, v_1297, v_1298, v_1299, v_1300, v_1301, v_1302, v_1303, v_1304, v_1305, v_1306, v_1307, v_1308, v_1309, v_1310, v_1311, v_1312, v_1313, v_1314, v_1315, v_1316, v_1317, v_1318, v_1319, v_1320, v_1321, v_1322, v_1323, v_1324, v_1325, v_1326, v_1327, v_1328, v_1329, v_1330, v_1331, v_1332, v_1333, v_1334, v_1335, v_1336, v_1337, v_1338, v_1339, v_1340, v_1341, v_1342, v_1343, v_1344, v_1345, v_1346, v_1347, v_1348, v_1349, v_1350, v_1351, v_1352, v_1353, v_1354, v_1355, v_1356, v_1357, v_1358, v_1359, v_1360, v_1361, v_1362, v_1363, v_1364, v_1365, v_1366, v_1367, v_1368, v_1369, v_1370, v_1371, v_1372, v_1373, v_1374, v_1375, v_1376, v_1377, v_1378, v_1379, v_1380, v_1381, v_1382, v_1383, v_1384, v_1385, v_1386, v_1387, v_1388, v_1389, v_1390, v_1391, v_1392, v_1393, v_1394, v_1395, v_1396, v_1397, v_1398, v_1399, v_1400, v_1401, v_1402, v_1403, v_1404, v_1405, v_1406, v_1407, v_1408, v_1409, v_1410, v_1411, v_1412, v_1413, v_1414, v_1415, v_1416, v_1417, v_1418, v_1419, v_1420, v_1421, v_1422, v_1423, v_1424, v_1425, v_1426, v_1427, v_1428, v_1429, v_1430, v_1431, v_1432, v_1433, v_1434, v_1435, v_1436, v_1437, v_1438, v_1439, v_1440, v_1441, v_1442, v_1443, v_1444, v_1445, v_1446, v_1447, v_1448, v_1449, v_1450, v_1451, v_1452, v_1453, v_1454, v_1455, v_1456, v_1457, v_1458, v_1459, v_1460, v_1461, v_1462, v_1463, v_1464, v_1465, v_1466, v_1467, v_1468, v_1469, v_1470, v_1471, v_1472, v_1473, v_1474, v_1475, v_1476, v_1477, v_1478, v_1479, v_1480, v_1481, v_1482, v_1483, v_1484, v_1485, v_1486, v_1487, v_1488, v_1489, v_1490, v_1491, v_1492, v_1493, v_1494, v_1495, v_1496, v_1497, v_1498, v_1499, v_1500, v_1501, v_1502, v_1503, v_1504, v_1505, v_1506, v_1507, v_1508, v_1509, v_1510, v_1511, v_1512, v_1513, v_1514, v_1515, v_1516, v_1517, v_1518, v_1519, v_1520, v_1521, v_1522, v_1523, v_1524, v_1525, v_1526, v_1527, v_1528, v_1529, v_1530, v_1531, v_1532, v_1533, v_1534, v_1535, v_1536, v_1537, v_1538, v_1539, v_1540, v_1541, v_1542, v_1543, v_1544, v_1545, v_1546, v_1547, v_1548, v_1549, v_1550, v_1551, v_1552, v_1553, v_1554, v_1555, v_1556, v_1557, v_1558, v_1559, v_1560, v_1561, v_1562, v_1563, v_1564, v_1565, v_1566, v_1567, v_1568, v_1569, v_1570, v_1571, v_1572, v_1573, v_1574, v_1575, v_1576, v_1577, v_1578, v_1579, v_1580, v_1581, v_1582, v_1583, v_1584, v_1585, v_1586, v_1587, v_1588, v_1589, v_1590, v_1591, v_1592, v_1593, v_1594, v_1595, v_1596, v_1597, v_1598, v_1599, v_1600, v_1601, v_1602, v_1603, v_1604, v_1605, v_1606, v_1607, v_1608, v_1609, v_1610, v_1611, v_1612, v_1613, v_1614, v_1615, v_1616, v_1617, v_1618, v_1619, v_1620, v_1621, v_1622, v_1623, v_1624, v_1625, v_1626, v_1627, v_1628, v_1629, v_1630, v_1631, v_1632, v_1633, v_1634, v_1635, v_1636, v_1637, v_1638, v_1639, v_1640, v_1641, v_1642, v_1643, v_1644, v_1645, v_1646, v_1647, v_1648, v_1649, v_1650, v_1651, v_1652, v_1653, v_1654, v_1655, v_1656, v_1657, v_1658, v_1659, v_1660, v_1661, v_1662, v_1663, v_1664, v_1665, v_1666, v_1667, v_1668, v_1669, v_1670, v_1671, v_1672, v_1673, v_1674, v_1675, v_1676, v_1677, v_1678, v_1679, v_1680, v_1681, v_1682, v_1683, v_1684, v_1685, v_1686, v_1687, v_1688, v_1689, v_1690, v_1691, v_1692, v_1693, v_1694, v_1695, v_1696, v_1697, v_1698, v_1699, v_1700, v_1701, v_1702, v_1703, v_1704, v_1705, v_1706, v_1707, v_1708, v_1709, v_1710, v_1711, v_1712, v_1713, v_1714, v_1715, v_1716, v_1717, v_1718, v_1719, v_1720, v_1721, v_1722, v_1723, v_1724, v_1725, v_1726, v_1727, v_1728, v_1729, v_1730, v_1731, v_1732, v_1733, v_1734, v_1735, v_1736, v_1737, v_1738, v_1739, v_1740, v_1741, v_1742, v_1743, v_1744, v_1745, v_1746, v_1747, v_1748, v_1749, v_1750, v_1751, v_1752, v_1753, v_1754, v_1755, v_1756, v_1757, v_1758, v_1759, v_1760, v_1761, v_1762, v_1763, v_1764, v_1765, v_1766, v_1767, v_1768, v_1769, v_1770, v_1771, v_1772, v_1773, v_1774, v_1775, v_1776, v_1777, v_1778, v_1779, v_1780, v_1781, v_1782, v_1783, v_1784, v_1785, v_1786, v_1787, v_1788, v_1789, v_1790, v_1791, v_1792, v_1793, v_1794, v_1795, v_1796, v_1797, v_1798, v_1799, v_1800, v_1801, v_1802, v_1803, v_1804, v_1805, v_1806, v_1807, v_1808, v_1809, v_1810, v_1811, v_1812, v_1813, v_1814, v_1815, v_1816, v_1817, v_1818, v_1819, v_1820, v_1821, v_1822, v_1823, v_1824, v_1825, v_1826, v_1827, v_1828, v_1829, v_1830, v_1831, v_1832, v_1833, v_1834, v_1835, v_1836, v_1837, v_1838, v_1839, v_1840, v_1841, v_1842, v_1843, v_1844, v_1845, v_1846, v_1847, v_1848, v_1849, v_1850, v_1851, v_1852, v_1853, v_1854, v_1855, v_1856, v_1857, v_1858, v_1859, v_1860, v_1861, v_1862, v_1863, v_1864, v_1865, v_1866, v_1867, v_1868, v_1869, v_1870, v_1871, v_1872, v_1873, v_1874, v_1875, v_1876, v_1877, v_1878, v_1879, v_1880, v_1881, v_1882, v_1883, v_1884, v_1885, v_1886, v_1887, v_1888, v_1889, v_1890, v_1891, v_1892, v_1893, v_1894, v_1895, v_1896, v_1897, v_1898, v_1899, v_1900, v_1901, v_1902, v_1903, v_1904, v_1905, v_1906, v_1907, v_1908, v_1909, v_1910, v_1911, v_1912, v_1913, v_1914, v_1915, v_1916, v_1917, v_1918, v_1919, v_1920, v_1921, v_1922, v_1923, v_1924, v_1925, v_1926, v_1927, v_1928, v_1929, v_1930, v_1931, v_1932, v_1933, v_1934, v_1935, v_1936, v_1937, v_1938, v_1939, v_1940, v_1941, v_1942, v_1943, v_1944, v_1945, v_1946, v_1947, v_1948, v_1949, v_1950, v_1951, v_1952, v_1953, v_1954, v_1955, v_1956, v_1957, v_1958, v_1959, v_1960, v_1961, v_1962, v_1963, v_1964, v_1965, v_1966, v_1967, v_1968, v_1969, v_1970, v_1971, v_1972, v_1973, v_1974, v_1975, v_1976, v_1977, v_1978, v_1979, v_1980, v_1981, v_1982, v_1983, v_1984, v_1985, v_1986, v_1987, v_1988, v_1989, v_1990, v_1991, v_1992, v_1993, v_1994, v_1995, v_1996, v_1997, v_1998, v_1999, v_2000, v_2001, v_2002, v_2003, v_2004, v_2005, v_2006, v_2007, v_2008, v_2009, v_2010, v_2011, v_2012, v_2013, v_2014, v_2015, v_2016, v_2017, v_2018, v_2019, v_2020, v_2021, v_2022, v_2023, v_2024, v_2025, v_2026, v_2027, v_2028, v_2029, v_2030, v_2031, v_2032, v_2033, v_2034, v_2035, v_2036, v_2037, v_2038, v_2039, v_2040, v_2041, v_2042, v_2043, v_2044, v_2045, v_2046, v_2047, v_2048, v_2049, v_2050, v_2051, v_2052, v_2053, v_2054, v_2055, v_2056, v_2057, v_2058, v_2059, v_2060, v_2061, v_2062, v_2063, v_2064, v_2065, v_2066, v_2067, v_2068, v_2069, v_2070, v_2071, v_2072, v_2073, v_2074, v_2075, v_2076, v_2077, v_2078, v_2079, v_2080, v_2081, v_2082, v_2083, v_2084, v_2085, v_2086, v_2087, v_2088, v_2089, v_2090, v_2091, v_2092, v_2093, v_2094, v_2095, v_2096, v_2097, v_2098, v_2099, v_2100, v_2101, v_2102, v_2103, v_2104, v_2105, v_2106, v_2107, v_2108, v_2109, v_2110, v_2111, v_2112, v_2113, v_2114, v_2115, v_2116, v_2117, v_2118, v_2119, v_2120, v_2121, v_2122, v_2123, v_2124, v_2125, v_2126, v_2127, v_2128, v_2129, v_2130, v_2131, v_2132, v_2133, v_2134, v_2135, v_2136, v_2137, v_2138, v_2139, v_2140, v_2141, v_2142, v_2143, v_2144, v_2145, v_2146, v_2147, v_2148, v_2149, v_2150, v_2151, v_2152, v_2153, v_2154, v_2155, v_2156, v_2157, v_2158, v_2159, v_2160, v_2161, v_2162, v_2163, v_2164, v_2165, v_2166, v_2167, v_2168, v_2169, v_2170, v_2171, v_2172, v_2173, v_2174, v_2175, v_2176, v_2177, v_2178, v_2179, v_2180, v_2181, v_2182, v_2183, v_2184, v_2185, v_2186, v_2187, v_2188, v_2189, v_2190, v_2191, v_2192, v_2193, v_2194, v_2195, v_2196, v_2197, v_2198, v_2199, v_2200, v_2201, v_2202, v_2203, v_2204, v_2205, v_2206, v_2207, v_2208, v_2209, v_2210, v_2211, v_2212, v_2213, v_2214, v_2215, v_2216, v_2217, v_2218, v_2219, v_2220, v_2221, v_2222, v_2223, v_2224, v_2225, v_2226, v_2227, v_2228, v_2229, v_2230, v_2231, v_2232, v_2233, v_2234, v_2235, v_2236, v_2237, v_2238, v_2239, v_2240, v_2241, v_2242, v_2243, v_2244, v_2245, v_2246, v_2247, v_2248, v_2249, v_2250, v_2251, v_2252, v_2253, v_2254, v_2255, v_2256, v_2257, v_2258, v_2259, v_2260, v_2261, v_2262, v_2263, v_2264, v_2265, v_2266, v_2267, v_2268, v_2269, v_2270, v_2271, v_2272, v_2273, v_2274, v_2275, v_2276, v_2277, v_2278, v_2279, v_2280, v_2281, v_2282, v_2283, v_2284, v_2285, v_2286, v_2287, v_2288, v_2289, v_2290, v_2291, v_2292, v_2293, v_2294, v_2295, v_2296, v_2297, v_2298, v_2299, v_2300, v_2301, v_2302, v_2303, v_2304, v_2305, v_2306, v_2307, v_2308, v_2309, v_2310, v_2311, v_2312, v_2313, v_2314, v_2315, v_2316, v_2317, v_2318, v_2319, v_2320, v_2321, v_2322, v_2323, v_2324, v_2325, v_2326, v_2327, v_2328, v_2329, v_2330, v_2331, v_2332, v_2333, v_2334, v_2335, v_2336, v_2337, v_2338, v_2339, v_2340, v_2341, v_2342, v_2343, v_2344, v_2345, v_2346, v_2347, v_2348, v_2349, v_2350, v_2351, v_2352, v_2353, v_2354, v_2355, v_2356, v_2357, v_2358, v_2359, v_2360, v_2361, v_2362, v_2363, v_2364, v_2365, v_2366, v_2367, v_2368, v_2369, v_2370, v_2371, v_2372, v_2373, v_2374, v_2375, v_2376, v_2377, v_2378, v_2379, v_2380, v_2381, v_2382, v_2383, v_2384, v_2385, v_2386, v_2387, v_2388, v_2389, v_2390, v_2391, v_2392, v_2393, v_2394, v_2395, v_2396, v_2397, v_2398, v_2399, v_2400, v_2401, v_2402, v_2403, v_2404, v_2405, v_2406, v_2407, v_2408, v_2409, v_2410, v_2411, v_2412, v_2413, v_2414, v_2415, v_2416, v_2417, v_2418, v_2419, v_2420, v_2421, v_2422, v_2423, v_2424, v_2425, v_2426, v_2427, v_2428, v_2429, v_2430, v_2431, v_2432, v_2433, v_2434, v_2435, v_2436, v_2437, v_2438, v_2439, v_2440, v_2441, v_2442, v_2443, v_2444, v_2445, v_2446, v_2447, v_2448, v_2449, v_2450, v_2451, v_2452, v_2453, v_2454, v_2455, v_2456, v_2457, v_2458, v_2459, v_2460, v_2461, v_2462, v_2463, v_2464, v_2465, v_2466, v_2467, v_2468, v_2469, v_2470, v_2471, v_2472, v_2473, v_2474, v_2475, v_2476, v_2477, v_2478, v_2479, v_2480, v_2481, v_2482, v_2483, v_2484, v_2485, v_2486, v_2487, v_2488, v_2489, v_2490, v_2491, v_2492, v_2493, v_2494, v_2495, v_2496, v_2497, v_2498, v_2499, v_2500, v_2501, v_2502, v_2503, v_2504, v_2505, v_2506, v_2507, v_2508, v_2509, v_2510, v_2511, v_2512, v_2513, v_2514, v_2515, v_2516, v_2517, v_2518, v_2519, v_2520, v_2521, v_2522, v_2523, v_2524, v_2525, v_2526, v_2527, v_2528, v_2529, v_2530, v_2531, v_2532, v_2533, v_2534, v_2535, v_2536, v_2537, v_2538, v_2539, v_2540, v_2541, v_2542, v_2543, v_2544, v_2545, v_2546, v_2547, v_2548, v_2549, v_2550, v_2551, v_2552, v_2553, v_2554, v_2555, v_2556, v_2557, v_2558, v_2559, v_2560, v_2561, v_2562, v_2563, v_2564, v_2565, v_2566, v_2567, v_2568, v_2569, v_2570, v_2571, v_2572, v_2573, v_2574, v_2575, v_2576, v_2577, v_2578, v_2579, v_2580, v_2581, v_2582, v_2583, v_2584, v_2585, v_2586, v_2587, v_2588, v_2589, v_2590, v_2591, v_2592, v_2593, v_2594, v_2595, v_2596, v_2597, v_2598, v_2599, v_2600, v_2601, v_2602, v_2603, v_2604, v_2605, v_2606, v_2607, v_2608, v_2609, v_2610, v_2611, v_2612, v_2613, v_2614, v_2615, v_2616, v_2617, v_2618, v_2619, v_2620, v_2621, v_2622, v_2623, v_2624, v_2625, v_2626, v_2627, v_2628, v_2629, v_2630, v_2631, v_2632, v_2633, v_2634, v_2635, v_2636, v_2637, v_2638, v_2639, v_2640, v_2641, v_2642, v_2643, v_2644, v_2645, v_2646, v_2647, v_2648, v_2649, v_2650, v_2651, v_2652, v_2653, v_2654, v_2655, v_2656, v_2657, v_2658, v_2659, v_2660, v_2661, v_2662, v_2663, v_2664, v_2665, v_2666, v_2667, v_2668, v_2669, v_2670, v_2671, v_2672, v_2673, v_2674, v_2675, v_2676, v_2677, v_2678, v_2679, v_2680, v_2681, v_2682, v_2683, v_2684, v_2685, v_2686, v_2687, v_2688, v_2689, v_2690, v_2691, v_2692, v_2693, v_2694, v_2695, v_2696, v_2697, v_2698, v_2699, v_2700, v_2701, v_2702, v_2703, v_2704, v_2705, v_2706, v_2707, v_2708, v_2709, v_2710, v_2711, v_2712, v_2713, v_2714, v_2715, v_2716, v_2717, v_2718, v_2719, v_2720, v_2721, v_2722, v_2723, v_2724, v_2725, v_2726, v_2727, v_2728, v_2729, v_2730, v_2731, v_2732, v_2733, v_2734, v_2735, v_2736, v_2737, v_2738, v_2739, v_2740, v_2741, v_2742, v_2743, v_2744, v_2745, v_2746, v_2747, v_2748, v_2749, v_2750, v_2751, v_2752, v_2753, v_2754, v_2755, v_2756, v_2757, v_2758, v_2759, v_2760, v_2761, v_2762, v_2763, v_2764, v_2765, v_2766, v_2767, v_2768, v_2769, v_2770, v_2771, v_2772, v_2773, v_2774, v_2775, v_2776, v_2777, v_2778, v_2779, v_2780, v_2781, v_2782, v_2783, v_2784, v_2785, v_2786, v_2787, v_2788, v_2789, v_2790, v_2791, v_2792, v_2793, v_2794, v_2795, v_2796, v_2797, v_2798, v_2799, v_2800, v_2801, v_2802, v_2803, v_2804, v_2805, v_2806, v_2807, v_2808, v_2809, v_2810, v_2811, v_2812, v_2813, v_2814, v_2815, v_2816, v_2817, v_2818, v_2819, v_2820, v_2821, v_2822, v_2823, v_2824, v_2825, v_2826, v_2827, v_2828, v_2829, v_2830, v_2831, v_2832, v_2833, v_2834, v_2835, v_2836, v_2837, v_2838, v_2839, v_2840, v_2841, v_2842, v_2843, v_2844, v_2845, v_2846, v_2847, v_2848, v_2849, v_2850, v_2851, v_2852, v_2853, v_2854, v_2855, v_2856, v_2857, v_2858, v_2859, v_2860, v_2861, v_2862, v_2863, v_2864, v_2865, v_2866, v_2867, v_2868, v_2869, v_2870, v_2871, v_2872, v_2873, v_2874, v_2875, v_2876, v_2877, v_2878, v_2879, v_2880, v_2881, v_2882, v_2883, v_2884, v_2885, v_2886, v_2887, v_2888, v_2889, v_2890, v_2891, v_2892, v_2893, v_2894, v_2895, v_2896, v_2897, v_2898, v_2899, v_2900, v_2901, v_2902, v_2903, v_2904, v_2905, v_2906, v_2907, v_2908, v_2909, v_2910, v_2911, v_2912, v_2913, v_2914, v_2915, v_2916, v_2917, v_2918, v_2919, v_2920, v_2921, v_2922, v_2923, v_2924, v_2925, v_2926, v_2927, v_2928, v_2929, v_2930, v_2931, v_2932, v_2933, v_2934, v_2935, v_2936, v_2937, v_2938, v_2939, v_2940, v_2941, v_2942, v_2943, v_2944, v_2945, v_2946, v_2947, v_2948, v_2949, v_2950, v_2951, v_2952, v_2953, v_2954, v_2955, v_2956, v_2957, v_2958, v_2959, v_2960, v_2961, v_2962, v_2963, v_2964, v_2965, v_2966, v_2967, v_2968, v_2969, v_2970, v_2971, v_2972, v_2973, v_2974, v_2975, v_2976, v_2977, v_2978, v_2979, v_2980, v_2981, v_2982, v_2983, v_2984, v_2985, v_2986, v_2987, v_2988, v_2989, v_2990, v_2991, v_2992, v_2993, v_2994, v_2995, v_2996, v_2997, v_2998, v_2999, v_3000, v_3001, v_3002, v_3003, v_3004, v_3005, v_3006, v_3007, v_3008, v_3009, v_3010, v_3011, v_3012, v_3013, v_3014, v_3015, v_3016, v_3017, v_3018, v_3019, v_3020, v_3021, v_3022, v_3023, v_3024, v_3025, v_3026, v_3027, v_3028, v_3029, v_3030, v_3031, v_3032, v_3033, v_3034, v_3035, v_3036, v_3037, v_3038, v_3039, v_3040, v_3041, v_3042, v_3043, v_3044, v_3045, v_3046, v_3047, v_3048, v_3049, v_3050, v_3051, v_3052, v_3053, v_3054, v_3055, v_3056, v_3057, v_3058, v_3059, v_3060, v_3061, v_3062, v_3063, v_3064, v_3065, v_3066, v_3067, v_3068, v_3069, v_3070, v_3071, v_3072, v_3073, v_3074, v_3075, v_3076, v_3077, v_3078, v_3079, v_3080, v_3081, v_3082, v_3083, v_3084, v_3085, v_3086, v_3087, v_3088, v_3089, v_3090, v_3091, v_3092, v_3093, v_3094, v_3095, v_3096, v_3097, v_3098, v_3099, v_3100, v_3101, v_3102, v_3103, v_3104, v_3105, v_3106, v_3107, v_3108, v_3109, v_3110, v_3111, v_3112, v_3113, v_3114, v_3115, v_3116, v_3117, v_3118, v_3119, v_3120, v_3121, v_3122, v_3123, v_3124, v_3125, v_3126, v_3127, v_3128, v_3129, v_3130, v_3131, v_3132, v_3133, v_3134, v_3135, v_3136, v_3137, v_3138, v_3139, v_3140, v_3141, v_3142, v_3143, v_3144, v_3145, v_3146, v_3147, v_3148, v_3149, v_3150, v_3151, v_3152, v_3153, v_3154, v_3155, v_3156, v_3157, v_3158, v_3159, v_3160, v_3161, v_3162, v_3163, v_3164, v_3165, v_3166, v_3167, v_3168, v_3169, v_3170, v_3171, v_3172, v_3173, v_3174, v_3175, v_3176, v_3177, v_3178, v_3179, v_3180, v_3181, v_3182, v_3183, v_3184, v_3185, v_3186, v_3187, v_3188, v_3189, v_3190, v_3191, v_3192, v_3193, v_3194, v_3195, v_3196, v_3197, v_3198, v_3199, v_3200, v_3201, v_3202, v_3203, v_3204, v_3205, v_3206, v_3207, v_3208, v_3209, v_3210, v_3211, v_3212, v_3213, v_3214, v_3215, v_3216, v_3217, v_3218, v_3219, v_3220, v_3221, v_3222, v_3223, v_3224, v_3225, v_3226, v_3227, v_3228, v_3229, v_3230, v_3231, v_3232, v_3233, v_3234, v_3235, v_3236, v_3237, v_3238, v_3239, v_3240, v_3241, v_3242, v_3243, v_3244, v_3245, v_3246, v_3247, v_3248, v_3249, v_3250, v_3251, v_3252, v_3253, v_3254, v_3255, v_3256, v_3257, v_3258, v_3259, v_3260, v_3261, v_3262, v_3263, v_3264, v_3265, v_3266, v_3267, v_3268, v_3269, v_3270, v_3271, v_3272, v_3273, v_3274, v_3275, v_3276, v_3277, v_3278, v_3279, v_3280, v_3281, v_3282, v_3283, v_3284, v_3285, v_3286, v_3287, v_3288, v_3289, v_3290, v_3291, v_3292, v_3293, v_3294, v_3295, v_3296, v_3297, v_3298, v_3299, v_3300, v_3301, v_3302, v_3303, v_3304, v_3305, v_3306, v_3307, v_3308, v_3309, v_3310, v_3311, v_3312, v_3313, v_3314, v_3315, v_3316, v_3317, v_3318, v_3319, v_3320, v_3321, v_3322, v_3323, v_3324, v_3325, v_3326, v_3327, v_3328, v_3329, v_3330, v_3331, v_3332, v_3333, v_3334, v_3335, v_3336, v_3337, v_3338, v_3339, v_3340, v_3341, v_3342, v_3343, v_3344, v_3345, v_3346, v_3347, v_3348, v_3349, v_3350, v_3351, v_3352, v_3353, v_3354, v_3355, v_3356, v_3357, v_3358, v_3359, v_3360, v_3361, v_3362, v_3363, v_3364, v_3365, v_3366, v_3367, v_3368, v_3369, v_3370, v_3371, v_3372, v_3373, v_3374, v_3375, v_3376, v_3377, v_3378, v_3379, v_3380, v_3381, v_3382, v_3383, v_3384, v_3385, v_3386, v_3387, v_3388, v_3389, v_3390, v_3391, v_3392, v_3393, v_3394, v_3395, v_3396, v_3397, v_3398, v_3399, v_3400, v_3401, v_3402, v_3403, v_3404, v_3405, v_3406, v_3407, v_3408, v_3409, v_3410, v_3411, v_3412, v_3413, v_3414, v_3415, v_3416, v_3417, v_3418, v_3419, v_3420, v_3421, v_3422, v_3423, v_3424, v_3425, v_3426, v_3427, v_3428, v_3429, v_3430, v_3431, v_3432, v_3433, v_3434, v_3435, v_3436, v_3437, v_3438, v_3439, v_3440, v_3441, v_3442, v_3443, v_3444, v_3445, v_3446, v_3447, v_3448, v_3449, v_3450, v_3451, v_3452, v_3453, v_3454, v_3455, v_3456, v_3457, v_3458, v_3459, v_3460, v_3461, v_3462, v_3463, v_3464, v_3465, v_3466, v_3467, v_3468, v_3469, v_3470, v_3471, v_3472, v_3473, v_3474, v_3475, v_3476, v_3477, v_3478, v_3479, v_3480, v_3481, v_3482, v_3483, v_3484, v_3485, v_3486, v_3487, v_3488, v_3489, v_3490, v_3491, v_3492, v_3493, v_3494, v_3495, v_3496, v_3497, v_3498, v_3499, v_3500, v_3501, v_3502, v_3503, v_3504, v_3505, v_3506, v_3507, v_3508, v_3509, v_3510, v_3511, v_3512, v_3513, v_3514, v_3515, v_3516, v_3517, v_3518, v_3519, v_3520, v_3521, v_3522, v_3523, v_3524, v_3525, v_3526, v_3527, v_3528, v_3529, v_3530, v_3531, v_3532, v_3533, v_3534, v_3535, v_3536, v_3537, v_3538, v_3539, v_3540, v_3541, v_3542, v_3543, v_3544, v_3545, v_3546, v_3547, v_3548, v_3549, v_3550, v_3551, v_3552, v_3553, v_3554, v_3555, v_3556, v_3557, v_3558, v_3559, v_3560, v_3561, v_3562, v_3563, v_3564, v_3565, v_3566, v_3567, v_3568, v_3569, v_3570, v_3571, v_3572, v_3573, v_3574, v_3575, v_3576, v_3577, v_3578, v_3579, v_3580, v_3581, v_3582, v_3583, v_3584, v_3585, v_3586, v_3587, v_3588, v_3589, v_3590, v_3591, v_3592, v_3593, v_3594, v_3595, v_3596, v_3597, v_3598, v_3599, v_3600, v_3601, v_3602, v_3603, v_3604, v_3605, v_3606, v_3607, v_3608, v_3609, v_3610, v_3611, v_3612, v_3613, v_3614, v_3615, v_3616, v_3617, v_3618, v_3619, v_3620, v_3621, v_3622, v_3623, v_3624, v_3625, v_3626, v_3627, v_3628, v_3629, v_3630, v_3631, v_3632, v_3633, v_3634, v_3635, v_3636, v_3637, v_3638, v_3639, v_3640, v_3641, v_3642, v_3643, v_3644, v_3645, v_3646, v_3647, v_3648, v_3649, v_3650, v_3651, v_3652, v_3653, v_3654, v_3655, v_3656, v_3657, v_3658, v_3659, v_3660, v_3661, v_3662, v_3663, v_3664, v_3665, v_3666, v_3667, v_3668, v_3669, v_3670, v_3671, v_3672, v_3673, v_3674, v_3675, v_3676, v_3677, v_3678, v_3679, v_3680, v_3681, v_3682, v_3683, v_3684, v_3685, v_3686, v_3687, v_3688, v_3689, v_3690, v_3691, v_3692, v_3693, v_3694, v_3695, v_3696, v_3697, v_3698, v_3699, v_3700, v_3701, v_3702, v_3703, v_3704, v_3705, v_3706, v_3707, v_3708, v_3709, v_3710, v_3711, v_3712, v_3713, v_3714, v_3715, v_3716, v_3717, v_3718, v_3719, v_3720, v_3721, v_3722, v_3723, v_3724, v_3725, v_3726, v_3727, v_3728, v_3729, v_3730, v_3731, v_3732, v_3733, v_3734, v_3735, v_3736, v_3737, v_3738, v_3739, v_3740, v_3741, v_3742, v_3743, v_3744, v_3745, v_3746, v_3747, v_3748, v_3749, v_3750, v_3751, v_3752, v_3753, v_3754, v_3755, v_3756, v_3757, v_3758, v_3759, v_3760, v_3761, v_3762, v_3763, v_3764, v_3765, v_3766, v_3767, v_3768, v_3769, v_3770, v_3771, v_3772, v_3773, v_3774, v_3775, v_3776, v_3777, v_3778, v_3779, v_3780, v_3781, v_3782, v_3783, v_3784, v_3785, v_3786, v_3787, v_3788, v_3789, v_3790, v_3791, v_3792, v_3793, v_3794, v_3795, v_3796, v_3797, v_3798, v_3799, v_3800, v_3801, v_3802, v_3803, v_3804, v_3805, v_3806, v_3807, v_3808, v_3809, v_3810, v_3811, v_3812, v_3813, v_3814, v_3815, v_3816, v_3817, v_3818, v_3819, v_3820, v_3821, v_3822, v_3823, v_3824, v_3825, v_3826, v_3827, v_3828, v_3829, v_3830, v_3831, v_3832, v_3833, v_3834, v_3835, v_3836, v_3837, v_3838, v_3839, v_3840, v_3841, v_3842, v_3843, v_3844, v_3845, v_3846, v_3847, v_3848, v_3849, v_3850, v_3851, v_3852, v_3853, v_3854, v_3855, v_3856, v_3857, v_3858, v_3859, v_3860, v_3861, v_3862, v_3863, v_3864, v_3865, v_3866, v_3867, v_3868, v_3869, v_3870, v_3871, v_3872, v_3873, v_3874, v_3875, v_3876, v_3877, v_3878, v_3879, v_3880, v_3881, v_3882, v_3883, v_3884, v_3885, v_3886, v_3887, v_3888, v_3889, v_3890, v_3891, v_3892, v_3893, v_3894, v_3895, v_3896, v_3897, v_3898, v_3899, v_3900, v_3901, v_3902, v_3903, v_3904, v_3905, v_3906, v_3907, v_3908, v_3909, v_3910, v_3911, v_3912, v_3913, v_3914, v_3915, v_3916, v_3917, v_3918, v_3919, v_3920, v_3921, v_3922, v_3923, v_3924, v_3925, v_3926, v_3927, v_3928, v_3929, v_3930, v_3931, v_3932, v_3933, v_3934, v_3935, v_3936, v_3937, v_3938, v_3939, v_3940, v_3941, v_3942, v_3943, v_3944, v_3945, v_3946, v_3947, v_3948, v_3949, v_3950, v_3951, v_3952, v_3953, v_3954, v_3955, v_3956, v_3957, v_3958, v_3959, v_3960, v_3961, v_3962, v_3963, v_3964, v_3965, v_3966, v_3967, v_3968, v_3969, v_3970, v_3971, v_3972, v_3973, v_3974, v_3975, v_3976, v_3977, v_3978, v_3979, v_3980, v_3981, v_3982, v_3983, v_3984, v_3985, v_3986, v_3987, v_3988, v_3989, v_3990, v_3991, v_3992, v_3993, v_3994, v_3995, v_3996, v_3997, v_3998, v_3999, v_4000, v_4001, v_4002, v_4003, v_4004, v_4005, v_4006, v_4007, v_4008, v_4009, v_4010, v_4011, v_4012, v_4013, v_4014, v_4015, v_4016, v_4017, v_4018, v_4019, v_4020, v_4021, v_4022, v_4023, v_4024, v_4025, v_4026, v_4027, v_4028, v_4029, v_4030, v_4031, v_4032, v_4033, v_4034, v_4035, v_4036, v_4037, v_4038, v_4039, v_4040, v_4041, v_4042, v_4043, v_4044, v_4045, v_4046, v_4047, v_4048, v_4049, v_4050, v_4051, v_4052, v_4053, v_4054, v_4055, v_4056, v_4057, v_4058, v_4059, v_4060, v_4061, v_4062, v_4063, v_4064, v_4065, v_4066, v_4067, v_4068, v_4069, v_4070, v_4071, v_4072, v_4073, v_4074, v_4075, v_4076, v_4077, v_4078, v_4079, v_4080, v_4081, v_4082, v_4083, v_4084, v_4085, v_4086, v_4087, v_4088, v_4089, v_4090, v_4091, v_4092, v_4093, v_4094, v_4095, v_4096, v_4097, v_4098, v_4099, v_4100, v_4101, v_4102, v_4103, v_4104, v_4105, v_4106, v_4107, v_4108, v_4109, v_4110, v_4111, v_4112, v_4113, v_4114, v_4115, v_4116, v_4117, v_4118, v_4119, v_4120, v_4121, v_4122, v_4123, v_4124, v_4125, v_4126, v_4127, v_4128, v_4129, v_4130, v_4131, v_4132, v_4133, v_4134, v_4135, v_4136, v_4137, v_4138, v_4139, v_4140, v_4141, v_4142, v_4143, v_4144, v_4145, v_4146, v_4147, v_4148, v_4149, v_4150, v_4151, v_4152, v_4153, v_4154, v_4155, v_4156, v_4157, v_4158, v_4159, v_4160, v_4161, v_4162, v_4163, v_4164, v_4165, v_4166, v_4167, v_4168, v_4169, v_4170, v_4171, v_4172, v_4173, v_4174, v_4175, v_4176, v_4177, v_4178, v_4179, v_4180, v_4181, v_4182, v_4183, v_4184, v_4185, v_4186, v_4187, v_4188, v_4189, v_4190, v_4191, v_4192, v_4193, v_4194, v_4195, v_4196, v_4197, v_4198, v_4199, v_4200, v_4201, v_4202, v_4203, v_4204, v_4205, v_4206, v_4207, v_4208, v_4209, v_4210, v_4211, v_4212, v_4213, v_4214, v_4215, v_4216, v_4217, v_4218, v_4219, v_4220, v_4221, v_4222, v_4223, v_4224, v_4225, v_4226, v_4227, v_4228, v_4229, v_4230, v_4231, v_4232, v_4233, v_4234, v_4235, v_4236, v_4237, v_4238, v_4239, v_4240, v_4241, v_4242, v_4243, v_4244, v_4245, v_4246, v_4247, v_4248, v_4249, v_4250, v_4251, v_4252, v_4253, v_4254, v_4255, v_4256, v_4257, v_4258, v_4259, v_4260, v_4261, v_4262, v_4263, v_4264, v_4265, v_4266, v_4267, v_4268, v_4269, v_4270, v_4271, v_4272, v_4273, v_4274, v_4275, v_4276, v_4277, v_4278, v_4279, v_4280, v_4281, v_4282, v_4283, v_4284, v_4285, v_4286, v_4287, v_4288, v_4289, v_4290, v_4291, v_4292, v_4293, v_4294, v_4295, v_4296, v_4297, v_4298, v_4299, v_4300, v_4301, v_4302, v_4303, v_4304, v_4305, v_4306, v_4307, v_4308, v_4309, v_4310, v_4311, v_4312, v_4313, v_4314, v_4315, v_4316, v_4317, v_4318, v_4319, v_4320, v_4321, v_4322, v_4323, v_4324, v_4325, v_4326, v_4327, v_4328, v_4329, v_4330, v_4331, v_4332, v_4333, v_4334, v_4335, v_4336, v_4337, v_4338, v_4339, v_4340, v_4341, v_4342, v_4343, v_4344, v_4345, v_4346, v_4347, v_4348, v_4349, v_4350, v_4351, v_4352, v_4353, v_4354, v_4355, v_4356, v_4357, v_4358, v_4359, v_4360, v_4361, v_4362, v_4363, v_4364, v_4365, v_4366, v_4367, v_4368, v_4369, v_4370, v_4371, v_4372, v_4373, v_4374, v_4375, v_4376, v_4377, v_4378, v_4379, v_4380, v_4381, v_4382, v_4383, v_4384, v_4385, v_4386, v_4387, v_4388, v_4389, v_4390, v_4391, v_4392, v_4393, v_4394, v_4395, v_4396, v_4397, v_4398, v_4399, v_4400, v_4401, v_4402, v_4403, v_4404, v_4405, v_4406, v_4407, v_4408, v_4409, v_4410, v_4411, v_4412, v_4413, v_4414, v_4415, v_4416, v_4417, v_4418, v_4419, v_4420, v_4421, v_4422, v_4423, v_4424, v_4425, v_4426, v_4427, v_4428, v_4429, v_4430, v_4431, v_4432, v_4433, v_4434, v_4435, v_4436, v_4437, v_4438, v_4439, v_4440, v_4441, v_4442, v_4443, v_4444, v_4445, v_4446, v_4447, v_4448, v_4449, v_4450, v_4451, v_4452, v_4453, v_4454, v_4455, v_4456, v_4457, v_4458, v_4459, v_4460, v_4461, v_4462, v_4463, v_4464, v_4465, v_4466, v_4467, v_4468, v_4469, v_4470, v_4471, v_4472, v_4473, v_4474, v_4475, v_4476, v_4477, v_4478, v_4479, v_4480, v_4481, v_4482, v_4483, v_4484, v_4485, v_4486, v_4487, v_4488, v_4489, v_4490, v_4491, v_4492, v_4493, v_4494, v_4495, v_4496, v_4497, v_4498, v_4499, v_4500, v_4501, v_4502, v_4503, v_4504, v_4505, v_4506, v_4507, v_4508, v_4509, v_4510, v_4511, v_4512, v_4513, v_4514, v_4515, v_4516, v_4517, v_4518, v_4519, v_4520, v_4521, v_4522, v_4523, v_4524, v_4525, v_4526, v_4527, v_4528, v_4529, v_4530, v_4531, v_4532, v_4533, v_4534, v_4535, v_4536, v_4537, v_4538, v_4539, v_4540, v_4541, v_4542, v_4543, v_4544, v_4545, v_4546, v_4547, v_4548, v_4549, v_4550, v_4551, v_4552, v_4553, v_4554, v_4555, v_4556, v_4557, v_4558, v_4559, v_4560, v_4561, v_4562, v_4563, v_4564, v_4565, v_4566, v_4567, v_4568, v_4569, v_4570, v_4571, v_4572, v_4573, v_4574, v_4575, v_4576, v_4577, v_4578, v_4579, v_4580, v_4581, v_4582, v_4583, v_4584, v_4585, v_4586, v_4587, v_4588, o_1);
input v_1;
input v_2;
input v_3;
input v_4;
input v_5;
input v_6;
input v_7;
input v_8;
input v_9;
input v_10;
input v_11;
input v_12;
input v_13;
input v_14;
input v_15;
input v_16;
input v_17;
input v_18;
input v_20;
input v_21;
input v_22;
input v_23;
input v_24;
input v_25;
input v_26;
input v_27;
input v_28;
input v_29;
input v_30;
input v_31;
input v_32;
input v_33;
input v_34;
input v_35;
input v_36;
input v_37;
input v_38;
input v_39;
input v_40;
input v_41;
input v_42;
input v_43;
input v_44;
input v_45;
input v_46;
input v_47;
input v_48;
input v_49;
input v_50;
input v_51;
input v_52;
input v_53;
input v_54;
input v_55;
input v_56;
input v_57;
input v_58;
input v_59;
input v_60;
input v_61;
input v_62;
input v_63;
input v_64;
input v_65;
input v_66;
input v_67;
input v_68;
input v_69;
input v_70;
input v_71;
input v_72;
input v_73;
input v_74;
input v_75;
input v_76;
input v_77;
input v_78;
input v_79;
input v_80;
input v_81;
input v_82;
input v_83;
input v_84;
input v_85;
input v_86;
input v_87;
input v_88;
input v_89;
input v_90;
input v_91;
input v_92;
input v_93;
input v_94;
input v_95;
input v_96;
input v_97;
input v_98;
input v_99;
input v_100;
input v_101;
input v_102;
input v_103;
input v_104;
input v_105;
input v_106;
input v_107;
input v_108;
input v_109;
input v_110;
input v_111;
input v_112;
input v_113;
input v_114;
input v_115;
input v_116;
input v_117;
input v_118;
input v_119;
input v_120;
input v_121;
input v_122;
input v_123;
input v_124;
input v_125;
input v_126;
input v_127;
input v_128;
input v_129;
input v_130;
input v_131;
input v_132;
input v_133;
input v_134;
input v_135;
input v_136;
input v_137;
input v_138;
input v_142;
input v_143;
input v_144;
input v_145;
input v_146;
input v_147;
input v_148;
input v_149;
input v_150;
input v_151;
input v_155;
input v_159;
input v_160;
input v_161;
input v_162;
input v_163;
input v_164;
input v_165;
input v_166;
input v_167;
input v_168;
input v_169;
input v_170;
input v_171;
input v_172;
input v_179;
input v_180;
input v_181;
input v_182;
input v_183;
input v_184;
input v_19;
input v_139;
input v_140;
input v_141;
input v_152;
input v_153;
input v_154;
input v_156;
input v_157;
input v_158;
input v_173;
input v_174;
input v_175;
input v_176;
input v_177;
input v_178;
input v_185;
input v_186;
input v_187;
input v_188;
input v_189;
input v_190;
input v_191;
input v_192;
input v_193;
input v_194;
input v_195;
input v_196;
input v_197;
input v_198;
input v_199;
input v_200;
input v_201;
input v_202;
input v_203;
input v_204;
input v_205;
input v_206;
input v_207;
input v_208;
input v_209;
input v_210;
input v_211;
input v_212;
input v_213;
input v_214;
input v_215;
input v_216;
input v_217;
input v_218;
input v_219;
input v_220;
input v_221;
input v_222;
input v_223;
input v_224;
input v_225;
input v_226;
input v_227;
input v_228;
input v_229;
input v_230;
input v_231;
input v_232;
input v_233;
input v_234;
input v_235;
input v_236;
input v_237;
input v_238;
input v_239;
input v_240;
input v_241;
input v_242;
input v_243;
input v_244;
input v_245;
input v_246;
input v_247;
input v_248;
input v_249;
input v_250;
input v_251;
input v_252;
input v_253;
input v_254;
input v_255;
input v_256;
input v_257;
input v_258;
input v_259;
input v_260;
input v_261;
input v_262;
input v_263;
input v_264;
input v_265;
input v_266;
input v_267;
input v_268;
input v_269;
input v_270;
input v_271;
input v_272;
input v_273;
input v_274;
input v_275;
input v_276;
input v_277;
input v_278;
input v_279;
input v_280;
input v_281;
input v_282;
input v_283;
input v_284;
input v_285;
input v_286;
input v_287;
input v_288;
input v_289;
input v_290;
input v_291;
input v_292;
input v_293;
input v_294;
input v_295;
input v_296;
input v_297;
input v_298;
input v_299;
input v_300;
input v_301;
input v_302;
input v_303;
input v_304;
input v_305;
input v_306;
input v_307;
input v_308;
input v_309;
input v_310;
input v_311;
input v_312;
input v_313;
input v_314;
input v_315;
input v_316;
input v_317;
input v_318;
input v_319;
input v_320;
input v_321;
input v_322;
input v_323;
input v_324;
input v_325;
input v_326;
input v_327;
input v_328;
input v_329;
input v_330;
input v_331;
input v_332;
input v_333;
input v_334;
input v_335;
input v_336;
input v_337;
input v_338;
input v_339;
input v_340;
input v_341;
input v_342;
input v_343;
input v_344;
input v_345;
input v_346;
input v_347;
input v_348;
input v_349;
input v_350;
input v_351;
input v_352;
input v_353;
input v_354;
input v_355;
input v_356;
input v_357;
input v_358;
input v_359;
input v_360;
input v_361;
input v_362;
input v_363;
input v_364;
input v_365;
input v_366;
input v_367;
input v_368;
input v_369;
input v_370;
input v_371;
input v_372;
input v_373;
input v_374;
input v_375;
input v_376;
input v_377;
input v_378;
input v_379;
input v_380;
input v_381;
input v_382;
input v_383;
input v_384;
input v_385;
input v_386;
input v_387;
input v_388;
input v_389;
input v_390;
input v_391;
input v_392;
input v_393;
input v_394;
input v_395;
input v_396;
input v_397;
input v_398;
input v_399;
input v_400;
input v_401;
input v_402;
input v_403;
input v_404;
input v_405;
input v_406;
input v_407;
input v_408;
input v_409;
input v_410;
input v_411;
input v_412;
input v_413;
input v_414;
input v_415;
input v_416;
input v_417;
input v_418;
input v_419;
input v_420;
input v_421;
input v_422;
input v_423;
input v_424;
input v_425;
input v_426;
input v_427;
input v_428;
input v_429;
input v_430;
input v_431;
input v_432;
input v_433;
input v_434;
input v_435;
input v_436;
input v_437;
input v_438;
input v_439;
input v_440;
input v_441;
input v_442;
input v_443;
input v_444;
input v_445;
input v_446;
input v_447;
input v_448;
input v_449;
input v_450;
input v_451;
input v_452;
input v_453;
input v_454;
input v_455;
input v_456;
input v_457;
input v_458;
input v_459;
input v_460;
input v_461;
input v_462;
input v_463;
input v_464;
input v_465;
input v_466;
input v_467;
input v_468;
input v_469;
input v_470;
input v_471;
input v_472;
input v_473;
input v_474;
input v_475;
input v_476;
input v_477;
input v_478;
input v_479;
input v_480;
input v_481;
input v_482;
input v_483;
input v_484;
input v_485;
input v_486;
input v_487;
input v_488;
input v_489;
input v_490;
input v_491;
input v_492;
input v_493;
input v_494;
input v_495;
input v_496;
input v_497;
input v_498;
input v_499;
input v_500;
input v_501;
input v_502;
input v_503;
input v_504;
input v_505;
input v_506;
input v_507;
input v_508;
input v_509;
input v_510;
input v_511;
input v_512;
input v_513;
input v_514;
input v_515;
input v_516;
input v_517;
input v_518;
input v_519;
input v_520;
input v_521;
input v_522;
input v_523;
input v_524;
input v_525;
input v_526;
input v_527;
input v_528;
input v_529;
input v_530;
input v_531;
input v_532;
input v_533;
input v_534;
input v_535;
input v_536;
input v_537;
input v_538;
input v_539;
input v_540;
input v_541;
input v_542;
input v_543;
input v_544;
input v_545;
input v_546;
input v_547;
input v_548;
input v_549;
input v_550;
input v_551;
input v_552;
input v_553;
input v_554;
input v_555;
input v_556;
input v_557;
input v_558;
input v_559;
input v_560;
input v_561;
input v_562;
input v_563;
input v_564;
input v_565;
input v_566;
input v_567;
input v_568;
input v_569;
input v_570;
input v_571;
input v_572;
input v_573;
input v_574;
input v_575;
input v_576;
input v_577;
input v_578;
input v_579;
input v_580;
input v_581;
input v_582;
input v_583;
input v_584;
input v_585;
input v_586;
input v_587;
input v_588;
input v_589;
input v_590;
input v_591;
input v_592;
input v_593;
input v_594;
input v_595;
input v_596;
input v_597;
input v_598;
input v_599;
input v_600;
input v_601;
input v_602;
input v_603;
input v_604;
input v_605;
input v_606;
input v_607;
input v_608;
input v_609;
input v_610;
input v_611;
input v_612;
input v_613;
input v_614;
input v_615;
input v_616;
input v_617;
input v_618;
input v_619;
input v_620;
input v_621;
input v_622;
input v_623;
input v_624;
input v_625;
input v_626;
input v_627;
input v_628;
input v_629;
input v_630;
input v_631;
input v_632;
input v_633;
input v_634;
input v_635;
input v_636;
input v_637;
input v_638;
input v_639;
input v_640;
input v_641;
input v_642;
input v_643;
input v_644;
input v_645;
input v_646;
input v_647;
input v_648;
input v_649;
input v_650;
input v_651;
input v_652;
input v_653;
input v_654;
input v_655;
input v_656;
input v_657;
input v_658;
input v_659;
input v_660;
input v_661;
input v_662;
input v_663;
input v_664;
input v_665;
input v_666;
input v_667;
input v_668;
input v_669;
input v_670;
input v_671;
input v_672;
input v_673;
input v_674;
input v_675;
input v_676;
input v_677;
input v_678;
input v_679;
input v_680;
input v_681;
input v_682;
input v_683;
input v_684;
input v_685;
input v_686;
input v_687;
input v_688;
input v_689;
input v_690;
input v_691;
input v_692;
input v_693;
input v_694;
input v_695;
input v_696;
input v_697;
input v_698;
input v_699;
input v_700;
input v_701;
input v_702;
input v_703;
input v_704;
input v_705;
input v_706;
input v_707;
input v_708;
input v_709;
input v_710;
input v_711;
input v_712;
input v_713;
input v_714;
input v_715;
input v_716;
input v_717;
input v_718;
input v_719;
input v_720;
input v_721;
input v_722;
input v_723;
input v_724;
input v_725;
input v_726;
input v_727;
input v_728;
input v_729;
input v_730;
input v_731;
input v_732;
input v_733;
input v_734;
input v_735;
input v_736;
input v_737;
input v_738;
input v_739;
input v_740;
input v_741;
input v_742;
input v_743;
input v_744;
input v_745;
input v_746;
input v_747;
input v_748;
input v_749;
input v_750;
input v_751;
input v_752;
input v_753;
input v_754;
input v_755;
input v_756;
input v_757;
input v_758;
input v_759;
input v_760;
input v_761;
input v_762;
input v_763;
input v_764;
input v_765;
input v_766;
input v_767;
input v_768;
input v_769;
input v_770;
input v_771;
input v_772;
input v_773;
input v_774;
input v_775;
input v_776;
input v_777;
input v_778;
input v_779;
input v_780;
input v_781;
input v_782;
input v_783;
input v_784;
input v_785;
input v_786;
input v_787;
input v_788;
input v_789;
input v_790;
input v_791;
input v_792;
input v_793;
input v_794;
input v_795;
input v_796;
input v_797;
input v_798;
input v_799;
input v_800;
input v_801;
input v_802;
input v_803;
input v_804;
input v_805;
input v_806;
input v_807;
input v_808;
input v_809;
input v_810;
input v_811;
input v_812;
input v_813;
input v_814;
input v_815;
input v_816;
input v_817;
input v_818;
input v_819;
input v_820;
input v_821;
input v_822;
input v_823;
input v_824;
input v_825;
input v_826;
input v_827;
input v_828;
input v_829;
input v_830;
input v_831;
input v_832;
input v_833;
input v_834;
input v_835;
input v_836;
input v_837;
input v_838;
input v_839;
input v_840;
input v_841;
input v_842;
input v_843;
input v_844;
input v_845;
input v_846;
input v_847;
input v_848;
input v_849;
input v_850;
input v_851;
input v_852;
input v_853;
input v_854;
input v_855;
input v_856;
input v_857;
input v_858;
input v_859;
input v_860;
input v_861;
input v_862;
input v_863;
input v_864;
input v_865;
input v_866;
input v_867;
input v_868;
input v_869;
input v_870;
input v_871;
input v_872;
input v_873;
input v_874;
input v_875;
input v_876;
input v_877;
input v_878;
input v_879;
input v_880;
input v_881;
input v_882;
input v_883;
input v_884;
input v_885;
input v_886;
input v_887;
input v_888;
input v_889;
input v_890;
input v_891;
input v_892;
input v_893;
input v_894;
input v_895;
input v_896;
input v_897;
input v_898;
input v_899;
input v_900;
input v_901;
input v_902;
input v_903;
input v_904;
input v_905;
input v_906;
input v_907;
input v_908;
input v_909;
input v_910;
input v_911;
input v_912;
input v_913;
input v_914;
input v_915;
input v_916;
input v_917;
input v_918;
input v_919;
input v_920;
input v_921;
input v_922;
input v_923;
input v_924;
input v_925;
input v_926;
input v_927;
input v_928;
input v_929;
input v_930;
input v_931;
input v_932;
input v_933;
input v_934;
input v_935;
input v_936;
input v_937;
input v_938;
input v_939;
input v_940;
input v_941;
input v_942;
input v_943;
input v_944;
input v_945;
input v_946;
input v_947;
input v_948;
input v_949;
input v_950;
input v_951;
input v_952;
input v_953;
input v_954;
input v_955;
input v_956;
input v_957;
input v_958;
input v_959;
input v_960;
input v_961;
input v_962;
input v_963;
input v_964;
input v_965;
input v_966;
input v_967;
input v_968;
input v_969;
input v_970;
input v_971;
input v_972;
input v_973;
input v_974;
input v_975;
input v_976;
input v_977;
input v_978;
input v_979;
input v_980;
input v_981;
input v_982;
input v_983;
input v_984;
input v_985;
input v_986;
input v_987;
input v_988;
input v_989;
input v_990;
input v_991;
input v_992;
input v_993;
input v_994;
input v_995;
input v_996;
input v_997;
input v_998;
input v_999;
input v_1000;
input v_1001;
input v_1002;
input v_1003;
input v_1004;
input v_1005;
input v_1006;
input v_1007;
input v_1008;
input v_1009;
input v_1010;
input v_1011;
input v_1012;
input v_1013;
input v_1014;
input v_1015;
input v_1016;
input v_1017;
input v_1018;
input v_1019;
input v_1020;
input v_1021;
input v_1022;
input v_1023;
input v_1024;
input v_1025;
input v_1026;
input v_1027;
input v_1028;
input v_1029;
input v_1030;
input v_1031;
input v_1032;
input v_1033;
input v_1034;
input v_1035;
input v_1036;
input v_1037;
input v_1038;
input v_1039;
input v_1040;
input v_1041;
input v_1042;
input v_1043;
input v_1044;
input v_1045;
input v_1046;
input v_1047;
input v_1048;
input v_1049;
input v_1050;
input v_1051;
input v_1052;
input v_1053;
input v_1054;
input v_1055;
input v_1056;
input v_1057;
input v_1058;
input v_1059;
input v_1060;
input v_1061;
input v_1062;
input v_1063;
input v_1064;
input v_1065;
input v_1066;
input v_1067;
input v_1068;
input v_1069;
input v_1070;
input v_1071;
input v_1072;
input v_1073;
input v_1074;
input v_1075;
input v_1076;
input v_1077;
input v_1078;
input v_1079;
input v_1080;
input v_1081;
input v_1082;
input v_1083;
input v_1084;
input v_1085;
input v_1086;
input v_1087;
input v_1088;
input v_1089;
input v_1090;
input v_1091;
input v_1092;
input v_1093;
input v_1094;
input v_1095;
input v_1096;
input v_1097;
input v_1098;
input v_1099;
input v_1100;
input v_1101;
input v_1102;
input v_1103;
input v_1104;
input v_1105;
input v_1106;
input v_1107;
input v_1108;
input v_1109;
input v_1110;
input v_1111;
input v_1112;
input v_1113;
input v_1114;
input v_1115;
input v_1116;
input v_1117;
input v_1118;
input v_1119;
input v_1120;
input v_1121;
input v_1122;
input v_1123;
input v_1124;
input v_1125;
input v_1126;
input v_1127;
input v_1128;
input v_1129;
input v_1130;
input v_1131;
input v_1132;
input v_1133;
input v_1134;
input v_1135;
input v_1136;
input v_1137;
input v_1138;
input v_1139;
input v_1140;
input v_1141;
input v_1142;
input v_1143;
input v_1144;
input v_1145;
input v_1146;
input v_1147;
input v_1148;
input v_1149;
input v_1150;
input v_1151;
input v_1152;
input v_1153;
input v_1154;
input v_1155;
input v_1156;
input v_1157;
input v_1158;
input v_1159;
input v_1160;
input v_1161;
input v_1162;
input v_1163;
input v_1164;
input v_1165;
input v_1166;
input v_1167;
input v_1168;
input v_1169;
input v_1170;
input v_1171;
input v_1172;
input v_1173;
input v_1174;
input v_1175;
input v_1176;
input v_1177;
input v_1178;
input v_1179;
input v_1180;
input v_1181;
input v_1182;
input v_1183;
input v_1184;
input v_1185;
input v_1186;
input v_1187;
input v_1188;
input v_1189;
input v_1190;
input v_1191;
input v_1192;
input v_1193;
input v_1194;
input v_1195;
input v_1196;
input v_1197;
input v_1198;
input v_1199;
input v_1200;
input v_1201;
input v_1202;
input v_1203;
input v_1204;
input v_1205;
input v_1206;
input v_1207;
input v_1208;
input v_1209;
input v_1210;
input v_1211;
input v_1212;
input v_1213;
input v_1214;
input v_1215;
input v_1216;
input v_1217;
input v_1218;
input v_1219;
input v_1220;
input v_1221;
input v_1222;
input v_1223;
input v_1224;
input v_1225;
input v_1226;
input v_1227;
input v_1228;
input v_1229;
input v_1230;
input v_1231;
input v_1232;
input v_1233;
input v_1234;
input v_1235;
input v_1236;
input v_1237;
input v_1238;
input v_1239;
input v_1240;
input v_1241;
input v_1242;
input v_1243;
input v_1244;
input v_1245;
input v_1246;
input v_1247;
input v_1248;
input v_1249;
input v_1250;
input v_1251;
input v_1252;
input v_1253;
input v_1254;
input v_1255;
input v_1256;
input v_1257;
input v_1258;
input v_1259;
input v_1260;
input v_1261;
input v_1262;
input v_1263;
input v_1264;
input v_1265;
input v_1266;
input v_1267;
input v_1268;
input v_1269;
input v_1270;
input v_1271;
input v_1272;
input v_1273;
input v_1274;
input v_1275;
input v_1276;
input v_1277;
input v_1278;
input v_1279;
input v_1280;
input v_1281;
input v_1282;
input v_1283;
input v_1284;
input v_1285;
input v_1286;
input v_1287;
input v_1288;
input v_1289;
input v_1290;
input v_1291;
input v_1292;
input v_1293;
input v_1294;
input v_1295;
input v_1296;
input v_1297;
input v_1298;
input v_1299;
input v_1300;
input v_1301;
input v_1302;
input v_1303;
input v_1304;
input v_1305;
input v_1306;
input v_1307;
input v_1308;
input v_1309;
input v_1310;
input v_1311;
input v_1312;
input v_1313;
input v_1314;
input v_1315;
input v_1316;
input v_1317;
input v_1318;
input v_1319;
input v_1320;
input v_1321;
input v_1322;
input v_1323;
input v_1324;
input v_1325;
input v_1326;
input v_1327;
input v_1328;
input v_1329;
input v_1330;
input v_1331;
input v_1332;
input v_1333;
input v_1334;
input v_1335;
input v_1336;
input v_1337;
input v_1338;
input v_1339;
input v_1340;
input v_1341;
input v_1342;
input v_1343;
input v_1344;
input v_1345;
input v_1346;
input v_1347;
input v_1348;
input v_1349;
input v_1350;
input v_1351;
input v_1352;
input v_1353;
input v_1354;
input v_1355;
input v_1356;
input v_1357;
input v_1358;
input v_1359;
input v_1360;
input v_1361;
input v_1362;
input v_1363;
input v_1364;
input v_1365;
input v_1366;
input v_1367;
input v_1368;
input v_1369;
input v_1370;
input v_1371;
input v_1372;
input v_1373;
input v_1374;
input v_1375;
input v_1376;
input v_1377;
input v_1378;
input v_1379;
input v_1380;
input v_1381;
input v_1382;
input v_1383;
input v_1384;
input v_1385;
input v_1386;
input v_1387;
input v_1388;
input v_1389;
input v_1390;
input v_1391;
input v_1392;
input v_1393;
input v_1394;
input v_1395;
input v_1396;
input v_1397;
input v_1398;
input v_1399;
input v_1400;
input v_1401;
input v_1402;
input v_1403;
input v_1404;
input v_1405;
input v_1406;
input v_1407;
input v_1408;
input v_1409;
input v_1410;
input v_1411;
input v_1412;
input v_1413;
input v_1414;
input v_1415;
input v_1416;
input v_1417;
input v_1418;
input v_1419;
input v_1420;
input v_1421;
input v_1422;
input v_1423;
input v_1424;
input v_1425;
input v_1426;
input v_1427;
input v_1428;
input v_1429;
input v_1430;
input v_1431;
input v_1432;
input v_1433;
input v_1434;
input v_1435;
input v_1436;
input v_1437;
input v_1438;
input v_1439;
input v_1440;
input v_1441;
input v_1442;
input v_1443;
input v_1444;
input v_1445;
input v_1446;
input v_1447;
input v_1448;
input v_1449;
input v_1450;
input v_1451;
input v_1452;
input v_1453;
input v_1454;
input v_1455;
input v_1456;
input v_1457;
input v_1458;
input v_1459;
input v_1460;
input v_1461;
input v_1462;
input v_1463;
input v_1464;
input v_1465;
input v_1466;
input v_1467;
input v_1468;
input v_1469;
input v_1470;
input v_1471;
input v_1472;
input v_1473;
input v_1474;
input v_1475;
input v_1476;
input v_1477;
input v_1478;
input v_1479;
input v_1480;
input v_1481;
input v_1482;
input v_1483;
input v_1484;
input v_1485;
input v_1486;
input v_1487;
input v_1488;
input v_1489;
input v_1490;
input v_1491;
input v_1492;
input v_1493;
input v_1494;
input v_1495;
input v_1496;
input v_1497;
input v_1498;
input v_1499;
input v_1500;
input v_1501;
input v_1502;
input v_1503;
input v_1504;
input v_1505;
input v_1506;
input v_1507;
input v_1508;
input v_1509;
input v_1510;
input v_1511;
input v_1512;
input v_1513;
input v_1514;
input v_1515;
input v_1516;
input v_1517;
input v_1518;
input v_1519;
input v_1520;
input v_1521;
input v_1522;
input v_1523;
input v_1524;
input v_1525;
input v_1526;
input v_1527;
input v_1528;
input v_1529;
input v_1530;
input v_1531;
input v_1532;
input v_1533;
input v_1534;
input v_1535;
input v_1536;
input v_1537;
input v_1538;
input v_1539;
input v_1540;
input v_1541;
input v_1542;
input v_1543;
input v_1544;
input v_1545;
input v_1546;
input v_1547;
input v_1548;
input v_1549;
input v_1550;
input v_1551;
input v_1552;
input v_1553;
input v_1554;
input v_1555;
input v_1556;
input v_1557;
input v_1558;
input v_1559;
input v_1560;
input v_1561;
input v_1562;
input v_1563;
input v_1564;
input v_1565;
input v_1566;
input v_1567;
input v_1568;
input v_1569;
input v_1570;
input v_1571;
input v_1572;
input v_1573;
input v_1574;
input v_1575;
input v_1576;
input v_1577;
input v_1578;
input v_1579;
input v_1580;
input v_1581;
input v_1582;
input v_1583;
input v_1584;
input v_1585;
input v_1586;
input v_1587;
input v_1588;
input v_1589;
input v_1590;
input v_1591;
input v_1592;
input v_1593;
input v_1594;
input v_1595;
input v_1596;
input v_1597;
input v_1598;
input v_1599;
input v_1600;
input v_1601;
input v_1602;
input v_1603;
input v_1604;
input v_1605;
input v_1606;
input v_1607;
input v_1608;
input v_1609;
input v_1610;
input v_1611;
input v_1612;
input v_1613;
input v_1614;
input v_1615;
input v_1616;
input v_1617;
input v_1618;
input v_1619;
input v_1620;
input v_1621;
input v_1622;
input v_1623;
input v_1624;
input v_1625;
input v_1626;
input v_1627;
input v_1628;
input v_1629;
input v_1630;
input v_1631;
input v_1632;
input v_1633;
input v_1634;
input v_1635;
input v_1636;
input v_1637;
input v_1638;
input v_1639;
input v_1640;
input v_1641;
input v_1642;
input v_1643;
input v_1644;
input v_1645;
input v_1646;
input v_1647;
input v_1648;
input v_1649;
input v_1650;
input v_1651;
input v_1652;
input v_1653;
input v_1654;
input v_1655;
input v_1656;
input v_1657;
input v_1658;
input v_1659;
input v_1660;
input v_1661;
input v_1662;
input v_1663;
input v_1664;
input v_1665;
input v_1666;
input v_1667;
input v_1668;
input v_1669;
input v_1670;
input v_1671;
input v_1672;
input v_1673;
input v_1674;
input v_1675;
input v_1676;
input v_1677;
input v_1678;
input v_1679;
input v_1680;
input v_1681;
input v_1682;
input v_1683;
input v_1684;
input v_1685;
input v_1686;
input v_1687;
input v_1688;
input v_1689;
input v_1690;
input v_1691;
input v_1692;
input v_1693;
input v_1694;
input v_1695;
input v_1696;
input v_1697;
input v_1698;
input v_1699;
input v_1700;
input v_1701;
input v_1702;
input v_1703;
input v_1704;
input v_1705;
input v_1706;
input v_1707;
input v_1708;
input v_1709;
input v_1710;
input v_1711;
input v_1712;
input v_1713;
input v_1714;
input v_1715;
input v_1716;
input v_1717;
input v_1718;
input v_1719;
input v_1720;
input v_1721;
input v_1722;
input v_1723;
input v_1724;
input v_1725;
input v_1726;
input v_1727;
input v_1728;
input v_1729;
input v_1730;
input v_1731;
input v_1732;
input v_1733;
input v_1734;
input v_1735;
input v_1736;
input v_1737;
input v_1738;
input v_1739;
input v_1740;
input v_1741;
input v_1742;
input v_1743;
input v_1744;
input v_1745;
input v_1746;
input v_1747;
input v_1748;
input v_1749;
input v_1750;
input v_1751;
input v_1752;
input v_1753;
input v_1754;
input v_1755;
input v_1756;
input v_1757;
input v_1758;
input v_1759;
input v_1760;
input v_1761;
input v_1762;
input v_1763;
input v_1764;
input v_1765;
input v_1766;
input v_1767;
input v_1768;
input v_1769;
input v_1770;
input v_1771;
input v_1772;
input v_1773;
input v_1774;
input v_1775;
input v_1776;
input v_1777;
input v_1778;
input v_1779;
input v_1780;
input v_1781;
input v_1782;
input v_1783;
input v_1784;
input v_1785;
input v_1786;
input v_1787;
input v_1788;
input v_1789;
input v_1790;
input v_1791;
input v_1792;
input v_1793;
input v_1794;
input v_1795;
input v_1796;
input v_1797;
input v_1798;
input v_1799;
input v_1800;
input v_1801;
input v_1802;
input v_1803;
input v_1804;
input v_1805;
input v_1806;
input v_1807;
input v_1808;
input v_1809;
input v_1810;
input v_1811;
input v_1812;
input v_1813;
input v_1814;
input v_1815;
input v_1816;
input v_1817;
input v_1818;
input v_1819;
input v_1820;
input v_1821;
input v_1822;
input v_1823;
input v_1824;
input v_1825;
input v_1826;
input v_1827;
input v_1828;
input v_1829;
input v_1830;
input v_1831;
input v_1832;
input v_1833;
input v_1834;
input v_1835;
input v_1836;
input v_1837;
input v_1838;
input v_1839;
input v_1840;
input v_1841;
input v_1842;
input v_1843;
input v_1844;
input v_1845;
input v_1846;
input v_1847;
input v_1848;
input v_1849;
input v_1850;
input v_1851;
input v_1852;
input v_1853;
input v_1854;
input v_1855;
input v_1856;
input v_1857;
input v_1858;
input v_1859;
input v_1860;
input v_1861;
input v_1862;
input v_1863;
input v_1864;
input v_1865;
input v_1866;
input v_1867;
input v_1868;
input v_1869;
input v_1870;
input v_1871;
input v_1872;
input v_1873;
input v_1874;
input v_1875;
input v_1876;
input v_1877;
input v_1878;
input v_1879;
input v_1880;
input v_1881;
input v_1882;
input v_1883;
input v_1884;
input v_1885;
input v_1886;
input v_1887;
input v_1888;
input v_1889;
input v_1890;
input v_1891;
input v_1892;
input v_1893;
input v_1894;
input v_1895;
input v_1896;
input v_1897;
input v_1898;
input v_1899;
input v_1900;
input v_1901;
input v_1902;
input v_1903;
input v_1904;
input v_1905;
input v_1906;
input v_1907;
input v_1908;
input v_1909;
input v_1910;
input v_1911;
input v_1912;
input v_1913;
input v_1914;
input v_1915;
input v_1916;
input v_1917;
input v_1918;
input v_1919;
input v_1920;
input v_1921;
input v_1922;
input v_1923;
input v_1924;
input v_1925;
input v_1926;
input v_1927;
input v_1928;
input v_1929;
input v_1930;
input v_1931;
input v_1932;
input v_1933;
input v_1934;
input v_1935;
input v_1936;
input v_1937;
input v_1938;
input v_1939;
input v_1940;
input v_1941;
input v_1942;
input v_1943;
input v_1944;
input v_1945;
input v_1946;
input v_1947;
input v_1948;
input v_1949;
input v_1950;
input v_1951;
input v_1952;
input v_1953;
input v_1954;
input v_1955;
input v_1956;
input v_1957;
input v_1958;
input v_1959;
input v_1960;
input v_1961;
input v_1962;
input v_1963;
input v_1964;
input v_1965;
input v_1966;
input v_1967;
input v_1968;
input v_1969;
input v_1970;
input v_1971;
input v_1972;
input v_1973;
input v_1974;
input v_1975;
input v_1976;
input v_1977;
input v_1978;
input v_1979;
input v_1980;
input v_1981;
input v_1982;
input v_1983;
input v_1984;
input v_1985;
input v_1986;
input v_1987;
input v_1988;
input v_1989;
input v_1990;
input v_1991;
input v_1992;
input v_1993;
input v_1994;
input v_1995;
input v_1996;
input v_1997;
input v_1998;
input v_1999;
input v_2000;
input v_2001;
input v_2002;
input v_2003;
input v_2004;
input v_2005;
input v_2006;
input v_2007;
input v_2008;
input v_2009;
input v_2010;
input v_2011;
input v_2012;
input v_2013;
input v_2014;
input v_2015;
input v_2016;
input v_2017;
input v_2018;
input v_2019;
input v_2020;
input v_2021;
input v_2022;
input v_2023;
input v_2024;
input v_2025;
input v_2026;
input v_2027;
input v_2028;
input v_2029;
input v_2030;
input v_2031;
input v_2032;
input v_2033;
input v_2034;
input v_2035;
input v_2036;
input v_2037;
input v_2038;
input v_2039;
input v_2040;
input v_2041;
input v_2042;
input v_2043;
input v_2044;
input v_2045;
input v_2046;
input v_2047;
input v_2048;
input v_2049;
input v_2050;
input v_2051;
input v_2052;
input v_2053;
input v_2054;
input v_2055;
input v_2056;
input v_2057;
input v_2058;
input v_2059;
input v_2060;
input v_2061;
input v_2062;
input v_2063;
input v_2064;
input v_2065;
input v_2066;
input v_2067;
input v_2068;
input v_2069;
input v_2070;
input v_2071;
input v_2072;
input v_2073;
input v_2074;
input v_2075;
input v_2076;
input v_2077;
input v_2078;
input v_2079;
input v_2080;
input v_2081;
input v_2082;
input v_2083;
input v_2084;
input v_2085;
input v_2086;
input v_2087;
input v_2088;
input v_2089;
input v_2090;
input v_2091;
input v_2092;
input v_2093;
input v_2094;
input v_2095;
input v_2096;
input v_2097;
input v_2098;
input v_2099;
input v_2100;
input v_2101;
input v_2102;
input v_2103;
input v_2104;
input v_2105;
input v_2106;
input v_2107;
input v_2108;
input v_2109;
input v_2110;
input v_2111;
input v_2112;
input v_2113;
input v_2114;
input v_2115;
input v_2116;
input v_2117;
input v_2118;
input v_2119;
input v_2120;
input v_2121;
input v_2122;
input v_2123;
input v_2124;
input v_2125;
input v_2126;
input v_2127;
input v_2128;
input v_2129;
input v_2130;
input v_2131;
input v_2132;
input v_2133;
input v_2134;
input v_2135;
input v_2136;
input v_2137;
input v_2138;
input v_2139;
input v_2140;
input v_2141;
input v_2142;
input v_2143;
input v_2144;
input v_2145;
input v_2146;
input v_2147;
input v_2148;
input v_2149;
input v_2150;
input v_2151;
input v_2152;
input v_2153;
input v_2154;
input v_2155;
input v_2156;
input v_2157;
input v_2158;
input v_2159;
input v_2160;
input v_2161;
input v_2162;
input v_2163;
input v_2164;
input v_2165;
input v_2166;
input v_2167;
input v_2168;
input v_2169;
input v_2170;
input v_2171;
input v_2172;
input v_2173;
input v_2174;
input v_2175;
input v_2176;
input v_2177;
input v_2178;
input v_2179;
input v_2180;
input v_2181;
input v_2182;
input v_2183;
input v_2184;
input v_2185;
input v_2186;
input v_2187;
input v_2188;
input v_2189;
input v_2190;
input v_2191;
input v_2192;
input v_2193;
input v_2194;
input v_2195;
input v_2196;
input v_2197;
input v_2198;
input v_2199;
input v_2200;
input v_2201;
input v_2202;
input v_2203;
input v_2204;
input v_2205;
input v_2206;
input v_2207;
input v_2208;
input v_2209;
input v_2210;
input v_2211;
input v_2212;
input v_2213;
input v_2214;
input v_2215;
input v_2216;
input v_2217;
input v_2218;
input v_2219;
input v_2220;
input v_2221;
input v_2222;
input v_2223;
input v_2224;
input v_2225;
input v_2226;
input v_2227;
input v_2228;
input v_2229;
input v_2230;
input v_2231;
input v_2232;
input v_2233;
input v_2234;
input v_2235;
input v_2236;
input v_2237;
input v_2238;
input v_2239;
input v_2240;
input v_2241;
input v_2242;
input v_2243;
input v_2244;
input v_2245;
input v_2246;
input v_2247;
input v_2248;
input v_2249;
input v_2250;
input v_2251;
input v_2252;
input v_2253;
input v_2254;
input v_2255;
input v_2256;
input v_2257;
input v_2258;
input v_2259;
input v_2260;
input v_2261;
input v_2262;
input v_2263;
input v_2264;
input v_2265;
input v_2266;
input v_2267;
input v_2268;
input v_2269;
input v_2270;
input v_2271;
input v_2272;
input v_2273;
input v_2274;
input v_2275;
input v_2276;
input v_2277;
input v_2278;
input v_2279;
input v_2280;
input v_2281;
input v_2282;
input v_2283;
input v_2284;
input v_2285;
input v_2286;
input v_2287;
input v_2288;
input v_2289;
input v_2290;
input v_2291;
input v_2292;
input v_2293;
input v_2294;
input v_2295;
input v_2296;
input v_2297;
input v_2298;
input v_2299;
input v_2300;
input v_2301;
input v_2302;
input v_2303;
input v_2304;
input v_2305;
input v_2306;
input v_2307;
input v_2308;
input v_2309;
input v_2310;
input v_2311;
input v_2312;
input v_2313;
input v_2314;
input v_2315;
input v_2316;
input v_2317;
input v_2318;
input v_2319;
input v_2320;
input v_2321;
input v_2322;
input v_2323;
input v_2324;
input v_2325;
input v_2326;
input v_2327;
input v_2328;
input v_2329;
input v_2330;
input v_2331;
input v_2332;
input v_2333;
input v_2334;
input v_2335;
input v_2336;
input v_2337;
input v_2338;
input v_2339;
input v_2340;
input v_2341;
input v_2342;
input v_2343;
input v_2344;
input v_2345;
input v_2346;
input v_2347;
input v_2348;
input v_2349;
input v_2350;
input v_2351;
input v_2352;
input v_2353;
input v_2354;
input v_2355;
input v_2356;
input v_2357;
input v_2358;
input v_2359;
input v_2360;
input v_2361;
input v_2362;
input v_2363;
input v_2364;
input v_2365;
input v_2366;
input v_2367;
input v_2368;
input v_2369;
input v_2370;
input v_2371;
input v_2372;
input v_2373;
input v_2374;
input v_2375;
input v_2376;
input v_2377;
input v_2378;
input v_2379;
input v_2380;
input v_2381;
input v_2382;
input v_2383;
input v_2384;
input v_2385;
input v_2386;
input v_2387;
input v_2388;
input v_2389;
input v_2390;
input v_2391;
input v_2392;
input v_2393;
input v_2394;
input v_2395;
input v_2396;
input v_2397;
input v_2398;
input v_2399;
input v_2400;
input v_2401;
input v_2402;
input v_2403;
input v_2404;
input v_2405;
input v_2406;
input v_2407;
input v_2408;
input v_2409;
input v_2410;
input v_2411;
input v_2412;
input v_2413;
input v_2414;
input v_2415;
input v_2416;
input v_2417;
input v_2418;
input v_2419;
input v_2420;
input v_2421;
input v_2422;
input v_2423;
input v_2424;
input v_2425;
input v_2426;
input v_2427;
input v_2428;
input v_2429;
input v_2430;
input v_2431;
input v_2432;
input v_2433;
input v_2434;
input v_2435;
input v_2436;
input v_2437;
input v_2438;
input v_2439;
input v_2440;
input v_2441;
input v_2442;
input v_2443;
input v_2444;
input v_2445;
input v_2446;
input v_2447;
input v_2448;
input v_2449;
input v_2450;
input v_2451;
input v_2452;
input v_2453;
input v_2454;
input v_2455;
input v_2456;
input v_2457;
input v_2458;
input v_2459;
input v_2460;
input v_2461;
input v_2462;
input v_2463;
input v_2464;
input v_2465;
input v_2466;
input v_2467;
input v_2468;
input v_2469;
input v_2470;
input v_2471;
input v_2472;
input v_2473;
input v_2474;
input v_2475;
input v_2476;
input v_2477;
input v_2478;
input v_2479;
input v_2480;
input v_2481;
input v_2482;
input v_2483;
input v_2484;
input v_2485;
input v_2486;
input v_2487;
input v_2488;
input v_2489;
input v_2490;
input v_2491;
input v_2492;
input v_2493;
input v_2494;
input v_2495;
input v_2496;
input v_2497;
input v_2498;
input v_2499;
input v_2500;
input v_2501;
input v_2502;
input v_2503;
input v_2504;
input v_2505;
input v_2506;
input v_2507;
input v_2508;
input v_2509;
input v_2510;
input v_2511;
input v_2512;
input v_2513;
input v_2514;
input v_2515;
input v_2516;
input v_2517;
input v_2518;
input v_2519;
input v_2520;
input v_2521;
input v_2522;
input v_2523;
input v_2524;
input v_2525;
input v_2526;
input v_2527;
input v_2528;
input v_2529;
input v_2530;
input v_2531;
input v_2532;
input v_2533;
input v_2534;
input v_2535;
input v_2536;
input v_2537;
input v_2538;
input v_2539;
input v_2540;
input v_2541;
input v_2542;
input v_2543;
input v_2544;
input v_2545;
input v_2546;
input v_2547;
input v_2548;
input v_2549;
input v_2550;
input v_2551;
input v_2552;
input v_2553;
input v_2554;
input v_2555;
input v_2556;
input v_2557;
input v_2558;
input v_2559;
input v_2560;
input v_2561;
input v_2562;
input v_2563;
input v_2564;
input v_2565;
input v_2566;
input v_2567;
input v_2568;
input v_2569;
input v_2570;
input v_2571;
input v_2572;
input v_2573;
input v_2574;
input v_2575;
input v_2576;
input v_2577;
input v_2578;
input v_2579;
input v_2580;
input v_2581;
input v_2582;
input v_2583;
input v_2584;
input v_2585;
input v_2586;
input v_2587;
input v_2588;
input v_2589;
input v_2590;
input v_2591;
input v_2592;
input v_2593;
input v_2594;
input v_2595;
input v_2596;
input v_2597;
input v_2598;
input v_2599;
input v_2600;
input v_2601;
input v_2602;
input v_2603;
input v_2604;
input v_2605;
input v_2606;
input v_2607;
input v_2608;
input v_2609;
input v_2610;
input v_2611;
input v_2612;
input v_2613;
input v_2614;
input v_2615;
input v_2616;
input v_2617;
input v_2618;
input v_2619;
input v_2620;
input v_2621;
input v_2622;
input v_2623;
input v_2624;
input v_2625;
input v_2626;
input v_2627;
input v_2628;
input v_2629;
input v_2630;
input v_2631;
input v_2632;
input v_2633;
input v_2634;
input v_2635;
input v_2636;
input v_2637;
input v_2638;
input v_2639;
input v_2640;
input v_2641;
input v_2642;
input v_2643;
input v_2644;
input v_2645;
input v_2646;
input v_2647;
input v_2648;
input v_2649;
input v_2650;
input v_2651;
input v_2652;
input v_2653;
input v_2654;
input v_2655;
input v_2656;
input v_2657;
input v_2658;
input v_2659;
input v_2660;
input v_2661;
input v_2662;
input v_2663;
input v_2664;
input v_2665;
input v_2666;
input v_2667;
input v_2668;
input v_2669;
input v_2670;
input v_2671;
input v_2672;
input v_2673;
input v_2674;
input v_2675;
input v_2676;
input v_2677;
input v_2678;
input v_2679;
input v_2680;
input v_2681;
input v_2682;
input v_2683;
input v_2684;
input v_2685;
input v_2686;
input v_2687;
input v_2688;
input v_2689;
input v_2690;
input v_2691;
input v_2692;
input v_2693;
input v_2694;
input v_2695;
input v_2696;
input v_2697;
input v_2698;
input v_2699;
input v_2700;
input v_2701;
input v_2702;
input v_2703;
input v_2704;
input v_2705;
input v_2706;
input v_2707;
input v_2708;
input v_2709;
input v_2710;
input v_2711;
input v_2712;
input v_2713;
input v_2714;
input v_2715;
input v_2716;
input v_2717;
input v_2718;
input v_2719;
input v_2720;
input v_2721;
input v_2722;
input v_2723;
input v_2724;
input v_2725;
input v_2726;
input v_2727;
input v_2728;
input v_2729;
input v_2730;
input v_2731;
input v_2732;
input v_2733;
input v_2734;
input v_2735;
input v_2736;
input v_2737;
input v_2738;
input v_2739;
input v_2740;
input v_2741;
input v_2742;
input v_2743;
input v_2744;
input v_2745;
input v_2746;
input v_2747;
input v_2748;
input v_2749;
input v_2750;
input v_2751;
input v_2752;
input v_2753;
input v_2754;
input v_2755;
input v_2756;
input v_2757;
input v_2758;
input v_2759;
input v_2760;
input v_2761;
input v_2762;
input v_2763;
input v_2764;
input v_2765;
input v_2766;
input v_2767;
input v_2768;
input v_2769;
input v_2770;
input v_2771;
input v_2772;
input v_2773;
input v_2774;
input v_2775;
input v_2776;
input v_2777;
input v_2778;
input v_2779;
input v_2780;
input v_2781;
input v_2782;
input v_2783;
input v_2784;
input v_2785;
input v_2786;
input v_2787;
input v_2788;
input v_2789;
input v_2790;
input v_2791;
input v_2792;
input v_2793;
input v_2794;
input v_2795;
input v_2796;
input v_2797;
input v_2798;
input v_2799;
input v_2800;
input v_2801;
input v_2802;
input v_2803;
input v_2804;
input v_2805;
input v_2806;
input v_2807;
input v_2808;
input v_2809;
input v_2810;
input v_2811;
input v_2812;
input v_2813;
input v_2814;
input v_2815;
input v_2816;
input v_2817;
input v_2818;
input v_2819;
input v_2820;
input v_2821;
input v_2822;
input v_2823;
input v_2824;
input v_2825;
input v_2826;
input v_2827;
input v_2828;
input v_2829;
input v_2830;
input v_2831;
input v_2832;
input v_2833;
input v_2834;
input v_2835;
input v_2836;
input v_2837;
input v_2838;
input v_2839;
input v_2840;
input v_2841;
input v_2842;
input v_2843;
input v_2844;
input v_2845;
input v_2846;
input v_2847;
input v_2848;
input v_2849;
input v_2850;
input v_2851;
input v_2852;
input v_2853;
input v_2854;
input v_2855;
input v_2856;
input v_2857;
input v_2858;
input v_2859;
input v_2860;
input v_2861;
input v_2862;
input v_2863;
input v_2864;
input v_2865;
input v_2866;
input v_2867;
input v_2868;
input v_2869;
input v_2870;
input v_2871;
input v_2872;
input v_2873;
input v_2874;
input v_2875;
input v_2876;
input v_2877;
input v_2878;
input v_2879;
input v_2880;
input v_2881;
input v_2882;
input v_2883;
input v_2884;
input v_2885;
input v_2886;
input v_2887;
input v_2888;
input v_2889;
input v_2890;
input v_2891;
input v_2892;
input v_2893;
input v_2894;
input v_2895;
input v_2896;
input v_2897;
input v_2898;
input v_2899;
input v_2900;
input v_2901;
input v_2902;
input v_2903;
input v_2904;
input v_2905;
input v_2906;
input v_2907;
input v_2908;
input v_2909;
input v_2910;
input v_2911;
input v_2912;
input v_2913;
input v_2914;
input v_2915;
input v_2916;
input v_2917;
input v_2918;
input v_2919;
input v_2920;
input v_2921;
input v_2922;
input v_2923;
input v_2924;
input v_2925;
input v_2926;
input v_2927;
input v_2928;
input v_2929;
input v_2930;
input v_2931;
input v_2932;
input v_2933;
input v_2934;
input v_2935;
input v_2936;
input v_2937;
input v_2938;
input v_2939;
input v_2940;
input v_2941;
input v_2942;
input v_2943;
input v_2944;
input v_2945;
input v_2946;
input v_2947;
input v_2948;
input v_2949;
input v_2950;
input v_2951;
input v_2952;
input v_2953;
input v_2954;
input v_2955;
input v_2956;
input v_2957;
input v_2958;
input v_2959;
input v_2960;
input v_2961;
input v_2962;
input v_2963;
input v_2964;
input v_2965;
input v_2966;
input v_2967;
input v_2968;
input v_2969;
input v_2970;
input v_2971;
input v_2972;
input v_2973;
input v_2974;
input v_2975;
input v_2976;
input v_2977;
input v_2978;
input v_2979;
input v_2980;
input v_2981;
input v_2982;
input v_2983;
input v_2984;
input v_2985;
input v_2986;
input v_2987;
input v_2988;
input v_2989;
input v_2990;
input v_2991;
input v_2992;
input v_2993;
input v_2994;
input v_2995;
input v_2996;
input v_2997;
input v_2998;
input v_2999;
input v_3000;
input v_3001;
input v_3002;
input v_3003;
input v_3004;
input v_3005;
input v_3006;
input v_3007;
input v_3008;
input v_3009;
input v_3010;
input v_3011;
input v_3012;
input v_3013;
input v_3014;
input v_3015;
input v_3016;
input v_3017;
input v_3018;
input v_3019;
input v_3020;
input v_3021;
input v_3022;
input v_3023;
input v_3024;
input v_3025;
input v_3026;
input v_3027;
input v_3028;
input v_3029;
input v_3030;
input v_3031;
input v_3032;
input v_3033;
input v_3034;
input v_3035;
input v_3036;
input v_3037;
input v_3038;
input v_3039;
input v_3040;
input v_3041;
input v_3042;
input v_3043;
input v_3044;
input v_3045;
input v_3046;
input v_3047;
input v_3048;
input v_3049;
input v_3050;
input v_3051;
input v_3052;
input v_3053;
input v_3054;
input v_3055;
input v_3056;
input v_3057;
input v_3058;
input v_3059;
input v_3060;
input v_3061;
input v_3062;
input v_3063;
input v_3064;
input v_3065;
input v_3066;
input v_3067;
input v_3068;
input v_3069;
input v_3070;
input v_3071;
input v_3072;
input v_3073;
input v_3074;
input v_3075;
input v_3076;
input v_3077;
input v_3078;
input v_3079;
input v_3080;
input v_3081;
input v_3082;
input v_3083;
input v_3084;
input v_3085;
input v_3086;
input v_3087;
input v_3088;
input v_3089;
input v_3090;
input v_3091;
input v_3092;
input v_3093;
input v_3094;
input v_3095;
input v_3096;
input v_3097;
input v_3098;
input v_3099;
input v_3100;
input v_3101;
input v_3102;
input v_3103;
input v_3104;
input v_3105;
input v_3106;
input v_3107;
input v_3108;
input v_3109;
input v_3110;
input v_3111;
input v_3112;
input v_3113;
input v_3114;
input v_3115;
input v_3116;
input v_3117;
input v_3118;
input v_3119;
input v_3120;
input v_3121;
input v_3122;
input v_3123;
input v_3124;
input v_3125;
input v_3126;
input v_3127;
input v_3128;
input v_3129;
input v_3130;
input v_3131;
input v_3132;
input v_3133;
input v_3134;
input v_3135;
input v_3136;
input v_3137;
input v_3138;
input v_3139;
input v_3140;
input v_3141;
input v_3142;
input v_3143;
input v_3144;
input v_3145;
input v_3146;
input v_3147;
input v_3148;
input v_3149;
input v_3150;
input v_3151;
input v_3152;
input v_3153;
input v_3154;
input v_3155;
input v_3156;
input v_3157;
input v_3158;
input v_3159;
input v_3160;
input v_3161;
input v_3162;
input v_3163;
input v_3164;
input v_3165;
input v_3166;
input v_3167;
input v_3168;
input v_3169;
input v_3170;
input v_3171;
input v_3172;
input v_3173;
input v_3174;
input v_3175;
input v_3176;
input v_3177;
input v_3178;
input v_3179;
input v_3180;
input v_3181;
input v_3182;
input v_3183;
input v_3184;
input v_3185;
input v_3186;
input v_3187;
input v_3188;
input v_3189;
input v_3190;
input v_3191;
input v_3192;
input v_3193;
input v_3194;
input v_3195;
input v_3196;
input v_3197;
input v_3198;
input v_3199;
input v_3200;
input v_3201;
input v_3202;
input v_3203;
input v_3204;
input v_3205;
input v_3206;
input v_3207;
input v_3208;
input v_3209;
input v_3210;
input v_3211;
input v_3212;
input v_3213;
input v_3214;
input v_3215;
input v_3216;
input v_3217;
input v_3218;
input v_3219;
input v_3220;
input v_3221;
input v_3222;
input v_3223;
input v_3224;
input v_3225;
input v_3226;
input v_3227;
input v_3228;
input v_3229;
input v_3230;
input v_3231;
input v_3232;
input v_3233;
input v_3234;
input v_3235;
input v_3236;
input v_3237;
input v_3238;
input v_3239;
input v_3240;
input v_3241;
input v_3242;
input v_3243;
input v_3244;
input v_3245;
input v_3246;
input v_3247;
input v_3248;
input v_3249;
input v_3250;
input v_3251;
input v_3252;
input v_3253;
input v_3254;
input v_3255;
input v_3256;
input v_3257;
input v_3258;
input v_3259;
input v_3260;
input v_3261;
input v_3262;
input v_3263;
input v_3264;
input v_3265;
input v_3266;
input v_3267;
input v_3268;
input v_3269;
input v_3270;
input v_3271;
input v_3272;
input v_3273;
input v_3274;
input v_3275;
input v_3276;
input v_3277;
input v_3278;
input v_3279;
input v_3280;
input v_3281;
input v_3282;
input v_3283;
input v_3284;
input v_3285;
input v_3286;
input v_3287;
input v_3288;
input v_3289;
input v_3290;
input v_3291;
input v_3292;
input v_3293;
input v_3294;
input v_3295;
input v_3296;
input v_3297;
input v_3298;
input v_3299;
input v_3300;
input v_3301;
input v_3302;
input v_3303;
input v_3304;
input v_3305;
input v_3306;
input v_3307;
input v_3308;
input v_3309;
input v_3310;
input v_3311;
input v_3312;
input v_3313;
input v_3314;
input v_3315;
input v_3316;
input v_3317;
input v_3318;
input v_3319;
input v_3320;
input v_3321;
input v_3322;
input v_3323;
input v_3324;
input v_3325;
input v_3326;
input v_3327;
input v_3328;
input v_3329;
input v_3330;
input v_3331;
input v_3332;
input v_3333;
input v_3334;
input v_3335;
input v_3336;
input v_3337;
input v_3338;
input v_3339;
input v_3340;
input v_3341;
input v_3342;
input v_3343;
input v_3344;
input v_3345;
input v_3346;
input v_3347;
input v_3348;
input v_3349;
input v_3350;
input v_3351;
input v_3352;
input v_3353;
input v_3354;
input v_3355;
input v_3356;
input v_3357;
input v_3358;
input v_3359;
input v_3360;
input v_3361;
input v_3362;
input v_3363;
input v_3364;
input v_3365;
input v_3366;
input v_3367;
input v_3368;
input v_3369;
input v_3370;
input v_3371;
input v_3372;
input v_3373;
input v_3374;
input v_3375;
input v_3376;
input v_3377;
input v_3378;
input v_3379;
input v_3380;
input v_3381;
input v_3382;
input v_3383;
input v_3384;
input v_3385;
input v_3386;
input v_3387;
input v_3388;
input v_3389;
input v_3390;
input v_3391;
input v_3392;
input v_3393;
input v_3394;
input v_3395;
input v_3396;
input v_3397;
input v_3398;
input v_3399;
input v_3400;
input v_3401;
input v_3402;
input v_3403;
input v_3404;
input v_3405;
input v_3406;
input v_3407;
input v_3408;
input v_3409;
input v_3410;
input v_3411;
input v_3412;
input v_3413;
input v_3414;
input v_3415;
input v_3416;
input v_3417;
input v_3418;
input v_3419;
input v_3420;
input v_3421;
input v_3422;
input v_3423;
input v_3424;
input v_3425;
input v_3426;
input v_3427;
input v_3428;
input v_3429;
input v_3430;
input v_3431;
input v_3432;
input v_3433;
input v_3434;
input v_3435;
input v_3436;
input v_3437;
input v_3438;
input v_3439;
input v_3440;
input v_3441;
input v_3442;
input v_3443;
input v_3444;
input v_3445;
input v_3446;
input v_3447;
input v_3448;
input v_3449;
input v_3450;
input v_3451;
input v_3452;
input v_3453;
input v_3454;
input v_3455;
input v_3456;
input v_3457;
input v_3458;
input v_3459;
input v_3460;
input v_3461;
input v_3462;
input v_3463;
input v_3464;
input v_3465;
input v_3466;
input v_3467;
input v_3468;
input v_3469;
input v_3470;
input v_3471;
input v_3472;
input v_3473;
input v_3474;
input v_3475;
input v_3476;
input v_3477;
input v_3478;
input v_3479;
input v_3480;
input v_3481;
input v_3482;
input v_3483;
input v_3484;
input v_3485;
input v_3486;
input v_3487;
input v_3488;
input v_3489;
input v_3490;
input v_3491;
input v_3492;
input v_3493;
input v_3494;
input v_3495;
input v_3496;
input v_3497;
input v_3498;
input v_3499;
input v_3500;
input v_3501;
input v_3502;
input v_3503;
input v_3504;
input v_3505;
input v_3506;
input v_3507;
input v_3508;
input v_3509;
input v_3510;
input v_3511;
input v_3512;
input v_3513;
input v_3514;
input v_3515;
input v_3516;
input v_3517;
input v_3518;
input v_3519;
input v_3520;
input v_3521;
input v_3522;
input v_3523;
input v_3524;
input v_3525;
input v_3526;
input v_3527;
input v_3528;
input v_3529;
input v_3530;
input v_3531;
input v_3532;
input v_3533;
input v_3534;
input v_3535;
input v_3536;
input v_3537;
input v_3538;
input v_3539;
input v_3540;
input v_3541;
input v_3542;
input v_3543;
input v_3544;
input v_3545;
input v_3546;
input v_3547;
input v_3548;
input v_3549;
input v_3550;
input v_3551;
input v_3552;
input v_3553;
input v_3554;
input v_3555;
input v_3556;
input v_3557;
input v_3558;
input v_3559;
input v_3560;
input v_3561;
input v_3562;
input v_3563;
input v_3564;
input v_3565;
input v_3566;
input v_3567;
input v_3568;
input v_3569;
input v_3570;
input v_3571;
input v_3572;
input v_3573;
input v_3574;
input v_3575;
input v_3576;
input v_3577;
input v_3578;
input v_3579;
input v_3580;
input v_3581;
input v_3582;
input v_3583;
input v_3584;
input v_3585;
input v_3586;
input v_3587;
input v_3588;
input v_3589;
input v_3590;
input v_3591;
input v_3592;
input v_3593;
input v_3594;
input v_3595;
input v_3596;
input v_3597;
input v_3598;
input v_3599;
input v_3600;
input v_3601;
input v_3602;
input v_3603;
input v_3604;
input v_3605;
input v_3606;
input v_3607;
input v_3608;
input v_3609;
input v_3610;
input v_3611;
input v_3612;
input v_3613;
input v_3614;
input v_3615;
input v_3616;
input v_3617;
input v_3618;
input v_3619;
input v_3620;
input v_3621;
input v_3622;
input v_3623;
input v_3624;
input v_3625;
input v_3626;
input v_3627;
input v_3628;
input v_3629;
input v_3630;
input v_3631;
input v_3632;
input v_3633;
input v_3634;
input v_3635;
input v_3636;
input v_3637;
input v_3638;
input v_3639;
input v_3640;
input v_3641;
input v_3642;
input v_3643;
input v_3644;
input v_3645;
input v_3646;
input v_3647;
input v_3648;
input v_3649;
input v_3650;
input v_3651;
input v_3652;
input v_3653;
input v_3654;
input v_3655;
input v_3656;
input v_3657;
input v_3658;
input v_3659;
input v_3660;
input v_3661;
input v_3662;
input v_3663;
input v_3664;
input v_3665;
input v_3666;
input v_3667;
input v_3668;
input v_3669;
input v_3670;
input v_3671;
input v_3672;
input v_3673;
input v_3674;
input v_3675;
input v_3676;
input v_3677;
input v_3678;
input v_3679;
input v_3680;
input v_3681;
input v_3682;
input v_3683;
input v_3684;
input v_3685;
input v_3686;
input v_3687;
input v_3688;
input v_3689;
input v_3690;
input v_3691;
input v_3692;
input v_3693;
input v_3694;
input v_3695;
input v_3696;
input v_3697;
input v_3698;
input v_3699;
input v_3700;
input v_3701;
input v_3702;
input v_3703;
input v_3704;
input v_3705;
input v_3706;
input v_3707;
input v_3708;
input v_3709;
input v_3710;
input v_3711;
input v_3712;
input v_3713;
input v_3714;
input v_3715;
input v_3716;
input v_3717;
input v_3718;
input v_3719;
input v_3720;
input v_3721;
input v_3722;
input v_3723;
input v_3724;
input v_3725;
input v_3726;
input v_3727;
input v_3728;
input v_3729;
input v_3730;
input v_3731;
input v_3732;
input v_3733;
input v_3734;
input v_3735;
input v_3736;
input v_3737;
input v_3738;
input v_3739;
input v_3740;
input v_3741;
input v_3742;
input v_3743;
input v_3744;
input v_3745;
input v_3746;
input v_3747;
input v_3748;
input v_3749;
input v_3750;
input v_3751;
input v_3752;
input v_3753;
input v_3754;
input v_3755;
input v_3756;
input v_3757;
input v_3758;
input v_3759;
input v_3760;
input v_3761;
input v_3762;
input v_3763;
input v_3764;
input v_3765;
input v_3766;
input v_3767;
input v_3768;
input v_3769;
input v_3770;
input v_3771;
input v_3772;
input v_3773;
input v_3774;
input v_3775;
input v_3776;
input v_3777;
input v_3778;
input v_3779;
input v_3780;
input v_3781;
input v_3782;
input v_3783;
input v_3784;
input v_3785;
input v_3786;
input v_3787;
input v_3788;
input v_3789;
input v_3790;
input v_3791;
input v_3792;
input v_3793;
input v_3794;
input v_3795;
input v_3796;
input v_3797;
input v_3798;
input v_3799;
input v_3800;
input v_3801;
input v_3802;
input v_3803;
input v_3804;
input v_3805;
input v_3806;
input v_3807;
input v_3808;
input v_3809;
input v_3810;
input v_3811;
input v_3812;
input v_3813;
input v_3814;
input v_3815;
input v_3816;
input v_3817;
input v_3818;
input v_3819;
input v_3820;
input v_3821;
input v_3822;
input v_3823;
input v_3824;
input v_3825;
input v_3826;
input v_3827;
input v_3828;
input v_3829;
input v_3830;
input v_3831;
input v_3832;
input v_3833;
input v_3834;
input v_3835;
input v_3836;
input v_3837;
input v_3838;
input v_3839;
input v_3840;
input v_3841;
input v_3842;
input v_3843;
input v_3844;
input v_3845;
input v_3846;
input v_3847;
input v_3848;
input v_3849;
input v_3850;
input v_3851;
input v_3852;
input v_3853;
input v_3854;
input v_3855;
input v_3856;
input v_3857;
input v_3858;
input v_3859;
input v_3860;
input v_3861;
input v_3862;
input v_3863;
input v_3864;
input v_3865;
input v_3866;
input v_3867;
input v_3868;
input v_3869;
input v_3870;
input v_3871;
input v_3872;
input v_3873;
input v_3874;
input v_3875;
input v_3876;
input v_3877;
input v_3878;
input v_3879;
input v_3880;
input v_3881;
input v_3882;
input v_3883;
input v_3884;
input v_3885;
input v_3886;
input v_3887;
input v_3888;
input v_3889;
input v_3890;
input v_3891;
input v_3892;
input v_3893;
input v_3894;
input v_3895;
input v_3896;
input v_3897;
input v_3898;
input v_3899;
input v_3900;
input v_3901;
input v_3902;
input v_3903;
input v_3904;
input v_3905;
input v_3906;
input v_3907;
input v_3908;
input v_3909;
input v_3910;
input v_3911;
input v_3912;
input v_3913;
input v_3914;
input v_3915;
input v_3916;
input v_3917;
input v_3918;
input v_3919;
input v_3920;
input v_3921;
input v_3922;
input v_3923;
input v_3924;
input v_3925;
input v_3926;
input v_3927;
input v_3928;
input v_3929;
input v_3930;
input v_3931;
input v_3932;
input v_3933;
input v_3934;
input v_3935;
input v_3936;
input v_3937;
input v_3938;
input v_3939;
input v_3940;
input v_3941;
input v_3942;
input v_3943;
input v_3944;
input v_3945;
input v_3946;
input v_3947;
input v_3948;
input v_3949;
input v_3950;
input v_3951;
input v_3952;
input v_3953;
input v_3954;
input v_3955;
input v_3956;
input v_3957;
input v_3958;
input v_3959;
input v_3960;
input v_3961;
input v_3962;
input v_3963;
input v_3964;
input v_3965;
input v_3966;
input v_3967;
input v_3968;
input v_3969;
input v_3970;
input v_3971;
input v_3972;
input v_3973;
input v_3974;
input v_3975;
input v_3976;
input v_3977;
input v_3978;
input v_3979;
input v_3980;
input v_3981;
input v_3982;
input v_3983;
input v_3984;
input v_3985;
input v_3986;
input v_3987;
input v_3988;
input v_3989;
input v_3990;
input v_3991;
input v_3992;
input v_3993;
input v_3994;
input v_3995;
input v_3996;
input v_3997;
input v_3998;
input v_3999;
input v_4000;
input v_4001;
input v_4002;
input v_4003;
input v_4004;
input v_4005;
input v_4006;
input v_4007;
input v_4008;
input v_4009;
input v_4010;
input v_4011;
input v_4012;
input v_4013;
input v_4014;
input v_4015;
input v_4016;
input v_4017;
input v_4018;
input v_4019;
input v_4020;
input v_4021;
input v_4022;
input v_4023;
input v_4024;
input v_4025;
input v_4026;
input v_4027;
input v_4028;
input v_4029;
input v_4030;
input v_4031;
input v_4032;
input v_4033;
input v_4034;
input v_4035;
input v_4036;
input v_4037;
input v_4038;
input v_4039;
input v_4040;
input v_4041;
input v_4042;
input v_4043;
input v_4044;
input v_4045;
input v_4046;
input v_4047;
input v_4048;
input v_4049;
input v_4050;
input v_4051;
input v_4052;
input v_4053;
input v_4054;
input v_4055;
input v_4056;
input v_4057;
input v_4058;
input v_4059;
input v_4060;
input v_4061;
input v_4062;
input v_4063;
input v_4064;
input v_4065;
input v_4066;
input v_4067;
input v_4068;
input v_4069;
input v_4070;
input v_4071;
input v_4072;
input v_4073;
input v_4074;
input v_4075;
input v_4076;
input v_4077;
input v_4078;
input v_4079;
input v_4080;
input v_4081;
input v_4082;
input v_4083;
input v_4084;
input v_4085;
input v_4086;
input v_4087;
input v_4088;
input v_4089;
input v_4090;
input v_4091;
input v_4092;
input v_4093;
input v_4094;
input v_4095;
input v_4096;
input v_4097;
input v_4098;
input v_4099;
input v_4100;
input v_4101;
input v_4102;
input v_4103;
input v_4104;
input v_4105;
input v_4106;
input v_4107;
input v_4108;
input v_4109;
input v_4110;
input v_4111;
input v_4112;
input v_4113;
input v_4114;
input v_4115;
input v_4116;
input v_4117;
input v_4118;
input v_4119;
input v_4120;
input v_4121;
input v_4122;
input v_4123;
input v_4124;
input v_4125;
input v_4126;
input v_4127;
input v_4128;
input v_4129;
input v_4130;
input v_4131;
input v_4132;
input v_4133;
input v_4134;
input v_4135;
input v_4136;
input v_4137;
input v_4138;
input v_4139;
input v_4140;
input v_4141;
input v_4142;
input v_4143;
input v_4144;
input v_4145;
input v_4146;
input v_4147;
input v_4148;
input v_4149;
input v_4150;
input v_4151;
input v_4152;
input v_4153;
input v_4154;
input v_4155;
input v_4156;
input v_4157;
input v_4158;
input v_4159;
input v_4160;
input v_4161;
input v_4162;
input v_4163;
input v_4164;
input v_4165;
input v_4166;
input v_4167;
input v_4168;
input v_4169;
input v_4170;
input v_4171;
input v_4172;
input v_4173;
input v_4174;
input v_4175;
input v_4176;
input v_4177;
input v_4178;
input v_4179;
input v_4180;
input v_4181;
input v_4182;
input v_4183;
input v_4184;
input v_4185;
input v_4186;
input v_4187;
input v_4188;
input v_4189;
input v_4190;
input v_4191;
input v_4192;
input v_4193;
input v_4194;
input v_4195;
input v_4196;
input v_4197;
input v_4198;
input v_4199;
input v_4200;
input v_4201;
input v_4202;
input v_4203;
input v_4204;
input v_4205;
input v_4206;
input v_4207;
input v_4208;
input v_4209;
input v_4210;
input v_4211;
input v_4212;
input v_4213;
input v_4214;
input v_4215;
input v_4216;
input v_4217;
input v_4218;
input v_4219;
input v_4220;
input v_4221;
input v_4222;
input v_4223;
input v_4224;
input v_4225;
input v_4226;
input v_4227;
input v_4228;
input v_4229;
input v_4230;
input v_4231;
input v_4232;
input v_4233;
input v_4234;
input v_4235;
input v_4236;
input v_4237;
input v_4238;
input v_4239;
input v_4240;
input v_4241;
input v_4242;
input v_4243;
input v_4244;
input v_4245;
input v_4246;
input v_4247;
input v_4248;
input v_4249;
input v_4250;
input v_4251;
input v_4252;
input v_4253;
input v_4254;
input v_4255;
input v_4256;
input v_4257;
input v_4258;
input v_4259;
input v_4260;
input v_4261;
input v_4262;
input v_4263;
input v_4264;
input v_4265;
input v_4266;
input v_4267;
input v_4268;
input v_4269;
input v_4270;
input v_4271;
input v_4272;
input v_4273;
input v_4274;
input v_4275;
input v_4276;
input v_4277;
input v_4278;
input v_4279;
input v_4280;
input v_4281;
input v_4282;
input v_4283;
input v_4284;
input v_4285;
input v_4286;
input v_4287;
input v_4288;
input v_4289;
input v_4290;
input v_4291;
input v_4292;
input v_4293;
input v_4294;
input v_4295;
input v_4296;
input v_4297;
input v_4298;
input v_4299;
input v_4300;
input v_4301;
input v_4302;
input v_4303;
input v_4304;
input v_4305;
input v_4306;
input v_4307;
input v_4308;
input v_4309;
input v_4310;
input v_4311;
input v_4312;
input v_4313;
input v_4314;
input v_4315;
input v_4316;
input v_4317;
input v_4318;
input v_4319;
input v_4320;
input v_4321;
input v_4322;
input v_4323;
input v_4324;
input v_4325;
input v_4326;
input v_4327;
input v_4328;
input v_4329;
input v_4330;
input v_4331;
input v_4332;
input v_4333;
input v_4334;
input v_4335;
input v_4336;
input v_4337;
input v_4338;
input v_4339;
input v_4340;
input v_4341;
input v_4342;
input v_4343;
input v_4344;
input v_4345;
input v_4346;
input v_4347;
input v_4348;
input v_4349;
input v_4350;
input v_4351;
input v_4352;
input v_4353;
input v_4354;
input v_4355;
input v_4356;
input v_4357;
input v_4358;
input v_4359;
input v_4360;
input v_4361;
input v_4362;
input v_4363;
input v_4364;
input v_4365;
input v_4366;
input v_4367;
input v_4368;
input v_4369;
input v_4370;
input v_4371;
input v_4372;
input v_4373;
input v_4374;
input v_4375;
input v_4376;
input v_4377;
input v_4378;
input v_4379;
input v_4380;
input v_4381;
input v_4382;
input v_4383;
input v_4384;
input v_4385;
input v_4386;
input v_4387;
input v_4388;
input v_4389;
input v_4390;
input v_4391;
input v_4392;
input v_4393;
input v_4394;
input v_4395;
input v_4396;
input v_4397;
input v_4398;
input v_4399;
input v_4400;
input v_4401;
input v_4402;
input v_4403;
input v_4404;
input v_4405;
input v_4406;
input v_4407;
input v_4408;
input v_4409;
input v_4410;
input v_4411;
input v_4412;
input v_4413;
input v_4414;
input v_4415;
input v_4416;
input v_4417;
input v_4418;
input v_4419;
input v_4420;
input v_4421;
input v_4422;
input v_4423;
input v_4424;
input v_4425;
input v_4426;
input v_4427;
input v_4428;
input v_4429;
input v_4430;
input v_4431;
input v_4432;
input v_4433;
input v_4434;
input v_4435;
input v_4436;
input v_4437;
input v_4438;
input v_4439;
input v_4440;
input v_4441;
input v_4442;
input v_4443;
input v_4444;
input v_4445;
input v_4446;
input v_4447;
input v_4448;
input v_4449;
input v_4450;
input v_4451;
input v_4452;
input v_4453;
input v_4454;
input v_4455;
input v_4456;
input v_4457;
input v_4458;
input v_4459;
input v_4460;
input v_4461;
input v_4462;
input v_4463;
input v_4464;
input v_4465;
input v_4466;
input v_4467;
input v_4468;
input v_4469;
input v_4470;
input v_4471;
input v_4472;
input v_4473;
input v_4474;
input v_4475;
input v_4476;
input v_4477;
input v_4478;
input v_4479;
input v_4480;
input v_4481;
input v_4482;
input v_4483;
input v_4484;
input v_4485;
input v_4486;
input v_4487;
input v_4488;
input v_4489;
input v_4490;
input v_4491;
input v_4492;
input v_4493;
input v_4494;
input v_4495;
input v_4496;
input v_4497;
input v_4498;
input v_4499;
input v_4500;
input v_4501;
input v_4502;
input v_4503;
input v_4504;
input v_4505;
input v_4506;
input v_4507;
input v_4508;
input v_4509;
input v_4510;
input v_4511;
input v_4512;
input v_4513;
input v_4514;
input v_4515;
input v_4516;
input v_4517;
input v_4518;
input v_4519;
input v_4520;
input v_4521;
input v_4522;
input v_4523;
input v_4524;
input v_4525;
input v_4526;
input v_4527;
input v_4528;
input v_4529;
input v_4530;
input v_4531;
input v_4532;
input v_4533;
input v_4534;
input v_4535;
input v_4536;
input v_4537;
input v_4538;
input v_4539;
input v_4540;
input v_4541;
input v_4542;
input v_4543;
input v_4544;
input v_4545;
input v_4546;
input v_4547;
input v_4548;
input v_4549;
input v_4550;
input v_4551;
input v_4552;
input v_4553;
input v_4554;
input v_4555;
input v_4556;
input v_4557;
input v_4558;
input v_4559;
input v_4560;
input v_4561;
input v_4562;
input v_4563;
input v_4564;
input v_4565;
input v_4566;
input v_4567;
input v_4568;
input v_4569;
input v_4570;
input v_4571;
input v_4572;
input v_4573;
input v_4574;
input v_4575;
input v_4576;
input v_4577;
input v_4578;
input v_4579;
input v_4580;
input v_4581;
input v_4582;
input v_4583;
input v_4584;
input v_4585;
input v_4586;
input v_4587;
input v_4588;
output o_1;
wire v_4589;
wire x_1;
wire x_2;
wire x_3;
wire x_4;
wire x_5;
wire x_6;
wire x_7;
wire x_8;
wire x_9;
wire x_10;
wire x_11;
wire x_12;
wire x_13;
wire x_14;
wire x_15;
wire x_16;
wire x_17;
wire x_18;
wire x_19;
wire x_20;
wire x_21;
wire x_22;
wire x_23;
wire x_24;
wire x_25;
wire x_26;
wire x_27;
wire x_28;
wire x_29;
wire x_30;
wire x_31;
wire x_32;
wire x_33;
wire x_34;
wire x_35;
wire x_36;
wire x_37;
wire x_38;
wire x_39;
wire x_40;
wire x_41;
wire x_42;
wire x_43;
wire x_44;
wire x_45;
wire x_46;
wire x_47;
wire x_48;
wire x_49;
wire x_50;
wire x_51;
wire x_52;
wire x_53;
wire x_54;
wire x_55;
wire x_56;
wire x_57;
wire x_58;
wire x_59;
wire x_60;
wire x_61;
wire x_62;
wire x_63;
wire x_64;
wire x_65;
wire x_66;
wire x_67;
wire x_68;
wire x_69;
wire x_70;
wire x_71;
wire x_72;
wire x_73;
wire x_74;
wire x_75;
wire x_76;
wire x_77;
wire x_78;
wire x_79;
wire x_80;
wire x_81;
wire x_82;
wire x_83;
wire x_84;
wire x_85;
wire x_86;
wire x_87;
wire x_88;
wire x_89;
wire x_90;
wire x_91;
wire x_92;
wire x_93;
wire x_94;
wire x_95;
wire x_96;
wire x_97;
wire x_98;
wire x_99;
wire x_100;
wire x_101;
wire x_102;
wire x_103;
wire x_104;
wire x_105;
wire x_106;
wire x_107;
wire x_108;
wire x_109;
wire x_110;
wire x_111;
wire x_112;
wire x_113;
wire x_114;
wire x_115;
wire x_116;
wire x_117;
wire x_118;
wire x_119;
wire x_120;
wire x_121;
wire x_122;
wire x_123;
wire x_124;
wire x_125;
wire x_126;
wire x_127;
wire x_128;
wire x_129;
wire x_130;
wire x_131;
wire x_132;
wire x_133;
wire x_134;
wire x_135;
wire x_136;
wire x_137;
wire x_138;
wire x_139;
wire x_140;
wire x_141;
wire x_142;
wire x_143;
wire x_144;
wire x_145;
wire x_146;
wire x_147;
wire x_148;
wire x_149;
wire x_150;
wire x_151;
wire x_152;
wire x_153;
wire x_154;
wire x_155;
wire x_156;
wire x_157;
wire x_158;
wire x_159;
wire x_160;
wire x_161;
wire x_162;
wire x_163;
wire x_164;
wire x_165;
wire x_166;
wire x_167;
wire x_168;
wire x_169;
wire x_170;
wire x_171;
wire x_172;
wire x_173;
wire x_174;
wire x_175;
wire x_176;
wire x_177;
wire x_178;
wire x_179;
wire x_180;
wire x_181;
wire x_182;
wire x_183;
wire x_184;
wire x_185;
wire x_186;
wire x_187;
wire x_188;
wire x_189;
wire x_190;
wire x_191;
wire x_192;
wire x_193;
wire x_194;
wire x_195;
wire x_196;
wire x_197;
wire x_198;
wire x_199;
wire x_200;
wire x_201;
wire x_202;
wire x_203;
wire x_204;
wire x_205;
wire x_206;
wire x_207;
wire x_208;
wire x_209;
wire x_210;
wire x_211;
wire x_212;
wire x_213;
wire x_214;
wire x_215;
wire x_216;
wire x_217;
wire x_218;
wire x_219;
wire x_220;
wire x_221;
wire x_222;
wire x_223;
wire x_224;
wire x_225;
wire x_226;
wire x_227;
wire x_228;
wire x_229;
wire x_230;
wire x_231;
wire x_232;
wire x_233;
wire x_234;
wire x_235;
wire x_236;
wire x_237;
wire x_238;
wire x_239;
wire x_240;
wire x_241;
wire x_242;
wire x_243;
wire x_244;
wire x_245;
wire x_246;
wire x_247;
wire x_248;
wire x_249;
wire x_250;
wire x_251;
wire x_252;
wire x_253;
wire x_254;
wire x_255;
wire x_256;
wire x_257;
wire x_258;
wire x_259;
wire x_260;
wire x_261;
wire x_262;
wire x_263;
wire x_264;
wire x_265;
wire x_266;
wire x_267;
wire x_268;
wire x_269;
wire x_270;
wire x_271;
wire x_272;
wire x_273;
wire x_274;
wire x_275;
wire x_276;
wire x_277;
wire x_278;
wire x_279;
wire x_280;
wire x_281;
wire x_282;
wire x_283;
wire x_284;
wire x_285;
wire x_286;
wire x_287;
wire x_288;
wire x_289;
wire x_290;
wire x_291;
wire x_292;
wire x_293;
wire x_294;
wire x_295;
wire x_296;
wire x_297;
wire x_298;
wire x_299;
wire x_300;
wire x_301;
wire x_302;
wire x_303;
wire x_304;
wire x_305;
wire x_306;
wire x_307;
wire x_308;
wire x_309;
wire x_310;
wire x_311;
wire x_312;
wire x_313;
wire x_314;
wire x_315;
wire x_316;
wire x_317;
wire x_318;
wire x_319;
wire x_320;
wire x_321;
wire x_322;
wire x_323;
wire x_324;
wire x_325;
wire x_326;
wire x_327;
wire x_328;
wire x_329;
wire x_330;
wire x_331;
wire x_332;
wire x_333;
wire x_334;
wire x_335;
wire x_336;
wire x_337;
wire x_338;
wire x_339;
wire x_340;
wire x_341;
wire x_342;
wire x_343;
wire x_344;
wire x_345;
wire x_346;
wire x_347;
wire x_348;
wire x_349;
wire x_350;
wire x_351;
wire x_352;
wire x_353;
wire x_354;
wire x_355;
wire x_356;
wire x_357;
wire x_358;
wire x_359;
wire x_360;
wire x_361;
wire x_362;
wire x_363;
wire x_364;
wire x_365;
wire x_366;
wire x_367;
wire x_368;
wire x_369;
wire x_370;
wire x_371;
wire x_372;
wire x_373;
wire x_374;
wire x_375;
wire x_376;
wire x_377;
wire x_378;
wire x_379;
wire x_380;
wire x_381;
wire x_382;
wire x_383;
wire x_384;
wire x_385;
wire x_386;
wire x_387;
wire x_388;
wire x_389;
wire x_390;
wire x_391;
wire x_392;
wire x_393;
wire x_394;
wire x_395;
wire x_396;
wire x_397;
wire x_398;
wire x_399;
wire x_400;
wire x_401;
wire x_402;
wire x_403;
wire x_404;
wire x_405;
wire x_406;
wire x_407;
wire x_408;
wire x_409;
wire x_410;
wire x_411;
wire x_412;
wire x_413;
wire x_414;
wire x_415;
wire x_416;
wire x_417;
wire x_418;
wire x_419;
wire x_420;
wire x_421;
wire x_422;
wire x_423;
wire x_424;
wire x_425;
wire x_426;
wire x_427;
wire x_428;
wire x_429;
wire x_430;
wire x_431;
wire x_432;
wire x_433;
wire x_434;
wire x_435;
wire x_436;
wire x_437;
wire x_438;
wire x_439;
wire x_440;
wire x_441;
wire x_442;
wire x_443;
wire x_444;
wire x_445;
wire x_446;
wire x_447;
wire x_448;
wire x_449;
wire x_450;
wire x_451;
wire x_452;
wire x_453;
wire x_454;
wire x_455;
wire x_456;
wire x_457;
wire x_458;
wire x_459;
wire x_460;
wire x_461;
wire x_462;
wire x_463;
wire x_464;
wire x_465;
wire x_466;
wire x_467;
wire x_468;
wire x_469;
wire x_470;
wire x_471;
wire x_472;
wire x_473;
wire x_474;
wire x_475;
wire x_476;
wire x_477;
wire x_478;
wire x_479;
wire x_480;
wire x_481;
wire x_482;
wire x_483;
wire x_484;
wire x_485;
wire x_486;
wire x_487;
wire x_488;
wire x_489;
wire x_490;
wire x_491;
wire x_492;
wire x_493;
wire x_494;
wire x_495;
wire x_496;
wire x_497;
wire x_498;
wire x_499;
wire x_500;
wire x_501;
wire x_502;
wire x_503;
wire x_504;
wire x_505;
wire x_506;
wire x_507;
wire x_508;
wire x_509;
wire x_510;
wire x_511;
wire x_512;
wire x_513;
wire x_514;
wire x_515;
wire x_516;
wire x_517;
wire x_518;
wire x_519;
wire x_520;
wire x_521;
wire x_522;
wire x_523;
wire x_524;
wire x_525;
wire x_526;
wire x_527;
wire x_528;
wire x_529;
wire x_530;
wire x_531;
wire x_532;
wire x_533;
wire x_534;
wire x_535;
wire x_536;
wire x_537;
wire x_538;
wire x_539;
wire x_540;
wire x_541;
wire x_542;
wire x_543;
wire x_544;
wire x_545;
wire x_546;
wire x_547;
wire x_548;
wire x_549;
wire x_550;
wire x_551;
wire x_552;
wire x_553;
wire x_554;
wire x_555;
wire x_556;
wire x_557;
wire x_558;
wire x_559;
wire x_560;
wire x_561;
wire x_562;
wire x_563;
wire x_564;
wire x_565;
wire x_566;
wire x_567;
wire x_568;
wire x_569;
wire x_570;
wire x_571;
wire x_572;
wire x_573;
wire x_574;
wire x_575;
wire x_576;
wire x_577;
wire x_578;
wire x_579;
wire x_580;
wire x_581;
wire x_582;
wire x_583;
wire x_584;
wire x_585;
wire x_586;
wire x_587;
wire x_588;
wire x_589;
wire x_590;
wire x_591;
wire x_592;
wire x_593;
wire x_594;
wire x_595;
wire x_596;
wire x_597;
wire x_598;
wire x_599;
wire x_600;
wire x_601;
wire x_602;
wire x_603;
wire x_604;
wire x_605;
wire x_606;
wire x_607;
wire x_608;
wire x_609;
wire x_610;
wire x_611;
wire x_612;
wire x_613;
wire x_614;
wire x_615;
wire x_616;
wire x_617;
wire x_618;
wire x_619;
wire x_620;
wire x_621;
wire x_622;
wire x_623;
wire x_624;
wire x_625;
wire x_626;
wire x_627;
wire x_628;
wire x_629;
wire x_630;
wire x_631;
wire x_632;
wire x_633;
wire x_634;
wire x_635;
wire x_636;
wire x_637;
wire x_638;
wire x_639;
wire x_640;
wire x_641;
wire x_642;
wire x_643;
wire x_644;
wire x_645;
wire x_646;
wire x_647;
wire x_648;
wire x_649;
wire x_650;
wire x_651;
wire x_652;
wire x_653;
wire x_654;
wire x_655;
wire x_656;
wire x_657;
wire x_658;
wire x_659;
wire x_660;
wire x_661;
wire x_662;
wire x_663;
wire x_664;
wire x_665;
wire x_666;
wire x_667;
wire x_668;
wire x_669;
wire x_670;
wire x_671;
wire x_672;
wire x_673;
wire x_674;
wire x_675;
wire x_676;
wire x_677;
wire x_678;
wire x_679;
wire x_680;
wire x_681;
wire x_682;
wire x_683;
wire x_684;
wire x_685;
wire x_686;
wire x_687;
wire x_688;
wire x_689;
wire x_690;
wire x_691;
wire x_692;
wire x_693;
wire x_694;
wire x_695;
wire x_696;
wire x_697;
wire x_698;
wire x_699;
wire x_700;
wire x_701;
wire x_702;
wire x_703;
wire x_704;
wire x_705;
wire x_706;
wire x_707;
wire x_708;
wire x_709;
wire x_710;
wire x_711;
wire x_712;
wire x_713;
wire x_714;
wire x_715;
wire x_716;
wire x_717;
wire x_718;
wire x_719;
wire x_720;
wire x_721;
wire x_722;
wire x_723;
wire x_724;
wire x_725;
wire x_726;
wire x_727;
wire x_728;
wire x_729;
wire x_730;
wire x_731;
wire x_732;
wire x_733;
wire x_734;
wire x_735;
wire x_736;
wire x_737;
wire x_738;
wire x_739;
wire x_740;
wire x_741;
wire x_742;
wire x_743;
wire x_744;
wire x_745;
wire x_746;
wire x_747;
wire x_748;
wire x_749;
wire x_750;
wire x_751;
wire x_752;
wire x_753;
wire x_754;
wire x_755;
wire x_756;
wire x_757;
wire x_758;
wire x_759;
wire x_760;
wire x_761;
wire x_762;
wire x_763;
wire x_764;
wire x_765;
wire x_766;
wire x_767;
wire x_768;
wire x_769;
wire x_770;
wire x_771;
wire x_772;
wire x_773;
wire x_774;
wire x_775;
wire x_776;
wire x_777;
wire x_778;
wire x_779;
wire x_780;
wire x_781;
wire x_782;
wire x_783;
wire x_784;
wire x_785;
wire x_786;
wire x_787;
wire x_788;
wire x_789;
wire x_790;
wire x_791;
wire x_792;
wire x_793;
wire x_794;
wire x_795;
wire x_796;
wire x_797;
wire x_798;
wire x_799;
wire x_800;
wire x_801;
wire x_802;
wire x_803;
wire x_804;
wire x_805;
wire x_806;
wire x_807;
wire x_808;
wire x_809;
wire x_810;
wire x_811;
wire x_812;
wire x_813;
wire x_814;
wire x_815;
wire x_816;
wire x_817;
wire x_818;
wire x_819;
wire x_820;
wire x_821;
wire x_822;
wire x_823;
wire x_824;
wire x_825;
wire x_826;
wire x_827;
wire x_828;
wire x_829;
wire x_830;
wire x_831;
wire x_832;
wire x_833;
wire x_834;
wire x_835;
wire x_836;
wire x_837;
wire x_838;
wire x_839;
wire x_840;
wire x_841;
wire x_842;
wire x_843;
wire x_844;
wire x_845;
wire x_846;
wire x_847;
wire x_848;
wire x_849;
wire x_850;
wire x_851;
wire x_852;
wire x_853;
wire x_854;
wire x_855;
wire x_856;
wire x_857;
wire x_858;
wire x_859;
wire x_860;
wire x_861;
wire x_862;
wire x_863;
wire x_864;
wire x_865;
wire x_866;
wire x_867;
wire x_868;
wire x_869;
wire x_870;
wire x_871;
wire x_872;
wire x_873;
wire x_874;
wire x_875;
wire x_876;
wire x_877;
wire x_878;
wire x_879;
wire x_880;
wire x_881;
wire x_882;
wire x_883;
wire x_884;
wire x_885;
wire x_886;
wire x_887;
wire x_888;
wire x_889;
wire x_890;
wire x_891;
wire x_892;
wire x_893;
wire x_894;
wire x_895;
wire x_896;
wire x_897;
wire x_898;
wire x_899;
wire x_900;
wire x_901;
wire x_902;
wire x_903;
wire x_904;
wire x_905;
wire x_906;
wire x_907;
wire x_908;
wire x_909;
wire x_910;
wire x_911;
wire x_912;
wire x_913;
wire x_914;
wire x_915;
wire x_916;
wire x_917;
wire x_918;
wire x_919;
wire x_920;
wire x_921;
wire x_922;
wire x_923;
wire x_924;
wire x_925;
wire x_926;
wire x_927;
wire x_928;
wire x_929;
wire x_930;
wire x_931;
wire x_932;
wire x_933;
wire x_934;
wire x_935;
wire x_936;
wire x_937;
wire x_938;
wire x_939;
wire x_940;
wire x_941;
wire x_942;
wire x_943;
wire x_944;
wire x_945;
wire x_946;
wire x_947;
wire x_948;
wire x_949;
wire x_950;
wire x_951;
wire x_952;
wire x_953;
wire x_954;
wire x_955;
wire x_956;
wire x_957;
wire x_958;
wire x_959;
wire x_960;
wire x_961;
wire x_962;
wire x_963;
wire x_964;
wire x_965;
wire x_966;
wire x_967;
wire x_968;
wire x_969;
wire x_970;
wire x_971;
wire x_972;
wire x_973;
wire x_974;
wire x_975;
wire x_976;
wire x_977;
wire x_978;
wire x_979;
wire x_980;
wire x_981;
wire x_982;
wire x_983;
wire x_984;
wire x_985;
wire x_986;
wire x_987;
wire x_988;
wire x_989;
wire x_990;
wire x_991;
wire x_992;
wire x_993;
wire x_994;
wire x_995;
wire x_996;
wire x_997;
wire x_998;
wire x_999;
wire x_1000;
wire x_1001;
wire x_1002;
wire x_1003;
wire x_1004;
wire x_1005;
wire x_1006;
wire x_1007;
wire x_1008;
wire x_1009;
wire x_1010;
wire x_1011;
wire x_1012;
wire x_1013;
wire x_1014;
wire x_1015;
wire x_1016;
wire x_1017;
wire x_1018;
wire x_1019;
wire x_1020;
wire x_1021;
wire x_1022;
wire x_1023;
wire x_1024;
wire x_1025;
wire x_1026;
wire x_1027;
wire x_1028;
wire x_1029;
wire x_1030;
wire x_1031;
wire x_1032;
wire x_1033;
wire x_1034;
wire x_1035;
wire x_1036;
wire x_1037;
wire x_1038;
wire x_1039;
wire x_1040;
wire x_1041;
wire x_1042;
wire x_1043;
wire x_1044;
wire x_1045;
wire x_1046;
wire x_1047;
wire x_1048;
wire x_1049;
wire x_1050;
wire x_1051;
wire x_1052;
wire x_1053;
wire x_1054;
wire x_1055;
wire x_1056;
wire x_1057;
wire x_1058;
wire x_1059;
wire x_1060;
wire x_1061;
wire x_1062;
wire x_1063;
wire x_1064;
wire x_1065;
wire x_1066;
wire x_1067;
wire x_1068;
wire x_1069;
wire x_1070;
wire x_1071;
wire x_1072;
wire x_1073;
wire x_1074;
wire x_1075;
wire x_1076;
wire x_1077;
wire x_1078;
wire x_1079;
wire x_1080;
wire x_1081;
wire x_1082;
wire x_1083;
wire x_1084;
wire x_1085;
wire x_1086;
wire x_1087;
wire x_1088;
wire x_1089;
wire x_1090;
wire x_1091;
wire x_1092;
wire x_1093;
wire x_1094;
wire x_1095;
wire x_1096;
wire x_1097;
wire x_1098;
wire x_1099;
wire x_1100;
wire x_1101;
wire x_1102;
wire x_1103;
wire x_1104;
wire x_1105;
wire x_1106;
wire x_1107;
wire x_1108;
wire x_1109;
wire x_1110;
wire x_1111;
wire x_1112;
wire x_1113;
wire x_1114;
wire x_1115;
wire x_1116;
wire x_1117;
wire x_1118;
wire x_1119;
wire x_1120;
wire x_1121;
wire x_1122;
wire x_1123;
wire x_1124;
wire x_1125;
wire x_1126;
wire x_1127;
wire x_1128;
wire x_1129;
wire x_1130;
wire x_1131;
wire x_1132;
wire x_1133;
wire x_1134;
wire x_1135;
wire x_1136;
wire x_1137;
wire x_1138;
wire x_1139;
wire x_1140;
wire x_1141;
wire x_1142;
wire x_1143;
wire x_1144;
wire x_1145;
wire x_1146;
wire x_1147;
wire x_1148;
wire x_1149;
wire x_1150;
wire x_1151;
wire x_1152;
wire x_1153;
wire x_1154;
wire x_1155;
wire x_1156;
wire x_1157;
wire x_1158;
wire x_1159;
wire x_1160;
wire x_1161;
wire x_1162;
wire x_1163;
wire x_1164;
wire x_1165;
wire x_1166;
wire x_1167;
wire x_1168;
wire x_1169;
wire x_1170;
wire x_1171;
wire x_1172;
wire x_1173;
wire x_1174;
wire x_1175;
wire x_1176;
wire x_1177;
wire x_1178;
wire x_1179;
wire x_1180;
wire x_1181;
wire x_1182;
wire x_1183;
wire x_1184;
wire x_1185;
wire x_1186;
wire x_1187;
wire x_1188;
wire x_1189;
wire x_1190;
wire x_1191;
wire x_1192;
wire x_1193;
wire x_1194;
wire x_1195;
wire x_1196;
wire x_1197;
wire x_1198;
wire x_1199;
wire x_1200;
wire x_1201;
wire x_1202;
wire x_1203;
wire x_1204;
wire x_1205;
wire x_1206;
wire x_1207;
wire x_1208;
wire x_1209;
wire x_1210;
wire x_1211;
wire x_1212;
wire x_1213;
wire x_1214;
wire x_1215;
wire x_1216;
wire x_1217;
wire x_1218;
wire x_1219;
wire x_1220;
wire x_1221;
wire x_1222;
wire x_1223;
wire x_1224;
wire x_1225;
wire x_1226;
wire x_1227;
wire x_1228;
wire x_1229;
wire x_1230;
wire x_1231;
wire x_1232;
wire x_1233;
wire x_1234;
wire x_1235;
wire x_1236;
wire x_1237;
wire x_1238;
wire x_1239;
wire x_1240;
wire x_1241;
wire x_1242;
wire x_1243;
wire x_1244;
wire x_1245;
wire x_1246;
wire x_1247;
wire x_1248;
wire x_1249;
wire x_1250;
wire x_1251;
wire x_1252;
wire x_1253;
wire x_1254;
wire x_1255;
wire x_1256;
wire x_1257;
wire x_1258;
wire x_1259;
wire x_1260;
wire x_1261;
wire x_1262;
wire x_1263;
wire x_1264;
wire x_1265;
wire x_1266;
wire x_1267;
wire x_1268;
wire x_1269;
wire x_1270;
wire x_1271;
wire x_1272;
wire x_1273;
wire x_1274;
wire x_1275;
wire x_1276;
wire x_1277;
wire x_1278;
wire x_1279;
wire x_1280;
wire x_1281;
wire x_1282;
wire x_1283;
wire x_1284;
wire x_1285;
wire x_1286;
wire x_1287;
wire x_1288;
wire x_1289;
wire x_1290;
wire x_1291;
wire x_1292;
wire x_1293;
wire x_1294;
wire x_1295;
wire x_1296;
wire x_1297;
wire x_1298;
wire x_1299;
wire x_1300;
wire x_1301;
wire x_1302;
wire x_1303;
wire x_1304;
wire x_1305;
wire x_1306;
wire x_1307;
wire x_1308;
wire x_1309;
wire x_1310;
wire x_1311;
wire x_1312;
wire x_1313;
wire x_1314;
wire x_1315;
wire x_1316;
wire x_1317;
wire x_1318;
wire x_1319;
wire x_1320;
wire x_1321;
wire x_1322;
wire x_1323;
wire x_1324;
wire x_1325;
wire x_1326;
wire x_1327;
wire x_1328;
wire x_1329;
wire x_1330;
wire x_1331;
wire x_1332;
wire x_1333;
wire x_1334;
wire x_1335;
wire x_1336;
wire x_1337;
wire x_1338;
wire x_1339;
wire x_1340;
wire x_1341;
wire x_1342;
wire x_1343;
wire x_1344;
wire x_1345;
wire x_1346;
wire x_1347;
wire x_1348;
wire x_1349;
wire x_1350;
wire x_1351;
wire x_1352;
wire x_1353;
wire x_1354;
wire x_1355;
wire x_1356;
wire x_1357;
wire x_1358;
wire x_1359;
wire x_1360;
wire x_1361;
wire x_1362;
wire x_1363;
wire x_1364;
wire x_1365;
wire x_1366;
wire x_1367;
wire x_1368;
wire x_1369;
wire x_1370;
wire x_1371;
wire x_1372;
wire x_1373;
wire x_1374;
wire x_1375;
wire x_1376;
wire x_1377;
wire x_1378;
wire x_1379;
wire x_1380;
wire x_1381;
wire x_1382;
wire x_1383;
wire x_1384;
wire x_1385;
wire x_1386;
wire x_1387;
wire x_1388;
wire x_1389;
wire x_1390;
wire x_1391;
wire x_1392;
wire x_1393;
wire x_1394;
wire x_1395;
wire x_1396;
wire x_1397;
wire x_1398;
wire x_1399;
wire x_1400;
wire x_1401;
wire x_1402;
wire x_1403;
wire x_1404;
wire x_1405;
wire x_1406;
wire x_1407;
wire x_1408;
wire x_1409;
wire x_1410;
wire x_1411;
wire x_1412;
wire x_1413;
wire x_1414;
wire x_1415;
wire x_1416;
wire x_1417;
wire x_1418;
wire x_1419;
wire x_1420;
wire x_1421;
wire x_1422;
wire x_1423;
wire x_1424;
wire x_1425;
wire x_1426;
wire x_1427;
wire x_1428;
wire x_1429;
wire x_1430;
wire x_1431;
wire x_1432;
wire x_1433;
wire x_1434;
wire x_1435;
wire x_1436;
wire x_1437;
wire x_1438;
wire x_1439;
wire x_1440;
wire x_1441;
wire x_1442;
wire x_1443;
wire x_1444;
wire x_1445;
wire x_1446;
wire x_1447;
wire x_1448;
wire x_1449;
wire x_1450;
wire x_1451;
wire x_1452;
wire x_1453;
wire x_1454;
wire x_1455;
wire x_1456;
wire x_1457;
wire x_1458;
wire x_1459;
wire x_1460;
wire x_1461;
wire x_1462;
wire x_1463;
wire x_1464;
wire x_1465;
wire x_1466;
wire x_1467;
wire x_1468;
wire x_1469;
wire x_1470;
wire x_1471;
wire x_1472;
wire x_1473;
wire x_1474;
wire x_1475;
wire x_1476;
wire x_1477;
wire x_1478;
wire x_1479;
wire x_1480;
wire x_1481;
wire x_1482;
wire x_1483;
wire x_1484;
wire x_1485;
wire x_1486;
wire x_1487;
wire x_1488;
wire x_1489;
wire x_1490;
wire x_1491;
wire x_1492;
wire x_1493;
wire x_1494;
wire x_1495;
wire x_1496;
wire x_1497;
wire x_1498;
wire x_1499;
wire x_1500;
wire x_1501;
wire x_1502;
wire x_1503;
wire x_1504;
wire x_1505;
wire x_1506;
wire x_1507;
wire x_1508;
wire x_1509;
wire x_1510;
wire x_1511;
wire x_1512;
wire x_1513;
wire x_1514;
wire x_1515;
wire x_1516;
wire x_1517;
wire x_1518;
wire x_1519;
wire x_1520;
wire x_1521;
wire x_1522;
wire x_1523;
wire x_1524;
wire x_1525;
wire x_1526;
wire x_1527;
wire x_1528;
wire x_1529;
wire x_1530;
wire x_1531;
wire x_1532;
wire x_1533;
wire x_1534;
wire x_1535;
wire x_1536;
wire x_1537;
wire x_1538;
wire x_1539;
wire x_1540;
wire x_1541;
wire x_1542;
wire x_1543;
wire x_1544;
wire x_1545;
wire x_1546;
wire x_1547;
wire x_1548;
wire x_1549;
wire x_1550;
wire x_1551;
wire x_1552;
wire x_1553;
wire x_1554;
wire x_1555;
wire x_1556;
wire x_1557;
wire x_1558;
wire x_1559;
wire x_1560;
wire x_1561;
wire x_1562;
wire x_1563;
wire x_1564;
wire x_1565;
wire x_1566;
wire x_1567;
wire x_1568;
wire x_1569;
wire x_1570;
wire x_1571;
wire x_1572;
wire x_1573;
wire x_1574;
wire x_1575;
wire x_1576;
wire x_1577;
wire x_1578;
wire x_1579;
wire x_1580;
wire x_1581;
wire x_1582;
wire x_1583;
wire x_1584;
wire x_1585;
wire x_1586;
wire x_1587;
wire x_1588;
wire x_1589;
wire x_1590;
wire x_1591;
wire x_1592;
wire x_1593;
wire x_1594;
wire x_1595;
wire x_1596;
wire x_1597;
wire x_1598;
wire x_1599;
wire x_1600;
wire x_1601;
wire x_1602;
wire x_1603;
wire x_1604;
wire x_1605;
wire x_1606;
wire x_1607;
wire x_1608;
wire x_1609;
wire x_1610;
wire x_1611;
wire x_1612;
wire x_1613;
wire x_1614;
wire x_1615;
wire x_1616;
wire x_1617;
wire x_1618;
wire x_1619;
wire x_1620;
wire x_1621;
wire x_1622;
wire x_1623;
wire x_1624;
wire x_1625;
wire x_1626;
wire x_1627;
wire x_1628;
wire x_1629;
wire x_1630;
wire x_1631;
wire x_1632;
wire x_1633;
wire x_1634;
wire x_1635;
wire x_1636;
wire x_1637;
wire x_1638;
wire x_1639;
wire x_1640;
wire x_1641;
wire x_1642;
wire x_1643;
wire x_1644;
wire x_1645;
wire x_1646;
wire x_1647;
wire x_1648;
wire x_1649;
wire x_1650;
wire x_1651;
wire x_1652;
wire x_1653;
wire x_1654;
wire x_1655;
wire x_1656;
wire x_1657;
wire x_1658;
wire x_1659;
wire x_1660;
wire x_1661;
wire x_1662;
wire x_1663;
wire x_1664;
wire x_1665;
wire x_1666;
wire x_1667;
wire x_1668;
wire x_1669;
wire x_1670;
wire x_1671;
wire x_1672;
wire x_1673;
wire x_1674;
wire x_1675;
wire x_1676;
wire x_1677;
wire x_1678;
wire x_1679;
wire x_1680;
wire x_1681;
wire x_1682;
wire x_1683;
wire x_1684;
wire x_1685;
wire x_1686;
wire x_1687;
wire x_1688;
wire x_1689;
wire x_1690;
wire x_1691;
wire x_1692;
wire x_1693;
wire x_1694;
wire x_1695;
wire x_1696;
wire x_1697;
wire x_1698;
wire x_1699;
wire x_1700;
wire x_1701;
wire x_1702;
wire x_1703;
wire x_1704;
wire x_1705;
wire x_1706;
wire x_1707;
wire x_1708;
wire x_1709;
wire x_1710;
wire x_1711;
wire x_1712;
wire x_1713;
wire x_1714;
wire x_1715;
wire x_1716;
wire x_1717;
wire x_1718;
wire x_1719;
wire x_1720;
wire x_1721;
wire x_1722;
wire x_1723;
wire x_1724;
wire x_1725;
wire x_1726;
wire x_1727;
wire x_1728;
wire x_1729;
wire x_1730;
wire x_1731;
wire x_1732;
wire x_1733;
wire x_1734;
wire x_1735;
wire x_1736;
wire x_1737;
wire x_1738;
wire x_1739;
wire x_1740;
wire x_1741;
wire x_1742;
wire x_1743;
wire x_1744;
wire x_1745;
wire x_1746;
wire x_1747;
wire x_1748;
wire x_1749;
wire x_1750;
wire x_1751;
wire x_1752;
wire x_1753;
wire x_1754;
wire x_1755;
wire x_1756;
wire x_1757;
wire x_1758;
wire x_1759;
wire x_1760;
wire x_1761;
wire x_1762;
wire x_1763;
wire x_1764;
wire x_1765;
wire x_1766;
wire x_1767;
wire x_1768;
wire x_1769;
wire x_1770;
wire x_1771;
wire x_1772;
wire x_1773;
wire x_1774;
wire x_1775;
wire x_1776;
wire x_1777;
wire x_1778;
wire x_1779;
wire x_1780;
wire x_1781;
wire x_1782;
wire x_1783;
wire x_1784;
wire x_1785;
wire x_1786;
wire x_1787;
wire x_1788;
wire x_1789;
wire x_1790;
wire x_1791;
wire x_1792;
wire x_1793;
wire x_1794;
wire x_1795;
wire x_1796;
wire x_1797;
wire x_1798;
wire x_1799;
wire x_1800;
wire x_1801;
wire x_1802;
wire x_1803;
wire x_1804;
wire x_1805;
wire x_1806;
wire x_1807;
wire x_1808;
wire x_1809;
wire x_1810;
wire x_1811;
wire x_1812;
wire x_1813;
wire x_1814;
wire x_1815;
wire x_1816;
wire x_1817;
wire x_1818;
wire x_1819;
wire x_1820;
wire x_1821;
wire x_1822;
wire x_1823;
wire x_1824;
wire x_1825;
wire x_1826;
wire x_1827;
wire x_1828;
wire x_1829;
wire x_1830;
wire x_1831;
wire x_1832;
wire x_1833;
wire x_1834;
wire x_1835;
wire x_1836;
wire x_1837;
wire x_1838;
wire x_1839;
wire x_1840;
wire x_1841;
wire x_1842;
wire x_1843;
wire x_1844;
wire x_1845;
wire x_1846;
wire x_1847;
wire x_1848;
wire x_1849;
wire x_1850;
wire x_1851;
wire x_1852;
wire x_1853;
wire x_1854;
wire x_1855;
wire x_1856;
wire x_1857;
wire x_1858;
wire x_1859;
wire x_1860;
wire x_1861;
wire x_1862;
wire x_1863;
wire x_1864;
wire x_1865;
wire x_1866;
wire x_1867;
wire x_1868;
wire x_1869;
wire x_1870;
wire x_1871;
wire x_1872;
wire x_1873;
wire x_1874;
wire x_1875;
wire x_1876;
wire x_1877;
wire x_1878;
wire x_1879;
wire x_1880;
wire x_1881;
wire x_1882;
wire x_1883;
wire x_1884;
wire x_1885;
wire x_1886;
wire x_1887;
wire x_1888;
wire x_1889;
wire x_1890;
wire x_1891;
wire x_1892;
wire x_1893;
wire x_1894;
wire x_1895;
wire x_1896;
wire x_1897;
wire x_1898;
wire x_1899;
wire x_1900;
wire x_1901;
wire x_1902;
wire x_1903;
wire x_1904;
wire x_1905;
wire x_1906;
wire x_1907;
wire x_1908;
wire x_1909;
wire x_1910;
wire x_1911;
wire x_1912;
wire x_1913;
wire x_1914;
wire x_1915;
wire x_1916;
wire x_1917;
wire x_1918;
wire x_1919;
wire x_1920;
wire x_1921;
wire x_1922;
wire x_1923;
wire x_1924;
wire x_1925;
wire x_1926;
wire x_1927;
wire x_1928;
wire x_1929;
wire x_1930;
wire x_1931;
wire x_1932;
wire x_1933;
wire x_1934;
wire x_1935;
wire x_1936;
wire x_1937;
wire x_1938;
wire x_1939;
wire x_1940;
wire x_1941;
wire x_1942;
wire x_1943;
wire x_1944;
wire x_1945;
wire x_1946;
wire x_1947;
wire x_1948;
wire x_1949;
wire x_1950;
wire x_1951;
wire x_1952;
wire x_1953;
wire x_1954;
wire x_1955;
wire x_1956;
wire x_1957;
wire x_1958;
wire x_1959;
wire x_1960;
wire x_1961;
wire x_1962;
wire x_1963;
wire x_1964;
wire x_1965;
wire x_1966;
wire x_1967;
wire x_1968;
wire x_1969;
wire x_1970;
wire x_1971;
wire x_1972;
wire x_1973;
wire x_1974;
wire x_1975;
wire x_1976;
wire x_1977;
wire x_1978;
wire x_1979;
wire x_1980;
wire x_1981;
wire x_1982;
wire x_1983;
wire x_1984;
wire x_1985;
wire x_1986;
wire x_1987;
wire x_1988;
wire x_1989;
wire x_1990;
wire x_1991;
wire x_1992;
wire x_1993;
wire x_1994;
wire x_1995;
wire x_1996;
wire x_1997;
wire x_1998;
wire x_1999;
wire x_2000;
wire x_2001;
wire x_2002;
wire x_2003;
wire x_2004;
wire x_2005;
wire x_2006;
wire x_2007;
wire x_2008;
wire x_2009;
wire x_2010;
wire x_2011;
wire x_2012;
wire x_2013;
wire x_2014;
wire x_2015;
wire x_2016;
wire x_2017;
wire x_2018;
wire x_2019;
wire x_2020;
wire x_2021;
wire x_2022;
wire x_2023;
wire x_2024;
wire x_2025;
wire x_2026;
wire x_2027;
wire x_2028;
wire x_2029;
wire x_2030;
wire x_2031;
wire x_2032;
wire x_2033;
wire x_2034;
wire x_2035;
wire x_2036;
wire x_2037;
wire x_2038;
wire x_2039;
wire x_2040;
wire x_2041;
wire x_2042;
wire x_2043;
wire x_2044;
wire x_2045;
wire x_2046;
wire x_2047;
wire x_2048;
wire x_2049;
wire x_2050;
wire x_2051;
wire x_2052;
wire x_2053;
wire x_2054;
wire x_2055;
wire x_2056;
wire x_2057;
wire x_2058;
wire x_2059;
wire x_2060;
wire x_2061;
wire x_2062;
wire x_2063;
wire x_2064;
wire x_2065;
wire x_2066;
wire x_2067;
wire x_2068;
wire x_2069;
wire x_2070;
wire x_2071;
wire x_2072;
wire x_2073;
wire x_2074;
wire x_2075;
wire x_2076;
wire x_2077;
wire x_2078;
wire x_2079;
wire x_2080;
wire x_2081;
wire x_2082;
wire x_2083;
wire x_2084;
wire x_2085;
wire x_2086;
wire x_2087;
wire x_2088;
wire x_2089;
wire x_2090;
wire x_2091;
wire x_2092;
wire x_2093;
wire x_2094;
wire x_2095;
wire x_2096;
wire x_2097;
wire x_2098;
wire x_2099;
wire x_2100;
wire x_2101;
wire x_2102;
wire x_2103;
wire x_2104;
wire x_2105;
wire x_2106;
wire x_2107;
wire x_2108;
wire x_2109;
wire x_2110;
wire x_2111;
wire x_2112;
wire x_2113;
wire x_2114;
wire x_2115;
wire x_2116;
wire x_2117;
wire x_2118;
wire x_2119;
wire x_2120;
wire x_2121;
wire x_2122;
wire x_2123;
wire x_2124;
wire x_2125;
wire x_2126;
wire x_2127;
wire x_2128;
wire x_2129;
wire x_2130;
wire x_2131;
wire x_2132;
wire x_2133;
wire x_2134;
wire x_2135;
wire x_2136;
wire x_2137;
wire x_2138;
wire x_2139;
wire x_2140;
wire x_2141;
wire x_2142;
wire x_2143;
wire x_2144;
wire x_2145;
wire x_2146;
wire x_2147;
wire x_2148;
wire x_2149;
wire x_2150;
wire x_2151;
wire x_2152;
wire x_2153;
wire x_2154;
wire x_2155;
wire x_2156;
wire x_2157;
wire x_2158;
wire x_2159;
wire x_2160;
wire x_2161;
wire x_2162;
wire x_2163;
wire x_2164;
wire x_2165;
wire x_2166;
wire x_2167;
wire x_2168;
wire x_2169;
wire x_2170;
wire x_2171;
wire x_2172;
wire x_2173;
wire x_2174;
wire x_2175;
wire x_2176;
wire x_2177;
wire x_2178;
wire x_2179;
wire x_2180;
wire x_2181;
wire x_2182;
wire x_2183;
wire x_2184;
wire x_2185;
wire x_2186;
wire x_2187;
wire x_2188;
wire x_2189;
wire x_2190;
wire x_2191;
wire x_2192;
wire x_2193;
wire x_2194;
wire x_2195;
wire x_2196;
wire x_2197;
wire x_2198;
wire x_2199;
wire x_2200;
wire x_2201;
wire x_2202;
wire x_2203;
wire x_2204;
wire x_2205;
wire x_2206;
wire x_2207;
wire x_2208;
wire x_2209;
wire x_2210;
wire x_2211;
wire x_2212;
wire x_2213;
wire x_2214;
wire x_2215;
wire x_2216;
wire x_2217;
wire x_2218;
wire x_2219;
wire x_2220;
wire x_2221;
wire x_2222;
wire x_2223;
wire x_2224;
wire x_2225;
wire x_2226;
wire x_2227;
wire x_2228;
wire x_2229;
wire x_2230;
wire x_2231;
wire x_2232;
wire x_2233;
wire x_2234;
wire x_2235;
wire x_2236;
wire x_2237;
wire x_2238;
wire x_2239;
wire x_2240;
wire x_2241;
wire x_2242;
wire x_2243;
wire x_2244;
wire x_2245;
wire x_2246;
wire x_2247;
wire x_2248;
wire x_2249;
wire x_2250;
wire x_2251;
wire x_2252;
wire x_2253;
wire x_2254;
wire x_2255;
wire x_2256;
wire x_2257;
wire x_2258;
wire x_2259;
wire x_2260;
wire x_2261;
wire x_2262;
wire x_2263;
wire x_2264;
wire x_2265;
wire x_2266;
wire x_2267;
wire x_2268;
wire x_2269;
wire x_2270;
wire x_2271;
wire x_2272;
wire x_2273;
wire x_2274;
wire x_2275;
wire x_2276;
wire x_2277;
wire x_2278;
wire x_2279;
wire x_2280;
wire x_2281;
wire x_2282;
wire x_2283;
wire x_2284;
wire x_2285;
wire x_2286;
wire x_2287;
wire x_2288;
wire x_2289;
wire x_2290;
wire x_2291;
wire x_2292;
wire x_2293;
wire x_2294;
wire x_2295;
wire x_2296;
wire x_2297;
wire x_2298;
wire x_2299;
wire x_2300;
wire x_2301;
wire x_2302;
wire x_2303;
wire x_2304;
wire x_2305;
wire x_2306;
wire x_2307;
wire x_2308;
wire x_2309;
wire x_2310;
wire x_2311;
wire x_2312;
wire x_2313;
wire x_2314;
wire x_2315;
wire x_2316;
wire x_2317;
wire x_2318;
wire x_2319;
wire x_2320;
wire x_2321;
wire x_2322;
wire x_2323;
wire x_2324;
wire x_2325;
wire x_2326;
wire x_2327;
wire x_2328;
wire x_2329;
wire x_2330;
wire x_2331;
wire x_2332;
wire x_2333;
wire x_2334;
wire x_2335;
wire x_2336;
wire x_2337;
wire x_2338;
wire x_2339;
wire x_2340;
wire x_2341;
wire x_2342;
wire x_2343;
wire x_2344;
wire x_2345;
wire x_2346;
wire x_2347;
wire x_2348;
wire x_2349;
wire x_2350;
wire x_2351;
wire x_2352;
wire x_2353;
wire x_2354;
wire x_2355;
wire x_2356;
wire x_2357;
wire x_2358;
wire x_2359;
wire x_2360;
wire x_2361;
wire x_2362;
wire x_2363;
wire x_2364;
wire x_2365;
wire x_2366;
wire x_2367;
wire x_2368;
wire x_2369;
wire x_2370;
wire x_2371;
wire x_2372;
wire x_2373;
wire x_2374;
wire x_2375;
wire x_2376;
wire x_2377;
wire x_2378;
wire x_2379;
wire x_2380;
wire x_2381;
wire x_2382;
wire x_2383;
wire x_2384;
wire x_2385;
wire x_2386;
wire x_2387;
wire x_2388;
wire x_2389;
wire x_2390;
wire x_2391;
wire x_2392;
wire x_2393;
wire x_2394;
wire x_2395;
wire x_2396;
wire x_2397;
wire x_2398;
wire x_2399;
wire x_2400;
wire x_2401;
wire x_2402;
wire x_2403;
wire x_2404;
wire x_2405;
wire x_2406;
wire x_2407;
wire x_2408;
wire x_2409;
wire x_2410;
wire x_2411;
wire x_2412;
wire x_2413;
wire x_2414;
wire x_2415;
wire x_2416;
wire x_2417;
wire x_2418;
wire x_2419;
wire x_2420;
wire x_2421;
wire x_2422;
wire x_2423;
wire x_2424;
wire x_2425;
wire x_2426;
wire x_2427;
wire x_2428;
wire x_2429;
wire x_2430;
wire x_2431;
wire x_2432;
wire x_2433;
wire x_2434;
wire x_2435;
wire x_2436;
wire x_2437;
wire x_2438;
wire x_2439;
wire x_2440;
wire x_2441;
wire x_2442;
wire x_2443;
wire x_2444;
wire x_2445;
wire x_2446;
wire x_2447;
wire x_2448;
wire x_2449;
wire x_2450;
wire x_2451;
wire x_2452;
wire x_2453;
wire x_2454;
wire x_2455;
wire x_2456;
wire x_2457;
wire x_2458;
wire x_2459;
wire x_2460;
wire x_2461;
wire x_2462;
wire x_2463;
wire x_2464;
wire x_2465;
wire x_2466;
wire x_2467;
wire x_2468;
wire x_2469;
wire x_2470;
wire x_2471;
wire x_2472;
wire x_2473;
wire x_2474;
wire x_2475;
wire x_2476;
wire x_2477;
wire x_2478;
wire x_2479;
wire x_2480;
wire x_2481;
wire x_2482;
wire x_2483;
wire x_2484;
wire x_2485;
wire x_2486;
wire x_2487;
wire x_2488;
wire x_2489;
wire x_2490;
wire x_2491;
wire x_2492;
wire x_2493;
wire x_2494;
wire x_2495;
wire x_2496;
wire x_2497;
wire x_2498;
wire x_2499;
wire x_2500;
wire x_2501;
wire x_2502;
wire x_2503;
wire x_2504;
wire x_2505;
wire x_2506;
wire x_2507;
wire x_2508;
wire x_2509;
wire x_2510;
wire x_2511;
wire x_2512;
wire x_2513;
wire x_2514;
wire x_2515;
wire x_2516;
wire x_2517;
wire x_2518;
wire x_2519;
wire x_2520;
wire x_2521;
wire x_2522;
wire x_2523;
wire x_2524;
wire x_2525;
wire x_2526;
wire x_2527;
wire x_2528;
wire x_2529;
wire x_2530;
wire x_2531;
wire x_2532;
wire x_2533;
wire x_2534;
wire x_2535;
wire x_2536;
wire x_2537;
wire x_2538;
wire x_2539;
wire x_2540;
wire x_2541;
wire x_2542;
wire x_2543;
wire x_2544;
wire x_2545;
wire x_2546;
wire x_2547;
wire x_2548;
wire x_2549;
wire x_2550;
wire x_2551;
wire x_2552;
wire x_2553;
wire x_2554;
wire x_2555;
wire x_2556;
wire x_2557;
wire x_2558;
wire x_2559;
wire x_2560;
wire x_2561;
wire x_2562;
wire x_2563;
wire x_2564;
wire x_2565;
wire x_2566;
wire x_2567;
wire x_2568;
wire x_2569;
wire x_2570;
wire x_2571;
wire x_2572;
wire x_2573;
wire x_2574;
wire x_2575;
wire x_2576;
wire x_2577;
wire x_2578;
wire x_2579;
wire x_2580;
wire x_2581;
wire x_2582;
wire x_2583;
wire x_2584;
wire x_2585;
wire x_2586;
wire x_2587;
wire x_2588;
wire x_2589;
wire x_2590;
wire x_2591;
wire x_2592;
wire x_2593;
wire x_2594;
wire x_2595;
wire x_2596;
wire x_2597;
wire x_2598;
wire x_2599;
wire x_2600;
wire x_2601;
wire x_2602;
wire x_2603;
wire x_2604;
wire x_2605;
wire x_2606;
wire x_2607;
wire x_2608;
wire x_2609;
wire x_2610;
wire x_2611;
wire x_2612;
wire x_2613;
wire x_2614;
wire x_2615;
wire x_2616;
wire x_2617;
wire x_2618;
wire x_2619;
wire x_2620;
wire x_2621;
wire x_2622;
wire x_2623;
wire x_2624;
wire x_2625;
wire x_2626;
wire x_2627;
wire x_2628;
wire x_2629;
wire x_2630;
wire x_2631;
wire x_2632;
wire x_2633;
wire x_2634;
wire x_2635;
wire x_2636;
wire x_2637;
wire x_2638;
wire x_2639;
wire x_2640;
wire x_2641;
wire x_2642;
wire x_2643;
wire x_2644;
wire x_2645;
wire x_2646;
wire x_2647;
wire x_2648;
wire x_2649;
wire x_2650;
wire x_2651;
wire x_2652;
wire x_2653;
wire x_2654;
wire x_2655;
wire x_2656;
wire x_2657;
wire x_2658;
wire x_2659;
wire x_2660;
wire x_2661;
wire x_2662;
wire x_2663;
wire x_2664;
wire x_2665;
wire x_2666;
wire x_2667;
wire x_2668;
wire x_2669;
wire x_2670;
wire x_2671;
wire x_2672;
wire x_2673;
wire x_2674;
wire x_2675;
wire x_2676;
wire x_2677;
wire x_2678;
wire x_2679;
wire x_2680;
wire x_2681;
wire x_2682;
wire x_2683;
wire x_2684;
wire x_2685;
wire x_2686;
wire x_2687;
wire x_2688;
wire x_2689;
wire x_2690;
wire x_2691;
wire x_2692;
wire x_2693;
wire x_2694;
wire x_2695;
wire x_2696;
wire x_2697;
wire x_2698;
wire x_2699;
wire x_2700;
wire x_2701;
wire x_2702;
wire x_2703;
wire x_2704;
wire x_2705;
wire x_2706;
wire x_2707;
wire x_2708;
wire x_2709;
wire x_2710;
wire x_2711;
wire x_2712;
wire x_2713;
wire x_2714;
wire x_2715;
wire x_2716;
wire x_2717;
wire x_2718;
wire x_2719;
wire x_2720;
wire x_2721;
wire x_2722;
wire x_2723;
wire x_2724;
wire x_2725;
wire x_2726;
wire x_2727;
wire x_2728;
wire x_2729;
wire x_2730;
wire x_2731;
wire x_2732;
wire x_2733;
wire x_2734;
wire x_2735;
wire x_2736;
wire x_2737;
wire x_2738;
wire x_2739;
wire x_2740;
wire x_2741;
wire x_2742;
wire x_2743;
wire x_2744;
wire x_2745;
wire x_2746;
wire x_2747;
wire x_2748;
wire x_2749;
wire x_2750;
wire x_2751;
wire x_2752;
wire x_2753;
wire x_2754;
wire x_2755;
wire x_2756;
wire x_2757;
wire x_2758;
wire x_2759;
wire x_2760;
wire x_2761;
wire x_2762;
wire x_2763;
wire x_2764;
wire x_2765;
wire x_2766;
wire x_2767;
wire x_2768;
wire x_2769;
wire x_2770;
wire x_2771;
wire x_2772;
wire x_2773;
wire x_2774;
wire x_2775;
wire x_2776;
wire x_2777;
wire x_2778;
wire x_2779;
wire x_2780;
wire x_2781;
wire x_2782;
wire x_2783;
wire x_2784;
wire x_2785;
wire x_2786;
wire x_2787;
wire x_2788;
wire x_2789;
wire x_2790;
wire x_2791;
wire x_2792;
wire x_2793;
wire x_2794;
wire x_2795;
wire x_2796;
wire x_2797;
wire x_2798;
wire x_2799;
wire x_2800;
wire x_2801;
wire x_2802;
wire x_2803;
wire x_2804;
wire x_2805;
wire x_2806;
wire x_2807;
wire x_2808;
wire x_2809;
wire x_2810;
wire x_2811;
wire x_2812;
wire x_2813;
wire x_2814;
wire x_2815;
wire x_2816;
wire x_2817;
wire x_2818;
wire x_2819;
wire x_2820;
wire x_2821;
wire x_2822;
wire x_2823;
wire x_2824;
wire x_2825;
wire x_2826;
wire x_2827;
wire x_2828;
wire x_2829;
wire x_2830;
wire x_2831;
wire x_2832;
wire x_2833;
wire x_2834;
wire x_2835;
wire x_2836;
wire x_2837;
wire x_2838;
wire x_2839;
wire x_2840;
wire x_2841;
wire x_2842;
wire x_2843;
wire x_2844;
wire x_2845;
wire x_2846;
wire x_2847;
wire x_2848;
wire x_2849;
wire x_2850;
wire x_2851;
wire x_2852;
wire x_2853;
wire x_2854;
wire x_2855;
wire x_2856;
wire x_2857;
wire x_2858;
wire x_2859;
wire x_2860;
wire x_2861;
wire x_2862;
wire x_2863;
wire x_2864;
wire x_2865;
wire x_2866;
wire x_2867;
wire x_2868;
wire x_2869;
wire x_2870;
wire x_2871;
wire x_2872;
wire x_2873;
wire x_2874;
wire x_2875;
wire x_2876;
wire x_2877;
wire x_2878;
wire x_2879;
wire x_2880;
wire x_2881;
wire x_2882;
wire x_2883;
wire x_2884;
wire x_2885;
wire x_2886;
wire x_2887;
wire x_2888;
wire x_2889;
wire x_2890;
wire x_2891;
wire x_2892;
wire x_2893;
wire x_2894;
wire x_2895;
wire x_2896;
wire x_2897;
wire x_2898;
wire x_2899;
wire x_2900;
wire x_2901;
wire x_2902;
wire x_2903;
wire x_2904;
wire x_2905;
wire x_2906;
wire x_2907;
wire x_2908;
wire x_2909;
wire x_2910;
wire x_2911;
wire x_2912;
wire x_2913;
wire x_2914;
wire x_2915;
wire x_2916;
wire x_2917;
wire x_2918;
wire x_2919;
wire x_2920;
wire x_2921;
wire x_2922;
wire x_2923;
wire x_2924;
wire x_2925;
wire x_2926;
wire x_2927;
wire x_2928;
wire x_2929;
wire x_2930;
wire x_2931;
wire x_2932;
wire x_2933;
wire x_2934;
wire x_2935;
wire x_2936;
wire x_2937;
wire x_2938;
wire x_2939;
wire x_2940;
wire x_2941;
wire x_2942;
wire x_2943;
wire x_2944;
wire x_2945;
wire x_2946;
wire x_2947;
wire x_2948;
wire x_2949;
wire x_2950;
wire x_2951;
wire x_2952;
wire x_2953;
wire x_2954;
wire x_2955;
wire x_2956;
wire x_2957;
wire x_2958;
wire x_2959;
wire x_2960;
wire x_2961;
wire x_2962;
wire x_2963;
wire x_2964;
wire x_2965;
wire x_2966;
wire x_2967;
wire x_2968;
wire x_2969;
wire x_2970;
wire x_2971;
wire x_2972;
wire x_2973;
wire x_2974;
wire x_2975;
wire x_2976;
wire x_2977;
wire x_2978;
wire x_2979;
wire x_2980;
wire x_2981;
wire x_2982;
wire x_2983;
wire x_2984;
wire x_2985;
wire x_2986;
wire x_2987;
wire x_2988;
wire x_2989;
wire x_2990;
wire x_2991;
wire x_2992;
wire x_2993;
wire x_2994;
wire x_2995;
wire x_2996;
wire x_2997;
wire x_2998;
wire x_2999;
wire x_3000;
wire x_3001;
wire x_3002;
wire x_3003;
wire x_3004;
wire x_3005;
wire x_3006;
wire x_3007;
wire x_3008;
wire x_3009;
wire x_3010;
wire x_3011;
wire x_3012;
wire x_3013;
wire x_3014;
wire x_3015;
wire x_3016;
wire x_3017;
wire x_3018;
wire x_3019;
wire x_3020;
wire x_3021;
wire x_3022;
wire x_3023;
wire x_3024;
wire x_3025;
wire x_3026;
wire x_3027;
wire x_3028;
wire x_3029;
wire x_3030;
wire x_3031;
wire x_3032;
wire x_3033;
wire x_3034;
wire x_3035;
wire x_3036;
wire x_3037;
wire x_3038;
wire x_3039;
wire x_3040;
wire x_3041;
wire x_3042;
wire x_3043;
wire x_3044;
wire x_3045;
wire x_3046;
wire x_3047;
wire x_3048;
wire x_3049;
wire x_3050;
wire x_3051;
wire x_3052;
wire x_3053;
wire x_3054;
wire x_3055;
wire x_3056;
wire x_3057;
wire x_3058;
wire x_3059;
wire x_3060;
wire x_3061;
wire x_3062;
wire x_3063;
wire x_3064;
wire x_3065;
wire x_3066;
wire x_3067;
wire x_3068;
wire x_3069;
wire x_3070;
wire x_3071;
wire x_3072;
wire x_3073;
wire x_3074;
wire x_3075;
wire x_3076;
wire x_3077;
wire x_3078;
wire x_3079;
wire x_3080;
wire x_3081;
wire x_3082;
wire x_3083;
wire x_3084;
wire x_3085;
wire x_3086;
wire x_3087;
wire x_3088;
wire x_3089;
wire x_3090;
wire x_3091;
wire x_3092;
wire x_3093;
wire x_3094;
wire x_3095;
wire x_3096;
wire x_3097;
wire x_3098;
wire x_3099;
wire x_3100;
wire x_3101;
wire x_3102;
wire x_3103;
wire x_3104;
wire x_3105;
wire x_3106;
wire x_3107;
wire x_3108;
wire x_3109;
wire x_3110;
wire x_3111;
wire x_3112;
wire x_3113;
wire x_3114;
wire x_3115;
wire x_3116;
wire x_3117;
wire x_3118;
wire x_3119;
wire x_3120;
wire x_3121;
wire x_3122;
wire x_3123;
wire x_3124;
wire x_3125;
wire x_3126;
wire x_3127;
wire x_3128;
wire x_3129;
wire x_3130;
wire x_3131;
wire x_3132;
wire x_3133;
wire x_3134;
wire x_3135;
wire x_3136;
wire x_3137;
wire x_3138;
wire x_3139;
wire x_3140;
wire x_3141;
wire x_3142;
wire x_3143;
wire x_3144;
wire x_3145;
wire x_3146;
wire x_3147;
wire x_3148;
wire x_3149;
wire x_3150;
wire x_3151;
wire x_3152;
wire x_3153;
wire x_3154;
wire x_3155;
wire x_3156;
wire x_3157;
wire x_3158;
wire x_3159;
wire x_3160;
wire x_3161;
wire x_3162;
wire x_3163;
wire x_3164;
wire x_3165;
wire x_3166;
wire x_3167;
wire x_3168;
wire x_3169;
wire x_3170;
wire x_3171;
wire x_3172;
wire x_3173;
wire x_3174;
wire x_3175;
wire x_3176;
wire x_3177;
wire x_3178;
wire x_3179;
wire x_3180;
wire x_3181;
wire x_3182;
wire x_3183;
wire x_3184;
wire x_3185;
wire x_3186;
wire x_3187;
wire x_3188;
wire x_3189;
wire x_3190;
wire x_3191;
wire x_3192;
wire x_3193;
wire x_3194;
wire x_3195;
wire x_3196;
wire x_3197;
wire x_3198;
wire x_3199;
wire x_3200;
wire x_3201;
wire x_3202;
wire x_3203;
wire x_3204;
wire x_3205;
wire x_3206;
wire x_3207;
wire x_3208;
wire x_3209;
wire x_3210;
wire x_3211;
wire x_3212;
wire x_3213;
wire x_3214;
wire x_3215;
wire x_3216;
wire x_3217;
wire x_3218;
wire x_3219;
wire x_3220;
wire x_3221;
wire x_3222;
wire x_3223;
wire x_3224;
wire x_3225;
wire x_3226;
wire x_3227;
wire x_3228;
wire x_3229;
wire x_3230;
wire x_3231;
wire x_3232;
wire x_3233;
wire x_3234;
wire x_3235;
wire x_3236;
wire x_3237;
wire x_3238;
wire x_3239;
wire x_3240;
wire x_3241;
wire x_3242;
wire x_3243;
wire x_3244;
wire x_3245;
wire x_3246;
wire x_3247;
wire x_3248;
wire x_3249;
wire x_3250;
wire x_3251;
wire x_3252;
wire x_3253;
wire x_3254;
wire x_3255;
wire x_3256;
wire x_3257;
wire x_3258;
wire x_3259;
wire x_3260;
wire x_3261;
wire x_3262;
wire x_3263;
wire x_3264;
wire x_3265;
wire x_3266;
wire x_3267;
wire x_3268;
wire x_3269;
wire x_3270;
wire x_3271;
wire x_3272;
wire x_3273;
wire x_3274;
wire x_3275;
wire x_3276;
wire x_3277;
wire x_3278;
wire x_3279;
wire x_3280;
wire x_3281;
wire x_3282;
wire x_3283;
wire x_3284;
wire x_3285;
wire x_3286;
wire x_3287;
wire x_3288;
wire x_3289;
wire x_3290;
wire x_3291;
wire x_3292;
wire x_3293;
wire x_3294;
wire x_3295;
wire x_3296;
wire x_3297;
wire x_3298;
wire x_3299;
wire x_3300;
wire x_3301;
wire x_3302;
wire x_3303;
wire x_3304;
wire x_3305;
wire x_3306;
wire x_3307;
wire x_3308;
wire x_3309;
wire x_3310;
wire x_3311;
wire x_3312;
wire x_3313;
wire x_3314;
wire x_3315;
wire x_3316;
wire x_3317;
wire x_3318;
wire x_3319;
wire x_3320;
wire x_3321;
wire x_3322;
wire x_3323;
wire x_3324;
wire x_3325;
wire x_3326;
wire x_3327;
wire x_3328;
wire x_3329;
wire x_3330;
wire x_3331;
wire x_3332;
wire x_3333;
wire x_3334;
wire x_3335;
wire x_3336;
wire x_3337;
wire x_3338;
wire x_3339;
wire x_3340;
wire x_3341;
wire x_3342;
wire x_3343;
wire x_3344;
wire x_3345;
wire x_3346;
wire x_3347;
wire x_3348;
wire x_3349;
wire x_3350;
wire x_3351;
wire x_3352;
wire x_3353;
wire x_3354;
wire x_3355;
wire x_3356;
wire x_3357;
wire x_3358;
wire x_3359;
wire x_3360;
wire x_3361;
wire x_3362;
wire x_3363;
wire x_3364;
wire x_3365;
wire x_3366;
wire x_3367;
wire x_3368;
wire x_3369;
wire x_3370;
wire x_3371;
wire x_3372;
wire x_3373;
wire x_3374;
wire x_3375;
wire x_3376;
wire x_3377;
wire x_3378;
wire x_3379;
wire x_3380;
wire x_3381;
wire x_3382;
wire x_3383;
wire x_3384;
wire x_3385;
wire x_3386;
wire x_3387;
wire x_3388;
wire x_3389;
wire x_3390;
wire x_3391;
wire x_3392;
wire x_3393;
wire x_3394;
wire x_3395;
wire x_3396;
wire x_3397;
wire x_3398;
wire x_3399;
wire x_3400;
wire x_3401;
wire x_3402;
wire x_3403;
wire x_3404;
wire x_3405;
wire x_3406;
wire x_3407;
wire x_3408;
wire x_3409;
wire x_3410;
wire x_3411;
wire x_3412;
wire x_3413;
wire x_3414;
wire x_3415;
wire x_3416;
wire x_3417;
wire x_3418;
wire x_3419;
wire x_3420;
wire x_3421;
wire x_3422;
wire x_3423;
wire x_3424;
wire x_3425;
wire x_3426;
wire x_3427;
wire x_3428;
wire x_3429;
wire x_3430;
wire x_3431;
wire x_3432;
wire x_3433;
wire x_3434;
wire x_3435;
wire x_3436;
wire x_3437;
wire x_3438;
wire x_3439;
wire x_3440;
wire x_3441;
wire x_3442;
wire x_3443;
wire x_3444;
wire x_3445;
wire x_3446;
wire x_3447;
wire x_3448;
wire x_3449;
wire x_3450;
wire x_3451;
wire x_3452;
wire x_3453;
wire x_3454;
wire x_3455;
wire x_3456;
wire x_3457;
wire x_3458;
wire x_3459;
wire x_3460;
wire x_3461;
wire x_3462;
wire x_3463;
wire x_3464;
wire x_3465;
wire x_3466;
wire x_3467;
wire x_3468;
wire x_3469;
wire x_3470;
wire x_3471;
wire x_3472;
wire x_3473;
wire x_3474;
wire x_3475;
wire x_3476;
wire x_3477;
wire x_3478;
wire x_3479;
wire x_3480;
wire x_3481;
wire x_3482;
wire x_3483;
wire x_3484;
wire x_3485;
wire x_3486;
wire x_3487;
wire x_3488;
wire x_3489;
wire x_3490;
wire x_3491;
wire x_3492;
wire x_3493;
wire x_3494;
wire x_3495;
wire x_3496;
wire x_3497;
wire x_3498;
wire x_3499;
wire x_3500;
wire x_3501;
wire x_3502;
wire x_3503;
wire x_3504;
wire x_3505;
wire x_3506;
wire x_3507;
wire x_3508;
wire x_3509;
wire x_3510;
wire x_3511;
wire x_3512;
wire x_3513;
wire x_3514;
wire x_3515;
wire x_3516;
wire x_3517;
wire x_3518;
wire x_3519;
wire x_3520;
wire x_3521;
wire x_3522;
wire x_3523;
wire x_3524;
wire x_3525;
wire x_3526;
wire x_3527;
wire x_3528;
wire x_3529;
wire x_3530;
wire x_3531;
wire x_3532;
wire x_3533;
wire x_3534;
wire x_3535;
wire x_3536;
wire x_3537;
wire x_3538;
wire x_3539;
wire x_3540;
wire x_3541;
wire x_3542;
wire x_3543;
wire x_3544;
wire x_3545;
wire x_3546;
wire x_3547;
wire x_3548;
wire x_3549;
wire x_3550;
wire x_3551;
wire x_3552;
wire x_3553;
wire x_3554;
wire x_3555;
wire x_3556;
wire x_3557;
wire x_3558;
wire x_3559;
wire x_3560;
wire x_3561;
wire x_3562;
wire x_3563;
wire x_3564;
wire x_3565;
wire x_3566;
wire x_3567;
wire x_3568;
wire x_3569;
wire x_3570;
wire x_3571;
wire x_3572;
wire x_3573;
wire x_3574;
wire x_3575;
wire x_3576;
wire x_3577;
wire x_3578;
wire x_3579;
wire x_3580;
wire x_3581;
wire x_3582;
wire x_3583;
wire x_3584;
wire x_3585;
wire x_3586;
wire x_3587;
wire x_3588;
wire x_3589;
wire x_3590;
wire x_3591;
wire x_3592;
wire x_3593;
wire x_3594;
wire x_3595;
wire x_3596;
wire x_3597;
wire x_3598;
wire x_3599;
wire x_3600;
wire x_3601;
wire x_3602;
wire x_3603;
wire x_3604;
wire x_3605;
wire x_3606;
wire x_3607;
wire x_3608;
wire x_3609;
wire x_3610;
wire x_3611;
wire x_3612;
wire x_3613;
wire x_3614;
wire x_3615;
wire x_3616;
wire x_3617;
wire x_3618;
wire x_3619;
wire x_3620;
wire x_3621;
wire x_3622;
wire x_3623;
wire x_3624;
wire x_3625;
wire x_3626;
wire x_3627;
wire x_3628;
wire x_3629;
wire x_3630;
wire x_3631;
wire x_3632;
wire x_3633;
wire x_3634;
wire x_3635;
wire x_3636;
wire x_3637;
wire x_3638;
wire x_3639;
wire x_3640;
wire x_3641;
wire x_3642;
wire x_3643;
wire x_3644;
wire x_3645;
wire x_3646;
wire x_3647;
wire x_3648;
wire x_3649;
wire x_3650;
wire x_3651;
wire x_3652;
wire x_3653;
wire x_3654;
wire x_3655;
wire x_3656;
wire x_3657;
wire x_3658;
wire x_3659;
wire x_3660;
wire x_3661;
wire x_3662;
wire x_3663;
wire x_3664;
wire x_3665;
wire x_3666;
wire x_3667;
wire x_3668;
wire x_3669;
wire x_3670;
wire x_3671;
wire x_3672;
wire x_3673;
wire x_3674;
wire x_3675;
wire x_3676;
wire x_3677;
wire x_3678;
wire x_3679;
wire x_3680;
wire x_3681;
wire x_3682;
wire x_3683;
wire x_3684;
wire x_3685;
wire x_3686;
wire x_3687;
wire x_3688;
wire x_3689;
wire x_3690;
wire x_3691;
wire x_3692;
wire x_3693;
wire x_3694;
wire x_3695;
wire x_3696;
wire x_3697;
wire x_3698;
wire x_3699;
wire x_3700;
wire x_3701;
wire x_3702;
wire x_3703;
wire x_3704;
wire x_3705;
wire x_3706;
wire x_3707;
wire x_3708;
wire x_3709;
wire x_3710;
wire x_3711;
wire x_3712;
wire x_3713;
wire x_3714;
wire x_3715;
wire x_3716;
wire x_3717;
wire x_3718;
wire x_3719;
wire x_3720;
wire x_3721;
wire x_3722;
wire x_3723;
wire x_3724;
wire x_3725;
wire x_3726;
wire x_3727;
wire x_3728;
wire x_3729;
wire x_3730;
wire x_3731;
wire x_3732;
wire x_3733;
wire x_3734;
wire x_3735;
wire x_3736;
wire x_3737;
wire x_3738;
wire x_3739;
wire x_3740;
wire x_3741;
wire x_3742;
wire x_3743;
wire x_3744;
wire x_3745;
wire x_3746;
wire x_3747;
wire x_3748;
wire x_3749;
wire x_3750;
wire x_3751;
wire x_3752;
wire x_3753;
wire x_3754;
wire x_3755;
wire x_3756;
wire x_3757;
wire x_3758;
wire x_3759;
wire x_3760;
wire x_3761;
wire x_3762;
wire x_3763;
wire x_3764;
wire x_3765;
wire x_3766;
wire x_3767;
wire x_3768;
wire x_3769;
wire x_3770;
wire x_3771;
wire x_3772;
wire x_3773;
wire x_3774;
wire x_3775;
wire x_3776;
wire x_3777;
wire x_3778;
wire x_3779;
wire x_3780;
wire x_3781;
wire x_3782;
wire x_3783;
wire x_3784;
wire x_3785;
wire x_3786;
wire x_3787;
wire x_3788;
wire x_3789;
wire x_3790;
wire x_3791;
wire x_3792;
wire x_3793;
wire x_3794;
wire x_3795;
wire x_3796;
wire x_3797;
wire x_3798;
wire x_3799;
wire x_3800;
wire x_3801;
wire x_3802;
wire x_3803;
wire x_3804;
wire x_3805;
wire x_3806;
wire x_3807;
wire x_3808;
wire x_3809;
wire x_3810;
wire x_3811;
wire x_3812;
wire x_3813;
wire x_3814;
wire x_3815;
wire x_3816;
wire x_3817;
wire x_3818;
wire x_3819;
wire x_3820;
wire x_3821;
wire x_3822;
wire x_3823;
wire x_3824;
wire x_3825;
wire x_3826;
wire x_3827;
wire x_3828;
wire x_3829;
wire x_3830;
wire x_3831;
wire x_3832;
wire x_3833;
wire x_3834;
wire x_3835;
wire x_3836;
wire x_3837;
wire x_3838;
wire x_3839;
wire x_3840;
wire x_3841;
wire x_3842;
wire x_3843;
wire x_3844;
wire x_3845;
wire x_3846;
wire x_3847;
wire x_3848;
wire x_3849;
wire x_3850;
wire x_3851;
wire x_3852;
wire x_3853;
wire x_3854;
wire x_3855;
wire x_3856;
wire x_3857;
wire x_3858;
wire x_3859;
wire x_3860;
wire x_3861;
wire x_3862;
wire x_3863;
wire x_3864;
wire x_3865;
wire x_3866;
wire x_3867;
wire x_3868;
wire x_3869;
wire x_3870;
wire x_3871;
wire x_3872;
wire x_3873;
wire x_3874;
wire x_3875;
wire x_3876;
wire x_3877;
wire x_3878;
wire x_3879;
wire x_3880;
wire x_3881;
wire x_3882;
wire x_3883;
wire x_3884;
wire x_3885;
wire x_3886;
wire x_3887;
wire x_3888;
wire x_3889;
wire x_3890;
wire x_3891;
wire x_3892;
wire x_3893;
wire x_3894;
wire x_3895;
wire x_3896;
wire x_3897;
wire x_3898;
wire x_3899;
wire x_3900;
wire x_3901;
wire x_3902;
wire x_3903;
wire x_3904;
wire x_3905;
wire x_3906;
wire x_3907;
wire x_3908;
wire x_3909;
wire x_3910;
wire x_3911;
wire x_3912;
wire x_3913;
wire x_3914;
wire x_3915;
wire x_3916;
wire x_3917;
wire x_3918;
wire x_3919;
wire x_3920;
wire x_3921;
wire x_3922;
wire x_3923;
wire x_3924;
wire x_3925;
wire x_3926;
wire x_3927;
wire x_3928;
wire x_3929;
wire x_3930;
wire x_3931;
wire x_3932;
wire x_3933;
wire x_3934;
wire x_3935;
wire x_3936;
wire x_3937;
wire x_3938;
wire x_3939;
wire x_3940;
wire x_3941;
wire x_3942;
wire x_3943;
wire x_3944;
wire x_3945;
wire x_3946;
wire x_3947;
wire x_3948;
wire x_3949;
wire x_3950;
wire x_3951;
wire x_3952;
wire x_3953;
wire x_3954;
wire x_3955;
wire x_3956;
wire x_3957;
wire x_3958;
wire x_3959;
wire x_3960;
wire x_3961;
wire x_3962;
wire x_3963;
wire x_3964;
wire x_3965;
wire x_3966;
wire x_3967;
wire x_3968;
wire x_3969;
wire x_3970;
wire x_3971;
wire x_3972;
wire x_3973;
wire x_3974;
wire x_3975;
wire x_3976;
wire x_3977;
wire x_3978;
wire x_3979;
wire x_3980;
wire x_3981;
wire x_3982;
wire x_3983;
wire x_3984;
wire x_3985;
wire x_3986;
wire x_3987;
wire x_3988;
wire x_3989;
wire x_3990;
wire x_3991;
wire x_3992;
wire x_3993;
wire x_3994;
wire x_3995;
wire x_3996;
wire x_3997;
wire x_3998;
wire x_3999;
wire x_4000;
wire x_4001;
wire x_4002;
wire x_4003;
wire x_4004;
wire x_4005;
wire x_4006;
wire x_4007;
wire x_4008;
wire x_4009;
wire x_4010;
wire x_4011;
wire x_4012;
wire x_4013;
wire x_4014;
wire x_4015;
wire x_4016;
wire x_4017;
wire x_4018;
wire x_4019;
wire x_4020;
wire x_4021;
wire x_4022;
wire x_4023;
wire x_4024;
wire x_4025;
wire x_4026;
wire x_4027;
wire x_4028;
wire x_4029;
wire x_4030;
wire x_4031;
wire x_4032;
wire x_4033;
wire x_4034;
wire x_4035;
wire x_4036;
wire x_4037;
wire x_4038;
wire x_4039;
wire x_4040;
wire x_4041;
wire x_4042;
wire x_4043;
wire x_4044;
wire x_4045;
wire x_4046;
wire x_4047;
wire x_4048;
wire x_4049;
wire x_4050;
wire x_4051;
wire x_4052;
wire x_4053;
wire x_4054;
wire x_4055;
wire x_4056;
wire x_4057;
wire x_4058;
wire x_4059;
wire x_4060;
wire x_4061;
wire x_4062;
wire x_4063;
wire x_4064;
wire x_4065;
wire x_4066;
wire x_4067;
wire x_4068;
wire x_4069;
wire x_4070;
wire x_4071;
wire x_4072;
wire x_4073;
wire x_4074;
wire x_4075;
wire x_4076;
wire x_4077;
wire x_4078;
wire x_4079;
wire x_4080;
wire x_4081;
wire x_4082;
wire x_4083;
wire x_4084;
wire x_4085;
wire x_4086;
wire x_4087;
wire x_4088;
wire x_4089;
wire x_4090;
wire x_4091;
wire x_4092;
wire x_4093;
wire x_4094;
wire x_4095;
wire x_4096;
wire x_4097;
wire x_4098;
wire x_4099;
wire x_4100;
wire x_4101;
wire x_4102;
wire x_4103;
wire x_4104;
wire x_4105;
wire x_4106;
wire x_4107;
wire x_4108;
wire x_4109;
wire x_4110;
wire x_4111;
wire x_4112;
wire x_4113;
wire x_4114;
wire x_4115;
wire x_4116;
wire x_4117;
wire x_4118;
wire x_4119;
wire x_4120;
wire x_4121;
wire x_4122;
wire x_4123;
wire x_4124;
wire x_4125;
wire x_4126;
wire x_4127;
wire x_4128;
wire x_4129;
wire x_4130;
wire x_4131;
wire x_4132;
wire x_4133;
wire x_4134;
wire x_4135;
wire x_4136;
wire x_4137;
wire x_4138;
wire x_4139;
wire x_4140;
wire x_4141;
wire x_4142;
wire x_4143;
wire x_4144;
wire x_4145;
wire x_4146;
wire x_4147;
wire x_4148;
wire x_4149;
wire x_4150;
wire x_4151;
wire x_4152;
wire x_4153;
wire x_4154;
wire x_4155;
wire x_4156;
wire x_4157;
wire x_4158;
wire x_4159;
wire x_4160;
wire x_4161;
wire x_4162;
wire x_4163;
wire x_4164;
wire x_4165;
wire x_4166;
wire x_4167;
wire x_4168;
wire x_4169;
wire x_4170;
wire x_4171;
wire x_4172;
wire x_4173;
wire x_4174;
wire x_4175;
wire x_4176;
wire x_4177;
wire x_4178;
wire x_4179;
wire x_4180;
wire x_4181;
wire x_4182;
wire x_4183;
wire x_4184;
wire x_4185;
wire x_4186;
wire x_4187;
wire x_4188;
wire x_4189;
wire x_4190;
wire x_4191;
wire x_4192;
wire x_4193;
wire x_4194;
wire x_4195;
wire x_4196;
wire x_4197;
wire x_4198;
wire x_4199;
wire x_4200;
wire x_4201;
wire x_4202;
wire x_4203;
wire x_4204;
wire x_4205;
wire x_4206;
wire x_4207;
wire x_4208;
wire x_4209;
wire x_4210;
wire x_4211;
wire x_4212;
wire x_4213;
wire x_4214;
wire x_4215;
wire x_4216;
wire x_4217;
wire x_4218;
wire x_4219;
wire x_4220;
wire x_4221;
wire x_4222;
wire x_4223;
wire x_4224;
wire x_4225;
wire x_4226;
wire x_4227;
wire x_4228;
wire x_4229;
wire x_4230;
wire x_4231;
wire x_4232;
wire x_4233;
wire x_4234;
wire x_4235;
wire x_4236;
wire x_4237;
wire x_4238;
wire x_4239;
wire x_4240;
wire x_4241;
wire x_4242;
wire x_4243;
wire x_4244;
wire x_4245;
wire x_4246;
wire x_4247;
wire x_4248;
wire x_4249;
wire x_4250;
wire x_4251;
wire x_4252;
wire x_4253;
wire x_4254;
wire x_4255;
wire x_4256;
wire x_4257;
wire x_4258;
wire x_4259;
wire x_4260;
wire x_4261;
wire x_4262;
wire x_4263;
wire x_4264;
wire x_4265;
wire x_4266;
wire x_4267;
wire x_4268;
wire x_4269;
wire x_4270;
wire x_4271;
wire x_4272;
wire x_4273;
wire x_4274;
wire x_4275;
wire x_4276;
wire x_4277;
wire x_4278;
wire x_4279;
wire x_4280;
wire x_4281;
wire x_4282;
wire x_4283;
wire x_4284;
wire x_4285;
wire x_4286;
wire x_4287;
wire x_4288;
wire x_4289;
wire x_4290;
wire x_4291;
wire x_4292;
wire x_4293;
wire x_4294;
wire x_4295;
wire x_4296;
wire x_4297;
wire x_4298;
wire x_4299;
wire x_4300;
wire x_4301;
wire x_4302;
wire x_4303;
wire x_4304;
wire x_4305;
wire x_4306;
wire x_4307;
wire x_4308;
wire x_4309;
wire x_4310;
wire x_4311;
wire x_4312;
wire x_4313;
wire x_4314;
wire x_4315;
wire x_4316;
wire x_4317;
wire x_4318;
wire x_4319;
wire x_4320;
wire x_4321;
wire x_4322;
wire x_4323;
wire x_4324;
wire x_4325;
wire x_4326;
wire x_4327;
wire x_4328;
wire x_4329;
wire x_4330;
wire x_4331;
wire x_4332;
wire x_4333;
wire x_4334;
wire x_4335;
wire x_4336;
wire x_4337;
wire x_4338;
wire x_4339;
wire x_4340;
wire x_4341;
wire x_4342;
wire x_4343;
wire x_4344;
wire x_4345;
wire x_4346;
wire x_4347;
wire x_4348;
wire x_4349;
wire x_4350;
wire x_4351;
wire x_4352;
wire x_4353;
wire x_4354;
wire x_4355;
wire x_4356;
wire x_4357;
wire x_4358;
wire x_4359;
wire x_4360;
wire x_4361;
wire x_4362;
wire x_4363;
wire x_4364;
wire x_4365;
wire x_4366;
wire x_4367;
wire x_4368;
wire x_4369;
wire x_4370;
wire x_4371;
wire x_4372;
wire x_4373;
wire x_4374;
wire x_4375;
wire x_4376;
wire x_4377;
wire x_4378;
wire x_4379;
wire x_4380;
wire x_4381;
wire x_4382;
wire x_4383;
wire x_4384;
wire x_4385;
wire x_4386;
wire x_4387;
wire x_4388;
wire x_4389;
wire x_4390;
wire x_4391;
wire x_4392;
wire x_4393;
wire x_4394;
wire x_4395;
wire x_4396;
wire x_4397;
wire x_4398;
wire x_4399;
wire x_4400;
wire x_4401;
wire x_4402;
wire x_4403;
wire x_4404;
wire x_4405;
wire x_4406;
wire x_4407;
wire x_4408;
wire x_4409;
wire x_4410;
wire x_4411;
wire x_4412;
wire x_4413;
wire x_4414;
wire x_4415;
wire x_4416;
wire x_4417;
wire x_4418;
wire x_4419;
wire x_4420;
wire x_4421;
wire x_4422;
wire x_4423;
wire x_4424;
wire x_4425;
wire x_4426;
wire x_4427;
wire x_4428;
wire x_4429;
wire x_4430;
wire x_4431;
wire x_4432;
wire x_4433;
wire x_4434;
wire x_4435;
wire x_4436;
wire x_4437;
wire x_4438;
wire x_4439;
wire x_4440;
wire x_4441;
wire x_4442;
wire x_4443;
wire x_4444;
wire x_4445;
wire x_4446;
wire x_4447;
wire x_4448;
wire x_4449;
wire x_4450;
wire x_4451;
wire x_4452;
wire x_4453;
wire x_4454;
wire x_4455;
wire x_4456;
wire x_4457;
wire x_4458;
wire x_4459;
wire x_4460;
wire x_4461;
wire x_4462;
wire x_4463;
wire x_4464;
wire x_4465;
wire x_4466;
wire x_4467;
wire x_4468;
wire x_4469;
wire x_4470;
wire x_4471;
wire x_4472;
wire x_4473;
wire x_4474;
wire x_4475;
wire x_4476;
wire x_4477;
wire x_4478;
wire x_4479;
wire x_4480;
wire x_4481;
wire x_4482;
wire x_4483;
wire x_4484;
wire x_4485;
wire x_4486;
wire x_4487;
wire x_4488;
wire x_4489;
wire x_4490;
wire x_4491;
wire x_4492;
wire x_4493;
wire x_4494;
wire x_4495;
wire x_4496;
wire x_4497;
wire x_4498;
wire x_4499;
wire x_4500;
wire x_4501;
wire x_4502;
wire x_4503;
wire x_4504;
wire x_4505;
wire x_4506;
wire x_4507;
wire x_4508;
wire x_4509;
wire x_4510;
wire x_4511;
wire x_4512;
wire x_4513;
wire x_4514;
wire x_4515;
wire x_4516;
wire x_4517;
wire x_4518;
wire x_4519;
wire x_4520;
wire x_4521;
wire x_4522;
wire x_4523;
wire x_4524;
wire x_4525;
wire x_4526;
wire x_4527;
wire x_4528;
wire x_4529;
wire x_4530;
wire x_4531;
wire x_4532;
wire x_4533;
wire x_4534;
wire x_4535;
wire x_4536;
wire x_4537;
wire x_4538;
wire x_4539;
wire x_4540;
wire x_4541;
wire x_4542;
wire x_4543;
wire x_4544;
wire x_4545;
wire x_4546;
wire x_4547;
wire x_4548;
wire x_4549;
wire x_4550;
wire x_4551;
wire x_4552;
wire x_4553;
wire x_4554;
wire x_4555;
wire x_4556;
wire x_4557;
wire x_4558;
wire x_4559;
wire x_4560;
wire x_4561;
wire x_4562;
wire x_4563;
wire x_4564;
wire x_4565;
wire x_4566;
wire x_4567;
wire x_4568;
wire x_4569;
wire x_4570;
wire x_4571;
wire x_4572;
wire x_4573;
wire x_4574;
wire x_4575;
wire x_4576;
wire x_4577;
wire x_4578;
wire x_4579;
wire x_4580;
wire x_4581;
wire x_4582;
wire x_4583;
wire x_4584;
wire x_4585;
wire x_4586;
wire x_4587;
wire x_4588;
wire x_4589;
wire x_4590;
wire x_4591;
wire x_4592;
wire x_4593;
wire x_4594;
wire x_4595;
wire x_4596;
wire x_4597;
wire x_4598;
wire x_4599;
wire x_4600;
wire x_4601;
wire x_4602;
wire x_4603;
wire x_4604;
wire x_4605;
wire x_4606;
wire x_4607;
wire x_4608;
wire x_4609;
wire x_4610;
wire x_4611;
wire x_4612;
wire x_4613;
wire x_4614;
wire x_4615;
wire x_4616;
wire x_4617;
wire x_4618;
wire x_4619;
wire x_4620;
wire x_4621;
wire x_4622;
wire x_4623;
wire x_4624;
wire x_4625;
wire x_4626;
wire x_4627;
wire x_4628;
wire x_4629;
wire x_4630;
wire x_4631;
wire x_4632;
wire x_4633;
wire x_4634;
wire x_4635;
wire x_4636;
wire x_4637;
wire x_4638;
wire x_4639;
wire x_4640;
wire x_4641;
wire x_4642;
wire x_4643;
wire x_4644;
wire x_4645;
wire x_4646;
wire x_4647;
wire x_4648;
wire x_4649;
wire x_4650;
wire x_4651;
wire x_4652;
wire x_4653;
wire x_4654;
wire x_4655;
wire x_4656;
wire x_4657;
wire x_4658;
wire x_4659;
wire x_4660;
wire x_4661;
wire x_4662;
wire x_4663;
wire x_4664;
wire x_4665;
wire x_4666;
wire x_4667;
wire x_4668;
wire x_4669;
wire x_4670;
wire x_4671;
wire x_4672;
wire x_4673;
wire x_4674;
wire x_4675;
wire x_4676;
wire x_4677;
wire x_4678;
wire x_4679;
wire x_4680;
wire x_4681;
wire x_4682;
wire x_4683;
wire x_4684;
wire x_4685;
wire x_4686;
wire x_4687;
wire x_4688;
wire x_4689;
wire x_4690;
wire x_4691;
wire x_4692;
wire x_4693;
wire x_4694;
wire x_4695;
wire x_4696;
wire x_4697;
wire x_4698;
wire x_4699;
wire x_4700;
wire x_4701;
wire x_4702;
wire x_4703;
wire x_4704;
wire x_4705;
wire x_4706;
wire x_4707;
wire x_4708;
wire x_4709;
wire x_4710;
wire x_4711;
wire x_4712;
wire x_4713;
wire x_4714;
wire x_4715;
wire x_4716;
wire x_4717;
wire x_4718;
wire x_4719;
wire x_4720;
wire x_4721;
wire x_4722;
wire x_4723;
wire x_4724;
wire x_4725;
wire x_4726;
wire x_4727;
wire x_4728;
wire x_4729;
wire x_4730;
wire x_4731;
wire x_4732;
wire x_4733;
wire x_4734;
wire x_4735;
wire x_4736;
wire x_4737;
wire x_4738;
wire x_4739;
wire x_4740;
wire x_4741;
wire x_4742;
wire x_4743;
wire x_4744;
wire x_4745;
wire x_4746;
wire x_4747;
wire x_4748;
wire x_4749;
wire x_4750;
wire x_4751;
wire x_4752;
wire x_4753;
wire x_4754;
wire x_4755;
wire x_4756;
wire x_4757;
wire x_4758;
wire x_4759;
wire x_4760;
wire x_4761;
wire x_4762;
wire x_4763;
wire x_4764;
wire x_4765;
wire x_4766;
wire x_4767;
wire x_4768;
wire x_4769;
wire x_4770;
wire x_4771;
wire x_4772;
wire x_4773;
wire x_4774;
wire x_4775;
wire x_4776;
wire x_4777;
wire x_4778;
wire x_4779;
wire x_4780;
wire x_4781;
wire x_4782;
wire x_4783;
wire x_4784;
wire x_4785;
wire x_4786;
wire x_4787;
wire x_4788;
wire x_4789;
wire x_4790;
wire x_4791;
wire x_4792;
wire x_4793;
wire x_4794;
wire x_4795;
wire x_4796;
wire x_4797;
wire x_4798;
wire x_4799;
wire x_4800;
wire x_4801;
wire x_4802;
wire x_4803;
wire x_4804;
wire x_4805;
wire x_4806;
wire x_4807;
wire x_4808;
wire x_4809;
wire x_4810;
wire x_4811;
wire x_4812;
wire x_4813;
wire x_4814;
wire x_4815;
wire x_4816;
wire x_4817;
wire x_4818;
wire x_4819;
wire x_4820;
wire x_4821;
wire x_4822;
wire x_4823;
wire x_4824;
wire x_4825;
wire x_4826;
wire x_4827;
wire x_4828;
wire x_4829;
wire x_4830;
wire x_4831;
wire x_4832;
wire x_4833;
wire x_4834;
wire x_4835;
wire x_4836;
wire x_4837;
wire x_4838;
wire x_4839;
wire x_4840;
wire x_4841;
wire x_4842;
wire x_4843;
wire x_4844;
wire x_4845;
wire x_4846;
wire x_4847;
wire x_4848;
wire x_4849;
wire x_4850;
wire x_4851;
wire x_4852;
wire x_4853;
wire x_4854;
wire x_4855;
wire x_4856;
wire x_4857;
wire x_4858;
wire x_4859;
wire x_4860;
wire x_4861;
wire x_4862;
wire x_4863;
wire x_4864;
wire x_4865;
wire x_4866;
wire x_4867;
wire x_4868;
wire x_4869;
wire x_4870;
wire x_4871;
wire x_4872;
wire x_4873;
wire x_4874;
wire x_4875;
wire x_4876;
wire x_4877;
wire x_4878;
wire x_4879;
wire x_4880;
wire x_4881;
wire x_4882;
wire x_4883;
wire x_4884;
wire x_4885;
wire x_4886;
wire x_4887;
wire x_4888;
wire x_4889;
wire x_4890;
wire x_4891;
wire x_4892;
wire x_4893;
wire x_4894;
wire x_4895;
wire x_4896;
wire x_4897;
wire x_4898;
wire x_4899;
wire x_4900;
wire x_4901;
wire x_4902;
wire x_4903;
wire x_4904;
wire x_4905;
wire x_4906;
wire x_4907;
wire x_4908;
wire x_4909;
wire x_4910;
wire x_4911;
wire x_4912;
wire x_4913;
wire x_4914;
wire x_4915;
wire x_4916;
wire x_4917;
wire x_4918;
wire x_4919;
wire x_4920;
wire x_4921;
wire x_4922;
wire x_4923;
wire x_4924;
wire x_4925;
wire x_4926;
wire x_4927;
wire x_4928;
wire x_4929;
wire x_4930;
wire x_4931;
wire x_4932;
wire x_4933;
wire x_4934;
wire x_4935;
wire x_4936;
wire x_4937;
wire x_4938;
wire x_4939;
wire x_4940;
wire x_4941;
wire x_4942;
wire x_4943;
wire x_4944;
wire x_4945;
wire x_4946;
wire x_4947;
wire x_4948;
wire x_4949;
wire x_4950;
wire x_4951;
wire x_4952;
wire x_4953;
wire x_4954;
wire x_4955;
wire x_4956;
wire x_4957;
wire x_4958;
wire x_4959;
wire x_4960;
wire x_4961;
wire x_4962;
wire x_4963;
wire x_4964;
wire x_4965;
wire x_4966;
wire x_4967;
wire x_4968;
wire x_4969;
wire x_4970;
wire x_4971;
wire x_4972;
wire x_4973;
wire x_4974;
wire x_4975;
wire x_4976;
wire x_4977;
wire x_4978;
wire x_4979;
wire x_4980;
wire x_4981;
wire x_4982;
wire x_4983;
wire x_4984;
wire x_4985;
wire x_4986;
wire x_4987;
wire x_4988;
wire x_4989;
wire x_4990;
wire x_4991;
wire x_4992;
wire x_4993;
wire x_4994;
wire x_4995;
wire x_4996;
wire x_4997;
wire x_4998;
wire x_4999;
wire x_5000;
wire x_5001;
wire x_5002;
wire x_5003;
wire x_5004;
wire x_5005;
wire x_5006;
wire x_5007;
wire x_5008;
wire x_5009;
wire x_5010;
wire x_5011;
wire x_5012;
wire x_5013;
wire x_5014;
wire x_5015;
wire x_5016;
wire x_5017;
wire x_5018;
wire x_5019;
wire x_5020;
wire x_5021;
wire x_5022;
wire x_5023;
wire x_5024;
wire x_5025;
wire x_5026;
wire x_5027;
wire x_5028;
wire x_5029;
wire x_5030;
wire x_5031;
wire x_5032;
wire x_5033;
wire x_5034;
wire x_5035;
wire x_5036;
wire x_5037;
wire x_5038;
wire x_5039;
wire x_5040;
wire x_5041;
wire x_5042;
wire x_5043;
wire x_5044;
wire x_5045;
wire x_5046;
wire x_5047;
wire x_5048;
wire x_5049;
wire x_5050;
wire x_5051;
wire x_5052;
wire x_5053;
wire x_5054;
wire x_5055;
wire x_5056;
wire x_5057;
wire x_5058;
wire x_5059;
wire x_5060;
wire x_5061;
wire x_5062;
wire x_5063;
wire x_5064;
wire x_5065;
wire x_5066;
wire x_5067;
wire x_5068;
wire x_5069;
wire x_5070;
wire x_5071;
wire x_5072;
wire x_5073;
wire x_5074;
wire x_5075;
wire x_5076;
wire x_5077;
wire x_5078;
wire x_5079;
wire x_5080;
wire x_5081;
wire x_5082;
wire x_5083;
wire x_5084;
wire x_5085;
wire x_5086;
wire x_5087;
wire x_5088;
wire x_5089;
wire x_5090;
wire x_5091;
wire x_5092;
wire x_5093;
wire x_5094;
wire x_5095;
wire x_5096;
wire x_5097;
wire x_5098;
wire x_5099;
wire x_5100;
wire x_5101;
wire x_5102;
wire x_5103;
wire x_5104;
wire x_5105;
wire x_5106;
wire x_5107;
wire x_5108;
wire x_5109;
wire x_5110;
wire x_5111;
wire x_5112;
wire x_5113;
wire x_5114;
wire x_5115;
wire x_5116;
wire x_5117;
wire x_5118;
wire x_5119;
wire x_5120;
wire x_5121;
wire x_5122;
wire x_5123;
wire x_5124;
wire x_5125;
wire x_5126;
wire x_5127;
wire x_5128;
wire x_5129;
wire x_5130;
wire x_5131;
wire x_5132;
wire x_5133;
wire x_5134;
wire x_5135;
wire x_5136;
wire x_5137;
wire x_5138;
wire x_5139;
wire x_5140;
wire x_5141;
wire x_5142;
wire x_5143;
wire x_5144;
wire x_5145;
wire x_5146;
wire x_5147;
wire x_5148;
wire x_5149;
wire x_5150;
wire x_5151;
wire x_5152;
wire x_5153;
wire x_5154;
wire x_5155;
wire x_5156;
wire x_5157;
wire x_5158;
wire x_5159;
wire x_5160;
wire x_5161;
wire x_5162;
wire x_5163;
wire x_5164;
wire x_5165;
wire x_5166;
wire x_5167;
wire x_5168;
wire x_5169;
wire x_5170;
wire x_5171;
wire x_5172;
wire x_5173;
wire x_5174;
wire x_5175;
wire x_5176;
wire x_5177;
wire x_5178;
wire x_5179;
wire x_5180;
wire x_5181;
wire x_5182;
wire x_5183;
wire x_5184;
wire x_5185;
wire x_5186;
wire x_5187;
wire x_5188;
wire x_5189;
wire x_5190;
wire x_5191;
wire x_5192;
wire x_5193;
wire x_5194;
wire x_5195;
wire x_5196;
wire x_5197;
wire x_5198;
wire x_5199;
wire x_5200;
wire x_5201;
wire x_5202;
wire x_5203;
wire x_5204;
wire x_5205;
wire x_5206;
wire x_5207;
wire x_5208;
wire x_5209;
wire x_5210;
wire x_5211;
wire x_5212;
wire x_5213;
wire x_5214;
wire x_5215;
wire x_5216;
wire x_5217;
wire x_5218;
wire x_5219;
wire x_5220;
wire x_5221;
wire x_5222;
wire x_5223;
wire x_5224;
wire x_5225;
wire x_5226;
wire x_5227;
wire x_5228;
wire x_5229;
wire x_5230;
wire x_5231;
wire x_5232;
wire x_5233;
wire x_5234;
wire x_5235;
wire x_5236;
wire x_5237;
wire x_5238;
wire x_5239;
wire x_5240;
wire x_5241;
wire x_5242;
wire x_5243;
wire x_5244;
wire x_5245;
wire x_5246;
wire x_5247;
wire x_5248;
wire x_5249;
wire x_5250;
wire x_5251;
wire x_5252;
wire x_5253;
wire x_5254;
wire x_5255;
wire x_5256;
wire x_5257;
wire x_5258;
wire x_5259;
wire x_5260;
wire x_5261;
wire x_5262;
wire x_5263;
wire x_5264;
wire x_5265;
wire x_5266;
wire x_5267;
wire x_5268;
wire x_5269;
wire x_5270;
wire x_5271;
wire x_5272;
wire x_5273;
wire x_5274;
wire x_5275;
wire x_5276;
wire x_5277;
wire x_5278;
wire x_5279;
wire x_5280;
wire x_5281;
wire x_5282;
wire x_5283;
wire x_5284;
wire x_5285;
wire x_5286;
wire x_5287;
wire x_5288;
wire x_5289;
wire x_5290;
wire x_5291;
wire x_5292;
wire x_5293;
wire x_5294;
wire x_5295;
wire x_5296;
wire x_5297;
wire x_5298;
wire x_5299;
wire x_5300;
wire x_5301;
wire x_5302;
wire x_5303;
wire x_5304;
wire x_5305;
wire x_5306;
wire x_5307;
wire x_5308;
wire x_5309;
wire x_5310;
wire x_5311;
wire x_5312;
wire x_5313;
wire x_5314;
wire x_5315;
wire x_5316;
wire x_5317;
wire x_5318;
wire x_5319;
wire x_5320;
wire x_5321;
wire x_5322;
wire x_5323;
wire x_5324;
wire x_5325;
wire x_5326;
wire x_5327;
wire x_5328;
wire x_5329;
wire x_5330;
wire x_5331;
wire x_5332;
wire x_5333;
wire x_5334;
wire x_5335;
wire x_5336;
wire x_5337;
wire x_5338;
wire x_5339;
wire x_5340;
wire x_5341;
wire x_5342;
wire x_5343;
wire x_5344;
wire x_5345;
wire x_5346;
wire x_5347;
wire x_5348;
wire x_5349;
wire x_5350;
wire x_5351;
wire x_5352;
wire x_5353;
wire x_5354;
wire x_5355;
wire x_5356;
wire x_5357;
wire x_5358;
wire x_5359;
wire x_5360;
wire x_5361;
wire x_5362;
wire x_5363;
wire x_5364;
wire x_5365;
wire x_5366;
wire x_5367;
wire x_5368;
wire x_5369;
wire x_5370;
wire x_5371;
wire x_5372;
wire x_5373;
wire x_5374;
wire x_5375;
wire x_5376;
wire x_5377;
wire x_5378;
wire x_5379;
wire x_5380;
wire x_5381;
wire x_5382;
wire x_5383;
wire x_5384;
wire x_5385;
wire x_5386;
wire x_5387;
wire x_5388;
wire x_5389;
wire x_5390;
wire x_5391;
wire x_5392;
wire x_5393;
wire x_5394;
wire x_5395;
wire x_5396;
wire x_5397;
wire x_5398;
wire x_5399;
wire x_5400;
wire x_5401;
wire x_5402;
wire x_5403;
wire x_5404;
wire x_5405;
wire x_5406;
wire x_5407;
wire x_5408;
wire x_5409;
wire x_5410;
wire x_5411;
wire x_5412;
wire x_5413;
wire x_5414;
wire x_5415;
wire x_5416;
wire x_5417;
wire x_5418;
wire x_5419;
wire x_5420;
wire x_5421;
wire x_5422;
wire x_5423;
wire x_5424;
wire x_5425;
wire x_5426;
wire x_5427;
wire x_5428;
wire x_5429;
wire x_5430;
wire x_5431;
wire x_5432;
wire x_5433;
wire x_5434;
wire x_5435;
wire x_5436;
wire x_5437;
wire x_5438;
wire x_5439;
wire x_5440;
wire x_5441;
wire x_5442;
wire x_5443;
wire x_5444;
wire x_5445;
wire x_5446;
wire x_5447;
wire x_5448;
wire x_5449;
wire x_5450;
wire x_5451;
wire x_5452;
wire x_5453;
wire x_5454;
wire x_5455;
wire x_5456;
wire x_5457;
wire x_5458;
wire x_5459;
wire x_5460;
wire x_5461;
wire x_5462;
wire x_5463;
wire x_5464;
wire x_5465;
wire x_5466;
wire x_5467;
wire x_5468;
wire x_5469;
wire x_5470;
wire x_5471;
wire x_5472;
wire x_5473;
wire x_5474;
wire x_5475;
wire x_5476;
wire x_5477;
wire x_5478;
wire x_5479;
wire x_5480;
wire x_5481;
wire x_5482;
wire x_5483;
wire x_5484;
wire x_5485;
wire x_5486;
wire x_5487;
wire x_5488;
wire x_5489;
wire x_5490;
wire x_5491;
wire x_5492;
wire x_5493;
wire x_5494;
wire x_5495;
wire x_5496;
wire x_5497;
wire x_5498;
wire x_5499;
wire x_5500;
wire x_5501;
wire x_5502;
wire x_5503;
wire x_5504;
wire x_5505;
wire x_5506;
wire x_5507;
wire x_5508;
wire x_5509;
wire x_5510;
wire x_5511;
wire x_5512;
wire x_5513;
wire x_5514;
wire x_5515;
wire x_5516;
wire x_5517;
wire x_5518;
wire x_5519;
wire x_5520;
wire x_5521;
wire x_5522;
wire x_5523;
wire x_5524;
wire x_5525;
wire x_5526;
wire x_5527;
wire x_5528;
wire x_5529;
wire x_5530;
wire x_5531;
wire x_5532;
wire x_5533;
wire x_5534;
wire x_5535;
wire x_5536;
wire x_5537;
wire x_5538;
wire x_5539;
wire x_5540;
wire x_5541;
wire x_5542;
wire x_5543;
wire x_5544;
wire x_5545;
wire x_5546;
wire x_5547;
wire x_5548;
wire x_5549;
wire x_5550;
wire x_5551;
wire x_5552;
wire x_5553;
wire x_5554;
wire x_5555;
wire x_5556;
wire x_5557;
wire x_5558;
wire x_5559;
wire x_5560;
wire x_5561;
wire x_5562;
wire x_5563;
wire x_5564;
wire x_5565;
wire x_5566;
wire x_5567;
wire x_5568;
wire x_5569;
wire x_5570;
wire x_5571;
wire x_5572;
wire x_5573;
wire x_5574;
wire x_5575;
wire x_5576;
wire x_5577;
wire x_5578;
wire x_5579;
wire x_5580;
wire x_5581;
wire x_5582;
wire x_5583;
wire x_5584;
wire x_5585;
wire x_5586;
wire x_5587;
wire x_5588;
wire x_5589;
wire x_5590;
wire x_5591;
wire x_5592;
wire x_5593;
wire x_5594;
wire x_5595;
wire x_5596;
wire x_5597;
wire x_5598;
wire x_5599;
wire x_5600;
wire x_5601;
wire x_5602;
wire x_5603;
wire x_5604;
wire x_5605;
wire x_5606;
wire x_5607;
wire x_5608;
wire x_5609;
wire x_5610;
wire x_5611;
wire x_5612;
wire x_5613;
wire x_5614;
wire x_5615;
wire x_5616;
wire x_5617;
wire x_5618;
wire x_5619;
wire x_5620;
wire x_5621;
wire x_5622;
wire x_5623;
wire x_5624;
wire x_5625;
wire x_5626;
wire x_5627;
wire x_5628;
wire x_5629;
wire x_5630;
wire x_5631;
wire x_5632;
wire x_5633;
wire x_5634;
wire x_5635;
wire x_5636;
wire x_5637;
wire x_5638;
wire x_5639;
wire x_5640;
wire x_5641;
wire x_5642;
wire x_5643;
wire x_5644;
wire x_5645;
wire x_5646;
wire x_5647;
wire x_5648;
wire x_5649;
wire x_5650;
wire x_5651;
wire x_5652;
wire x_5653;
wire x_5654;
wire x_5655;
wire x_5656;
wire x_5657;
wire x_5658;
wire x_5659;
wire x_5660;
wire x_5661;
wire x_5662;
wire x_5663;
wire x_5664;
wire x_5665;
wire x_5666;
wire x_5667;
wire x_5668;
wire x_5669;
wire x_5670;
wire x_5671;
wire x_5672;
wire x_5673;
wire x_5674;
wire x_5675;
wire x_5676;
wire x_5677;
wire x_5678;
wire x_5679;
wire x_5680;
wire x_5681;
wire x_5682;
wire x_5683;
wire x_5684;
wire x_5685;
wire x_5686;
wire x_5687;
wire x_5688;
wire x_5689;
wire x_5690;
wire x_5691;
wire x_5692;
wire x_5693;
wire x_5694;
wire x_5695;
wire x_5696;
wire x_5697;
wire x_5698;
wire x_5699;
wire x_5700;
wire x_5701;
wire x_5702;
wire x_5703;
wire x_5704;
wire x_5705;
wire x_5706;
wire x_5707;
wire x_5708;
wire x_5709;
wire x_5710;
wire x_5711;
wire x_5712;
wire x_5713;
wire x_5714;
wire x_5715;
wire x_5716;
wire x_5717;
wire x_5718;
wire x_5719;
wire x_5720;
wire x_5721;
wire x_5722;
wire x_5723;
wire x_5724;
wire x_5725;
wire x_5726;
wire x_5727;
wire x_5728;
wire x_5729;
wire x_5730;
wire x_5731;
wire x_5732;
wire x_5733;
wire x_5734;
wire x_5735;
wire x_5736;
wire x_5737;
wire x_5738;
wire x_5739;
wire x_5740;
wire x_5741;
wire x_5742;
wire x_5743;
wire x_5744;
wire x_5745;
wire x_5746;
wire x_5747;
wire x_5748;
wire x_5749;
wire x_5750;
wire x_5751;
wire x_5752;
wire x_5753;
wire x_5754;
wire x_5755;
wire x_5756;
wire x_5757;
wire x_5758;
wire x_5759;
wire x_5760;
wire x_5761;
wire x_5762;
wire x_5763;
wire x_5764;
wire x_5765;
wire x_5766;
wire x_5767;
wire x_5768;
wire x_5769;
wire x_5770;
wire x_5771;
wire x_5772;
wire x_5773;
wire x_5774;
wire x_5775;
wire x_5776;
wire x_5777;
wire x_5778;
wire x_5779;
wire x_5780;
wire x_5781;
wire x_5782;
wire x_5783;
wire x_5784;
wire x_5785;
wire x_5786;
wire x_5787;
wire x_5788;
wire x_5789;
wire x_5790;
wire x_5791;
wire x_5792;
wire x_5793;
wire x_5794;
wire x_5795;
wire x_5796;
wire x_5797;
wire x_5798;
wire x_5799;
wire x_5800;
wire x_5801;
wire x_5802;
wire x_5803;
wire x_5804;
wire x_5805;
wire x_5806;
wire x_5807;
wire x_5808;
wire x_5809;
wire x_5810;
wire x_5811;
wire x_5812;
wire x_5813;
wire x_5814;
wire x_5815;
wire x_5816;
wire x_5817;
wire x_5818;
wire x_5819;
wire x_5820;
wire x_5821;
wire x_5822;
wire x_5823;
wire x_5824;
wire x_5825;
wire x_5826;
wire x_5827;
wire x_5828;
wire x_5829;
wire x_5830;
wire x_5831;
wire x_5832;
wire x_5833;
wire x_5834;
wire x_5835;
wire x_5836;
wire x_5837;
wire x_5838;
wire x_5839;
wire x_5840;
wire x_5841;
wire x_5842;
wire x_5843;
wire x_5844;
wire x_5845;
wire x_5846;
wire x_5847;
wire x_5848;
wire x_5849;
wire x_5850;
wire x_5851;
wire x_5852;
wire x_5853;
wire x_5854;
wire x_5855;
wire x_5856;
wire x_5857;
wire x_5858;
wire x_5859;
wire x_5860;
wire x_5861;
wire x_5862;
wire x_5863;
wire x_5864;
wire x_5865;
wire x_5866;
wire x_5867;
wire x_5868;
wire x_5869;
wire x_5870;
wire x_5871;
wire x_5872;
wire x_5873;
wire x_5874;
wire x_5875;
wire x_5876;
wire x_5877;
wire x_5878;
wire x_5879;
wire x_5880;
wire x_5881;
wire x_5882;
wire x_5883;
wire x_5884;
wire x_5885;
wire x_5886;
wire x_5887;
wire x_5888;
wire x_5889;
wire x_5890;
wire x_5891;
wire x_5892;
wire x_5893;
wire x_5894;
wire x_5895;
wire x_5896;
wire x_5897;
wire x_5898;
wire x_5899;
wire x_5900;
wire x_5901;
wire x_5902;
wire x_5903;
wire x_5904;
wire x_5905;
wire x_5906;
wire x_5907;
wire x_5908;
wire x_5909;
wire x_5910;
wire x_5911;
wire x_5912;
wire x_5913;
wire x_5914;
wire x_5915;
wire x_5916;
wire x_5917;
wire x_5918;
wire x_5919;
wire x_5920;
wire x_5921;
wire x_5922;
wire x_5923;
wire x_5924;
wire x_5925;
wire x_5926;
wire x_5927;
wire x_5928;
wire x_5929;
wire x_5930;
wire x_5931;
wire x_5932;
wire x_5933;
wire x_5934;
wire x_5935;
wire x_5936;
wire x_5937;
wire x_5938;
wire x_5939;
wire x_5940;
wire x_5941;
wire x_5942;
wire x_5943;
wire x_5944;
wire x_5945;
wire x_5946;
wire x_5947;
wire x_5948;
wire x_5949;
wire x_5950;
wire x_5951;
wire x_5952;
wire x_5953;
wire x_5954;
wire x_5955;
wire x_5956;
wire x_5957;
wire x_5958;
wire x_5959;
wire x_5960;
wire x_5961;
wire x_5962;
wire x_5963;
wire x_5964;
wire x_5965;
wire x_5966;
wire x_5967;
wire x_5968;
wire x_5969;
wire x_5970;
wire x_5971;
wire x_5972;
wire x_5973;
wire x_5974;
wire x_5975;
wire x_5976;
wire x_5977;
wire x_5978;
wire x_5979;
wire x_5980;
wire x_5981;
wire x_5982;
wire x_5983;
wire x_5984;
wire x_5985;
wire x_5986;
wire x_5987;
wire x_5988;
wire x_5989;
wire x_5990;
wire x_5991;
wire x_5992;
wire x_5993;
wire x_5994;
wire x_5995;
wire x_5996;
wire x_5997;
wire x_5998;
wire x_5999;
wire x_6000;
wire x_6001;
wire x_6002;
wire x_6003;
wire x_6004;
wire x_6005;
wire x_6006;
wire x_6007;
wire x_6008;
wire x_6009;
wire x_6010;
wire x_6011;
wire x_6012;
wire x_6013;
wire x_6014;
wire x_6015;
wire x_6016;
wire x_6017;
wire x_6018;
wire x_6019;
wire x_6020;
wire x_6021;
wire x_6022;
wire x_6023;
wire x_6024;
wire x_6025;
wire x_6026;
wire x_6027;
wire x_6028;
wire x_6029;
wire x_6030;
wire x_6031;
wire x_6032;
wire x_6033;
wire x_6034;
wire x_6035;
wire x_6036;
wire x_6037;
wire x_6038;
wire x_6039;
wire x_6040;
wire x_6041;
wire x_6042;
wire x_6043;
wire x_6044;
wire x_6045;
wire x_6046;
wire x_6047;
wire x_6048;
wire x_6049;
wire x_6050;
wire x_6051;
wire x_6052;
wire x_6053;
wire x_6054;
wire x_6055;
wire x_6056;
wire x_6057;
wire x_6058;
wire x_6059;
wire x_6060;
wire x_6061;
wire x_6062;
wire x_6063;
wire x_6064;
wire x_6065;
wire x_6066;
wire x_6067;
wire x_6068;
wire x_6069;
wire x_6070;
wire x_6071;
wire x_6072;
wire x_6073;
wire x_6074;
wire x_6075;
wire x_6076;
wire x_6077;
wire x_6078;
wire x_6079;
wire x_6080;
wire x_6081;
wire x_6082;
wire x_6083;
wire x_6084;
wire x_6085;
wire x_6086;
wire x_6087;
wire x_6088;
wire x_6089;
wire x_6090;
wire x_6091;
wire x_6092;
wire x_6093;
wire x_6094;
wire x_6095;
wire x_6096;
wire x_6097;
wire x_6098;
wire x_6099;
wire x_6100;
wire x_6101;
wire x_6102;
wire x_6103;
wire x_6104;
wire x_6105;
wire x_6106;
wire x_6107;
wire x_6108;
wire x_6109;
wire x_6110;
wire x_6111;
wire x_6112;
wire x_6113;
wire x_6114;
wire x_6115;
wire x_6116;
wire x_6117;
wire x_6118;
wire x_6119;
wire x_6120;
wire x_6121;
wire x_6122;
wire x_6123;
wire x_6124;
wire x_6125;
wire x_6126;
wire x_6127;
wire x_6128;
wire x_6129;
wire x_6130;
wire x_6131;
wire x_6132;
wire x_6133;
wire x_6134;
wire x_6135;
wire x_6136;
wire x_6137;
wire x_6138;
wire x_6139;
wire x_6140;
wire x_6141;
wire x_6142;
wire x_6143;
wire x_6144;
wire x_6145;
wire x_6146;
wire x_6147;
wire x_6148;
wire x_6149;
wire x_6150;
wire x_6151;
wire x_6152;
wire x_6153;
wire x_6154;
wire x_6155;
wire x_6156;
wire x_6157;
wire x_6158;
wire x_6159;
wire x_6160;
wire x_6161;
wire x_6162;
wire x_6163;
wire x_6164;
wire x_6165;
wire x_6166;
wire x_6167;
wire x_6168;
wire x_6169;
wire x_6170;
wire x_6171;
wire x_6172;
wire x_6173;
wire x_6174;
wire x_6175;
wire x_6176;
wire x_6177;
wire x_6178;
wire x_6179;
wire x_6180;
wire x_6181;
wire x_6182;
wire x_6183;
wire x_6184;
wire x_6185;
wire x_6186;
wire x_6187;
wire x_6188;
wire x_6189;
wire x_6190;
wire x_6191;
wire x_6192;
wire x_6193;
wire x_6194;
wire x_6195;
wire x_6196;
wire x_6197;
wire x_6198;
wire x_6199;
wire x_6200;
wire x_6201;
wire x_6202;
wire x_6203;
wire x_6204;
wire x_6205;
wire x_6206;
wire x_6207;
wire x_6208;
wire x_6209;
wire x_6210;
wire x_6211;
wire x_6212;
wire x_6213;
wire x_6214;
wire x_6215;
wire x_6216;
wire x_6217;
wire x_6218;
wire x_6219;
wire x_6220;
wire x_6221;
wire x_6222;
wire x_6223;
wire x_6224;
wire x_6225;
wire x_6226;
wire x_6227;
wire x_6228;
wire x_6229;
wire x_6230;
wire x_6231;
wire x_6232;
wire x_6233;
wire x_6234;
wire x_6235;
wire x_6236;
wire x_6237;
wire x_6238;
wire x_6239;
wire x_6240;
wire x_6241;
wire x_6242;
wire x_6243;
wire x_6244;
wire x_6245;
wire x_6246;
wire x_6247;
wire x_6248;
wire x_6249;
wire x_6250;
wire x_6251;
wire x_6252;
wire x_6253;
wire x_6254;
wire x_6255;
wire x_6256;
wire x_6257;
wire x_6258;
wire x_6259;
wire x_6260;
wire x_6261;
wire x_6262;
wire x_6263;
wire x_6264;
wire x_6265;
wire x_6266;
wire x_6267;
wire x_6268;
wire x_6269;
wire x_6270;
wire x_6271;
wire x_6272;
wire x_6273;
wire x_6274;
wire x_6275;
wire x_6276;
wire x_6277;
wire x_6278;
wire x_6279;
wire x_6280;
wire x_6281;
wire x_6282;
wire x_6283;
wire x_6284;
wire x_6285;
wire x_6286;
wire x_6287;
wire x_6288;
wire x_6289;
wire x_6290;
wire x_6291;
wire x_6292;
wire x_6293;
wire x_6294;
wire x_6295;
wire x_6296;
wire x_6297;
wire x_6298;
wire x_6299;
wire x_6300;
wire x_6301;
wire x_6302;
wire x_6303;
wire x_6304;
wire x_6305;
wire x_6306;
wire x_6307;
wire x_6308;
wire x_6309;
wire x_6310;
wire x_6311;
wire x_6312;
wire x_6313;
wire x_6314;
wire x_6315;
wire x_6316;
wire x_6317;
wire x_6318;
wire x_6319;
wire x_6320;
wire x_6321;
wire x_6322;
wire x_6323;
wire x_6324;
wire x_6325;
wire x_6326;
wire x_6327;
wire x_6328;
wire x_6329;
wire x_6330;
wire x_6331;
wire x_6332;
wire x_6333;
wire x_6334;
wire x_6335;
wire x_6336;
wire x_6337;
wire x_6338;
wire x_6339;
wire x_6340;
wire x_6341;
wire x_6342;
wire x_6343;
wire x_6344;
wire x_6345;
wire x_6346;
wire x_6347;
wire x_6348;
wire x_6349;
wire x_6350;
wire x_6351;
wire x_6352;
wire x_6353;
wire x_6354;
wire x_6355;
wire x_6356;
wire x_6357;
wire x_6358;
wire x_6359;
wire x_6360;
wire x_6361;
wire x_6362;
wire x_6363;
wire x_6364;
wire x_6365;
wire x_6366;
wire x_6367;
wire x_6368;
wire x_6369;
wire x_6370;
wire x_6371;
wire x_6372;
wire x_6373;
wire x_6374;
wire x_6375;
wire x_6376;
wire x_6377;
wire x_6378;
wire x_6379;
wire x_6380;
wire x_6381;
wire x_6382;
wire x_6383;
wire x_6384;
wire x_6385;
wire x_6386;
wire x_6387;
wire x_6388;
wire x_6389;
wire x_6390;
wire x_6391;
wire x_6392;
wire x_6393;
wire x_6394;
wire x_6395;
wire x_6396;
wire x_6397;
wire x_6398;
wire x_6399;
wire x_6400;
wire x_6401;
wire x_6402;
wire x_6403;
wire x_6404;
wire x_6405;
wire x_6406;
wire x_6407;
wire x_6408;
wire x_6409;
wire x_6410;
wire x_6411;
wire x_6412;
wire x_6413;
wire x_6414;
wire x_6415;
wire x_6416;
wire x_6417;
wire x_6418;
wire x_6419;
wire x_6420;
wire x_6421;
wire x_6422;
wire x_6423;
wire x_6424;
wire x_6425;
wire x_6426;
wire x_6427;
wire x_6428;
wire x_6429;
wire x_6430;
wire x_6431;
wire x_6432;
wire x_6433;
wire x_6434;
wire x_6435;
wire x_6436;
wire x_6437;
wire x_6438;
wire x_6439;
wire x_6440;
wire x_6441;
wire x_6442;
wire x_6443;
wire x_6444;
wire x_6445;
wire x_6446;
wire x_6447;
wire x_6448;
wire x_6449;
wire x_6450;
wire x_6451;
wire x_6452;
wire x_6453;
wire x_6454;
wire x_6455;
wire x_6456;
wire x_6457;
wire x_6458;
wire x_6459;
wire x_6460;
wire x_6461;
wire x_6462;
wire x_6463;
wire x_6464;
wire x_6465;
wire x_6466;
wire x_6467;
wire x_6468;
wire x_6469;
wire x_6470;
wire x_6471;
wire x_6472;
wire x_6473;
wire x_6474;
wire x_6475;
wire x_6476;
wire x_6477;
wire x_6478;
wire x_6479;
wire x_6480;
wire x_6481;
wire x_6482;
wire x_6483;
wire x_6484;
wire x_6485;
wire x_6486;
wire x_6487;
wire x_6488;
wire x_6489;
wire x_6490;
wire x_6491;
wire x_6492;
wire x_6493;
wire x_6494;
wire x_6495;
wire x_6496;
wire x_6497;
wire x_6498;
wire x_6499;
wire x_6500;
wire x_6501;
wire x_6502;
wire x_6503;
wire x_6504;
wire x_6505;
wire x_6506;
wire x_6507;
wire x_6508;
wire x_6509;
wire x_6510;
wire x_6511;
wire x_6512;
wire x_6513;
wire x_6514;
wire x_6515;
wire x_6516;
wire x_6517;
wire x_6518;
wire x_6519;
wire x_6520;
wire x_6521;
wire x_6522;
wire x_6523;
wire x_6524;
wire x_6525;
wire x_6526;
wire x_6527;
wire x_6528;
wire x_6529;
wire x_6530;
wire x_6531;
wire x_6532;
wire x_6533;
wire x_6534;
wire x_6535;
wire x_6536;
wire x_6537;
wire x_6538;
wire x_6539;
wire x_6540;
wire x_6541;
wire x_6542;
wire x_6543;
wire x_6544;
wire x_6545;
wire x_6546;
wire x_6547;
wire x_6548;
wire x_6549;
wire x_6550;
wire x_6551;
wire x_6552;
wire x_6553;
wire x_6554;
wire x_6555;
wire x_6556;
wire x_6557;
wire x_6558;
wire x_6559;
wire x_6560;
wire x_6561;
wire x_6562;
wire x_6563;
wire x_6564;
wire x_6565;
wire x_6566;
wire x_6567;
wire x_6568;
wire x_6569;
wire x_6570;
wire x_6571;
wire x_6572;
wire x_6573;
wire x_6574;
wire x_6575;
wire x_6576;
wire x_6577;
wire x_6578;
wire x_6579;
wire x_6580;
wire x_6581;
wire x_6582;
wire x_6583;
wire x_6584;
wire x_6585;
wire x_6586;
wire x_6587;
wire x_6588;
wire x_6589;
wire x_6590;
wire x_6591;
wire x_6592;
wire x_6593;
wire x_6594;
wire x_6595;
wire x_6596;
wire x_6597;
wire x_6598;
wire x_6599;
wire x_6600;
wire x_6601;
wire x_6602;
wire x_6603;
wire x_6604;
wire x_6605;
wire x_6606;
wire x_6607;
wire x_6608;
wire x_6609;
wire x_6610;
wire x_6611;
wire x_6612;
wire x_6613;
wire x_6614;
wire x_6615;
wire x_6616;
wire x_6617;
wire x_6618;
wire x_6619;
wire x_6620;
wire x_6621;
wire x_6622;
wire x_6623;
wire x_6624;
wire x_6625;
wire x_6626;
wire x_6627;
wire x_6628;
wire x_6629;
wire x_6630;
wire x_6631;
wire x_6632;
wire x_6633;
wire x_6634;
wire x_6635;
wire x_6636;
wire x_6637;
wire x_6638;
wire x_6639;
wire x_6640;
wire x_6641;
wire x_6642;
wire x_6643;
wire x_6644;
wire x_6645;
wire x_6646;
wire x_6647;
wire x_6648;
wire x_6649;
wire x_6650;
wire x_6651;
wire x_6652;
wire x_6653;
wire x_6654;
wire x_6655;
wire x_6656;
wire x_6657;
wire x_6658;
wire x_6659;
wire x_6660;
wire x_6661;
wire x_6662;
wire x_6663;
wire x_6664;
wire x_6665;
wire x_6666;
wire x_6667;
wire x_6668;
wire x_6669;
wire x_6670;
wire x_6671;
wire x_6672;
wire x_6673;
wire x_6674;
wire x_6675;
wire x_6676;
wire x_6677;
wire x_6678;
wire x_6679;
wire x_6680;
wire x_6681;
wire x_6682;
wire x_6683;
wire x_6684;
wire x_6685;
wire x_6686;
wire x_6687;
wire x_6688;
wire x_6689;
wire x_6690;
wire x_6691;
wire x_6692;
wire x_6693;
wire x_6694;
wire x_6695;
wire x_6696;
wire x_6697;
wire x_6698;
wire x_6699;
wire x_6700;
wire x_6701;
wire x_6702;
wire x_6703;
wire x_6704;
wire x_6705;
wire x_6706;
wire x_6707;
wire x_6708;
wire x_6709;
wire x_6710;
wire x_6711;
wire x_6712;
wire x_6713;
wire x_6714;
wire x_6715;
wire x_6716;
wire x_6717;
wire x_6718;
wire x_6719;
wire x_6720;
wire x_6721;
wire x_6722;
wire x_6723;
wire x_6724;
wire x_6725;
wire x_6726;
wire x_6727;
wire x_6728;
wire x_6729;
wire x_6730;
wire x_6731;
wire x_6732;
wire x_6733;
wire x_6734;
wire x_6735;
wire x_6736;
wire x_6737;
wire x_6738;
wire x_6739;
wire x_6740;
wire x_6741;
wire x_6742;
wire x_6743;
wire x_6744;
wire x_6745;
wire x_6746;
wire x_6747;
wire x_6748;
wire x_6749;
wire x_6750;
wire x_6751;
wire x_6752;
wire x_6753;
wire x_6754;
wire x_6755;
wire x_6756;
wire x_6757;
wire x_6758;
wire x_6759;
wire x_6760;
wire x_6761;
wire x_6762;
wire x_6763;
wire x_6764;
wire x_6765;
wire x_6766;
wire x_6767;
wire x_6768;
wire x_6769;
wire x_6770;
wire x_6771;
wire x_6772;
wire x_6773;
wire x_6774;
wire x_6775;
wire x_6776;
wire x_6777;
wire x_6778;
wire x_6779;
wire x_6780;
wire x_6781;
wire x_6782;
wire x_6783;
wire x_6784;
wire x_6785;
wire x_6786;
wire x_6787;
wire x_6788;
wire x_6789;
wire x_6790;
wire x_6791;
wire x_6792;
wire x_6793;
wire x_6794;
wire x_6795;
wire x_6796;
wire x_6797;
wire x_6798;
wire x_6799;
wire x_6800;
wire x_6801;
wire x_6802;
wire x_6803;
wire x_6804;
wire x_6805;
wire x_6806;
wire x_6807;
wire x_6808;
wire x_6809;
wire x_6810;
wire x_6811;
wire x_6812;
wire x_6813;
wire x_6814;
wire x_6815;
wire x_6816;
wire x_6817;
wire x_6818;
wire x_6819;
wire x_6820;
wire x_6821;
wire x_6822;
wire x_6823;
wire x_6824;
wire x_6825;
wire x_6826;
wire x_6827;
wire x_6828;
wire x_6829;
wire x_6830;
wire x_6831;
wire x_6832;
wire x_6833;
wire x_6834;
wire x_6835;
wire x_6836;
wire x_6837;
wire x_6838;
wire x_6839;
wire x_6840;
wire x_6841;
wire x_6842;
wire x_6843;
wire x_6844;
wire x_6845;
wire x_6846;
wire x_6847;
wire x_6848;
wire x_6849;
wire x_6850;
wire x_6851;
wire x_6852;
wire x_6853;
wire x_6854;
wire x_6855;
wire x_6856;
wire x_6857;
wire x_6858;
wire x_6859;
wire x_6860;
wire x_6861;
wire x_6862;
wire x_6863;
wire x_6864;
wire x_6865;
wire x_6866;
wire x_6867;
wire x_6868;
wire x_6869;
wire x_6870;
wire x_6871;
wire x_6872;
wire x_6873;
wire x_6874;
wire x_6875;
wire x_6876;
wire x_6877;
wire x_6878;
wire x_6879;
wire x_6880;
wire x_6881;
wire x_6882;
wire x_6883;
wire x_6884;
wire x_6885;
wire x_6886;
wire x_6887;
wire x_6888;
wire x_6889;
wire x_6890;
wire x_6891;
wire x_6892;
wire x_6893;
wire x_6894;
wire x_6895;
wire x_6896;
wire x_6897;
wire x_6898;
wire x_6899;
wire x_6900;
wire x_6901;
wire x_6902;
wire x_6903;
wire x_6904;
wire x_6905;
wire x_6906;
wire x_6907;
wire x_6908;
wire x_6909;
wire x_6910;
wire x_6911;
wire x_6912;
wire x_6913;
wire x_6914;
wire x_6915;
wire x_6916;
wire x_6917;
wire x_6918;
wire x_6919;
wire x_6920;
wire x_6921;
wire x_6922;
wire x_6923;
wire x_6924;
wire x_6925;
wire x_6926;
wire x_6927;
wire x_6928;
wire x_6929;
wire x_6930;
wire x_6931;
wire x_6932;
wire x_6933;
wire x_6934;
wire x_6935;
wire x_6936;
wire x_6937;
wire x_6938;
wire x_6939;
wire x_6940;
wire x_6941;
wire x_6942;
wire x_6943;
wire x_6944;
wire x_6945;
wire x_6946;
wire x_6947;
wire x_6948;
wire x_6949;
wire x_6950;
wire x_6951;
wire x_6952;
wire x_6953;
wire x_6954;
wire x_6955;
wire x_6956;
wire x_6957;
wire x_6958;
wire x_6959;
wire x_6960;
wire x_6961;
wire x_6962;
wire x_6963;
wire x_6964;
wire x_6965;
wire x_6966;
wire x_6967;
wire x_6968;
wire x_6969;
wire x_6970;
wire x_6971;
wire x_6972;
wire x_6973;
wire x_6974;
wire x_6975;
wire x_6976;
wire x_6977;
wire x_6978;
wire x_6979;
wire x_6980;
wire x_6981;
wire x_6982;
wire x_6983;
wire x_6984;
wire x_6985;
wire x_6986;
wire x_6987;
wire x_6988;
wire x_6989;
wire x_6990;
wire x_6991;
wire x_6992;
wire x_6993;
wire x_6994;
wire x_6995;
wire x_6996;
wire x_6997;
wire x_6998;
wire x_6999;
wire x_7000;
wire x_7001;
wire x_7002;
wire x_7003;
wire x_7004;
wire x_7005;
wire x_7006;
wire x_7007;
wire x_7008;
wire x_7009;
wire x_7010;
wire x_7011;
wire x_7012;
wire x_7013;
wire x_7014;
wire x_7015;
wire x_7016;
wire x_7017;
wire x_7018;
wire x_7019;
wire x_7020;
wire x_7021;
wire x_7022;
wire x_7023;
wire x_7024;
wire x_7025;
wire x_7026;
wire x_7027;
wire x_7028;
wire x_7029;
wire x_7030;
wire x_7031;
wire x_7032;
wire x_7033;
wire x_7034;
wire x_7035;
wire x_7036;
wire x_7037;
wire x_7038;
wire x_7039;
wire x_7040;
wire x_7041;
wire x_7042;
wire x_7043;
wire x_7044;
wire x_7045;
wire x_7046;
wire x_7047;
wire x_7048;
wire x_7049;
wire x_7050;
wire x_7051;
wire x_7052;
wire x_7053;
wire x_7054;
wire x_7055;
wire x_7056;
wire x_7057;
wire x_7058;
wire x_7059;
wire x_7060;
wire x_7061;
wire x_7062;
wire x_7063;
wire x_7064;
wire x_7065;
wire x_7066;
wire x_7067;
wire x_7068;
wire x_7069;
wire x_7070;
wire x_7071;
wire x_7072;
wire x_7073;
wire x_7074;
wire x_7075;
wire x_7076;
wire x_7077;
wire x_7078;
wire x_7079;
wire x_7080;
wire x_7081;
wire x_7082;
wire x_7083;
wire x_7084;
wire x_7085;
wire x_7086;
wire x_7087;
wire x_7088;
wire x_7089;
wire x_7090;
wire x_7091;
wire x_7092;
wire x_7093;
wire x_7094;
wire x_7095;
wire x_7096;
wire x_7097;
wire x_7098;
wire x_7099;
wire x_7100;
wire x_7101;
wire x_7102;
wire x_7103;
wire x_7104;
wire x_7105;
wire x_7106;
wire x_7107;
wire x_7108;
wire x_7109;
wire x_7110;
wire x_7111;
wire x_7112;
wire x_7113;
wire x_7114;
wire x_7115;
wire x_7116;
wire x_7117;
wire x_7118;
wire x_7119;
wire x_7120;
wire x_7121;
wire x_7122;
wire x_7123;
wire x_7124;
wire x_7125;
wire x_7126;
wire x_7127;
wire x_7128;
wire x_7129;
wire x_7130;
wire x_7131;
wire x_7132;
wire x_7133;
wire x_7134;
wire x_7135;
wire x_7136;
wire x_7137;
wire x_7138;
wire x_7139;
wire x_7140;
wire x_7141;
wire x_7142;
wire x_7143;
wire x_7144;
wire x_7145;
wire x_7146;
wire x_7147;
wire x_7148;
wire x_7149;
wire x_7150;
wire x_7151;
wire x_7152;
wire x_7153;
wire x_7154;
wire x_7155;
wire x_7156;
wire x_7157;
wire x_7158;
wire x_7159;
wire x_7160;
wire x_7161;
wire x_7162;
wire x_7163;
wire x_7164;
wire x_7165;
wire x_7166;
wire x_7167;
wire x_7168;
wire x_7169;
wire x_7170;
wire x_7171;
wire x_7172;
wire x_7173;
wire x_7174;
wire x_7175;
wire x_7176;
wire x_7177;
wire x_7178;
wire x_7179;
wire x_7180;
wire x_7181;
wire x_7182;
wire x_7183;
wire x_7184;
wire x_7185;
wire x_7186;
wire x_7187;
wire x_7188;
wire x_7189;
wire x_7190;
wire x_7191;
wire x_7192;
wire x_7193;
wire x_7194;
wire x_7195;
wire x_7196;
wire x_7197;
wire x_7198;
wire x_7199;
wire x_7200;
wire x_7201;
wire x_7202;
wire x_7203;
wire x_7204;
wire x_7205;
wire x_7206;
wire x_7207;
wire x_7208;
wire x_7209;
wire x_7210;
wire x_7211;
wire x_7212;
wire x_7213;
wire x_7214;
wire x_7215;
wire x_7216;
wire x_7217;
wire x_7218;
wire x_7219;
wire x_7220;
wire x_7221;
wire x_7222;
wire x_7223;
wire x_7224;
wire x_7225;
wire x_7226;
wire x_7227;
wire x_7228;
wire x_7229;
wire x_7230;
wire x_7231;
wire x_7232;
wire x_7233;
wire x_7234;
wire x_7235;
wire x_7236;
wire x_7237;
wire x_7238;
wire x_7239;
wire x_7240;
wire x_7241;
wire x_7242;
wire x_7243;
wire x_7244;
wire x_7245;
wire x_7246;
wire x_7247;
wire x_7248;
wire x_7249;
wire x_7250;
wire x_7251;
wire x_7252;
wire x_7253;
wire x_7254;
wire x_7255;
wire x_7256;
wire x_7257;
wire x_7258;
wire x_7259;
wire x_7260;
wire x_7261;
wire x_7262;
wire x_7263;
wire x_7264;
wire x_7265;
wire x_7266;
wire x_7267;
wire x_7268;
wire x_7269;
wire x_7270;
wire x_7271;
wire x_7272;
wire x_7273;
wire x_7274;
wire x_7275;
wire x_7276;
wire x_7277;
wire x_7278;
wire x_7279;
wire x_7280;
wire x_7281;
wire x_7282;
wire x_7283;
wire x_7284;
wire x_7285;
wire x_7286;
wire x_7287;
wire x_7288;
wire x_7289;
wire x_7290;
wire x_7291;
wire x_7292;
wire x_7293;
wire x_7294;
wire x_7295;
wire x_7296;
wire x_7297;
wire x_7298;
wire x_7299;
wire x_7300;
wire x_7301;
wire x_7302;
wire x_7303;
wire x_7304;
wire x_7305;
wire x_7306;
wire x_7307;
wire x_7308;
wire x_7309;
wire x_7310;
wire x_7311;
wire x_7312;
wire x_7313;
wire x_7314;
wire x_7315;
wire x_7316;
wire x_7317;
wire x_7318;
wire x_7319;
wire x_7320;
wire x_7321;
wire x_7322;
wire x_7323;
wire x_7324;
wire x_7325;
wire x_7326;
wire x_7327;
wire x_7328;
wire x_7329;
wire x_7330;
wire x_7331;
wire x_7332;
wire x_7333;
wire x_7334;
wire x_7335;
wire x_7336;
wire x_7337;
wire x_7338;
wire x_7339;
wire x_7340;
wire x_7341;
wire x_7342;
wire x_7343;
wire x_7344;
wire x_7345;
wire x_7346;
wire x_7347;
wire x_7348;
wire x_7349;
wire x_7350;
wire x_7351;
wire x_7352;
wire x_7353;
wire x_7354;
wire x_7355;
wire x_7356;
wire x_7357;
wire x_7358;
wire x_7359;
wire x_7360;
wire x_7361;
wire x_7362;
wire x_7363;
wire x_7364;
wire x_7365;
wire x_7366;
wire x_7367;
wire x_7368;
wire x_7369;
wire x_7370;
wire x_7371;
wire x_7372;
wire x_7373;
wire x_7374;
wire x_7375;
wire x_7376;
wire x_7377;
wire x_7378;
wire x_7379;
wire x_7380;
wire x_7381;
wire x_7382;
wire x_7383;
wire x_7384;
wire x_7385;
wire x_7386;
wire x_7387;
wire x_7388;
wire x_7389;
wire x_7390;
wire x_7391;
wire x_7392;
wire x_7393;
wire x_7394;
wire x_7395;
wire x_7396;
wire x_7397;
wire x_7398;
wire x_7399;
wire x_7400;
wire x_7401;
wire x_7402;
wire x_7403;
wire x_7404;
wire x_7405;
wire x_7406;
wire x_7407;
wire x_7408;
wire x_7409;
wire x_7410;
wire x_7411;
wire x_7412;
wire x_7413;
wire x_7414;
wire x_7415;
wire x_7416;
wire x_7417;
wire x_7418;
wire x_7419;
wire x_7420;
wire x_7421;
wire x_7422;
wire x_7423;
wire x_7424;
wire x_7425;
wire x_7426;
wire x_7427;
wire x_7428;
wire x_7429;
wire x_7430;
wire x_7431;
wire x_7432;
wire x_7433;
wire x_7434;
wire x_7435;
wire x_7436;
wire x_7437;
wire x_7438;
wire x_7439;
wire x_7440;
wire x_7441;
wire x_7442;
wire x_7443;
wire x_7444;
wire x_7445;
wire x_7446;
wire x_7447;
wire x_7448;
wire x_7449;
wire x_7450;
wire x_7451;
wire x_7452;
wire x_7453;
wire x_7454;
wire x_7455;
wire x_7456;
wire x_7457;
wire x_7458;
wire x_7459;
wire x_7460;
wire x_7461;
wire x_7462;
wire x_7463;
wire x_7464;
wire x_7465;
wire x_7466;
wire x_7467;
wire x_7468;
wire x_7469;
wire x_7470;
wire x_7471;
wire x_7472;
wire x_7473;
wire x_7474;
wire x_7475;
wire x_7476;
wire x_7477;
wire x_7478;
wire x_7479;
wire x_7480;
wire x_7481;
wire x_7482;
wire x_7483;
wire x_7484;
wire x_7485;
wire x_7486;
wire x_7487;
wire x_7488;
wire x_7489;
wire x_7490;
wire x_7491;
wire x_7492;
wire x_7493;
wire x_7494;
wire x_7495;
wire x_7496;
wire x_7497;
wire x_7498;
wire x_7499;
wire x_7500;
wire x_7501;
wire x_7502;
wire x_7503;
wire x_7504;
wire x_7505;
wire x_7506;
wire x_7507;
wire x_7508;
wire x_7509;
wire x_7510;
wire x_7511;
wire x_7512;
wire x_7513;
wire x_7514;
wire x_7515;
wire x_7516;
wire x_7517;
wire x_7518;
wire x_7519;
wire x_7520;
wire x_7521;
wire x_7522;
wire x_7523;
wire x_7524;
wire x_7525;
wire x_7526;
wire x_7527;
wire x_7528;
wire x_7529;
wire x_7530;
wire x_7531;
wire x_7532;
wire x_7533;
wire x_7534;
wire x_7535;
wire x_7536;
wire x_7537;
wire x_7538;
wire x_7539;
wire x_7540;
wire x_7541;
wire x_7542;
wire x_7543;
wire x_7544;
wire x_7545;
wire x_7546;
wire x_7547;
wire x_7548;
wire x_7549;
wire x_7550;
wire x_7551;
wire x_7552;
wire x_7553;
wire x_7554;
wire x_7555;
wire x_7556;
wire x_7557;
wire x_7558;
wire x_7559;
wire x_7560;
wire x_7561;
wire x_7562;
wire x_7563;
wire x_7564;
wire x_7565;
wire x_7566;
wire x_7567;
wire x_7568;
wire x_7569;
wire x_7570;
wire x_7571;
wire x_7572;
wire x_7573;
wire x_7574;
wire x_7575;
wire x_7576;
wire x_7577;
wire x_7578;
wire x_7579;
wire x_7580;
wire x_7581;
wire x_7582;
wire x_7583;
wire x_7584;
wire x_7585;
wire x_7586;
wire x_7587;
wire x_7588;
wire x_7589;
wire x_7590;
wire x_7591;
wire x_7592;
wire x_7593;
wire x_7594;
wire x_7595;
wire x_7596;
wire x_7597;
wire x_7598;
wire x_7599;
wire x_7600;
wire x_7601;
wire x_7602;
wire x_7603;
wire x_7604;
wire x_7605;
wire x_7606;
wire x_7607;
wire x_7608;
wire x_7609;
wire x_7610;
wire x_7611;
wire x_7612;
wire x_7613;
wire x_7614;
wire x_7615;
wire x_7616;
wire x_7617;
wire x_7618;
wire x_7619;
wire x_7620;
wire x_7621;
wire x_7622;
wire x_7623;
wire x_7624;
wire x_7625;
wire x_7626;
wire x_7627;
wire x_7628;
wire x_7629;
wire x_7630;
wire x_7631;
wire x_7632;
wire x_7633;
wire x_7634;
wire x_7635;
wire x_7636;
wire x_7637;
wire x_7638;
wire x_7639;
wire x_7640;
wire x_7641;
wire x_7642;
wire x_7643;
wire x_7644;
wire x_7645;
wire x_7646;
wire x_7647;
wire x_7648;
wire x_7649;
wire x_7650;
wire x_7651;
wire x_7652;
wire x_7653;
wire x_7654;
wire x_7655;
wire x_7656;
wire x_7657;
wire x_7658;
wire x_7659;
wire x_7660;
wire x_7661;
wire x_7662;
wire x_7663;
wire x_7664;
wire x_7665;
wire x_7666;
wire x_7667;
wire x_7668;
wire x_7669;
wire x_7670;
wire x_7671;
wire x_7672;
wire x_7673;
wire x_7674;
wire x_7675;
wire x_7676;
wire x_7677;
wire x_7678;
wire x_7679;
wire x_7680;
wire x_7681;
wire x_7682;
wire x_7683;
wire x_7684;
wire x_7685;
wire x_7686;
wire x_7687;
wire x_7688;
wire x_7689;
wire x_7690;
wire x_7691;
wire x_7692;
wire x_7693;
wire x_7694;
wire x_7695;
wire x_7696;
wire x_7697;
wire x_7698;
wire x_7699;
wire x_7700;
wire x_7701;
wire x_7702;
wire x_7703;
wire x_7704;
wire x_7705;
wire x_7706;
wire x_7707;
wire x_7708;
wire x_7709;
wire x_7710;
wire x_7711;
wire x_7712;
wire x_7713;
wire x_7714;
wire x_7715;
wire x_7716;
wire x_7717;
wire x_7718;
wire x_7719;
wire x_7720;
wire x_7721;
wire x_7722;
wire x_7723;
wire x_7724;
wire x_7725;
wire x_7726;
wire x_7727;
wire x_7728;
wire x_7729;
wire x_7730;
wire x_7731;
wire x_7732;
wire x_7733;
wire x_7734;
wire x_7735;
wire x_7736;
wire x_7737;
wire x_7738;
wire x_7739;
wire x_7740;
wire x_7741;
wire x_7742;
wire x_7743;
wire x_7744;
wire x_7745;
wire x_7746;
wire x_7747;
wire x_7748;
wire x_7749;
wire x_7750;
wire x_7751;
wire x_7752;
wire x_7753;
wire x_7754;
wire x_7755;
wire x_7756;
wire x_7757;
wire x_7758;
wire x_7759;
wire x_7760;
wire x_7761;
wire x_7762;
wire x_7763;
wire x_7764;
wire x_7765;
wire x_7766;
wire x_7767;
wire x_7768;
wire x_7769;
wire x_7770;
wire x_7771;
wire x_7772;
wire x_7773;
wire x_7774;
wire x_7775;
wire x_7776;
wire x_7777;
wire x_7778;
wire x_7779;
wire x_7780;
wire x_7781;
wire x_7782;
wire x_7783;
wire x_7784;
wire x_7785;
wire x_7786;
wire x_7787;
wire x_7788;
wire x_7789;
wire x_7790;
wire x_7791;
wire x_7792;
wire x_7793;
wire x_7794;
wire x_7795;
wire x_7796;
wire x_7797;
wire x_7798;
wire x_7799;
wire x_7800;
wire x_7801;
wire x_7802;
wire x_7803;
wire x_7804;
wire x_7805;
wire x_7806;
wire x_7807;
wire x_7808;
wire x_7809;
wire x_7810;
wire x_7811;
wire x_7812;
wire x_7813;
wire x_7814;
wire x_7815;
wire x_7816;
wire x_7817;
wire x_7818;
wire x_7819;
wire x_7820;
wire x_7821;
wire x_7822;
wire x_7823;
wire x_7824;
wire x_7825;
wire x_7826;
wire x_7827;
wire x_7828;
wire x_7829;
wire x_7830;
wire x_7831;
wire x_7832;
wire x_7833;
wire x_7834;
wire x_7835;
wire x_7836;
wire x_7837;
wire x_7838;
wire x_7839;
wire x_7840;
wire x_7841;
wire x_7842;
wire x_7843;
wire x_7844;
wire x_7845;
wire x_7846;
wire x_7847;
wire x_7848;
wire x_7849;
wire x_7850;
wire x_7851;
wire x_7852;
wire x_7853;
wire x_7854;
wire x_7855;
wire x_7856;
wire x_7857;
wire x_7858;
wire x_7859;
wire x_7860;
wire x_7861;
wire x_7862;
wire x_7863;
wire x_7864;
wire x_7865;
wire x_7866;
wire x_7867;
wire x_7868;
wire x_7869;
wire x_7870;
wire x_7871;
wire x_7872;
wire x_7873;
wire x_7874;
wire x_7875;
wire x_7876;
wire x_7877;
wire x_7878;
wire x_7879;
wire x_7880;
wire x_7881;
wire x_7882;
wire x_7883;
wire x_7884;
wire x_7885;
wire x_7886;
wire x_7887;
wire x_7888;
wire x_7889;
wire x_7890;
wire x_7891;
wire x_7892;
wire x_7893;
wire x_7894;
wire x_7895;
wire x_7896;
wire x_7897;
wire x_7898;
wire x_7899;
wire x_7900;
wire x_7901;
wire x_7902;
wire x_7903;
wire x_7904;
wire x_7905;
wire x_7906;
wire x_7907;
wire x_7908;
wire x_7909;
wire x_7910;
wire x_7911;
wire x_7912;
wire x_7913;
wire x_7914;
wire x_7915;
wire x_7916;
wire x_7917;
wire x_7918;
wire x_7919;
wire x_7920;
wire x_7921;
wire x_7922;
wire x_7923;
wire x_7924;
wire x_7925;
wire x_7926;
wire x_7927;
wire x_7928;
wire x_7929;
wire x_7930;
wire x_7931;
wire x_7932;
wire x_7933;
wire x_7934;
wire x_7935;
wire x_7936;
wire x_7937;
wire x_7938;
wire x_7939;
wire x_7940;
wire x_7941;
wire x_7942;
wire x_7943;
wire x_7944;
wire x_7945;
wire x_7946;
wire x_7947;
wire x_7948;
wire x_7949;
wire x_7950;
wire x_7951;
wire x_7952;
wire x_7953;
wire x_7954;
wire x_7955;
wire x_7956;
wire x_7957;
wire x_7958;
wire x_7959;
wire x_7960;
wire x_7961;
wire x_7962;
wire x_7963;
wire x_7964;
wire x_7965;
wire x_7966;
wire x_7967;
wire x_7968;
wire x_7969;
wire x_7970;
wire x_7971;
wire x_7972;
wire x_7973;
wire x_7974;
wire x_7975;
wire x_7976;
wire x_7977;
wire x_7978;
wire x_7979;
wire x_7980;
wire x_7981;
wire x_7982;
wire x_7983;
wire x_7984;
wire x_7985;
wire x_7986;
wire x_7987;
wire x_7988;
wire x_7989;
wire x_7990;
wire x_7991;
wire x_7992;
wire x_7993;
wire x_7994;
wire x_7995;
wire x_7996;
wire x_7997;
wire x_7998;
wire x_7999;
wire x_8000;
wire x_8001;
wire x_8002;
wire x_8003;
wire x_8004;
wire x_8005;
wire x_8006;
wire x_8007;
wire x_8008;
wire x_8009;
wire x_8010;
wire x_8011;
wire x_8012;
wire x_8013;
wire x_8014;
wire x_8015;
wire x_8016;
wire x_8017;
wire x_8018;
wire x_8019;
wire x_8020;
wire x_8021;
wire x_8022;
wire x_8023;
wire x_8024;
wire x_8025;
wire x_8026;
wire x_8027;
wire x_8028;
wire x_8029;
wire x_8030;
wire x_8031;
wire x_8032;
wire x_8033;
wire x_8034;
wire x_8035;
wire x_8036;
wire x_8037;
wire x_8038;
wire x_8039;
wire x_8040;
wire x_8041;
wire x_8042;
wire x_8043;
wire x_8044;
wire x_8045;
wire x_8046;
wire x_8047;
wire x_8048;
wire x_8049;
wire x_8050;
wire x_8051;
wire x_8052;
wire x_8053;
wire x_8054;
wire x_8055;
wire x_8056;
wire x_8057;
wire x_8058;
wire x_8059;
wire x_8060;
wire x_8061;
wire x_8062;
wire x_8063;
wire x_8064;
wire x_8065;
wire x_8066;
wire x_8067;
wire x_8068;
wire x_8069;
wire x_8070;
wire x_8071;
wire x_8072;
wire x_8073;
wire x_8074;
wire x_8075;
wire x_8076;
wire x_8077;
wire x_8078;
wire x_8079;
wire x_8080;
wire x_8081;
wire x_8082;
wire x_8083;
wire x_8084;
wire x_8085;
wire x_8086;
wire x_8087;
wire x_8088;
wire x_8089;
wire x_8090;
wire x_8091;
wire x_8092;
wire x_8093;
wire x_8094;
wire x_8095;
wire x_8096;
wire x_8097;
wire x_8098;
wire x_8099;
wire x_8100;
wire x_8101;
wire x_8102;
wire x_8103;
wire x_8104;
wire x_8105;
wire x_8106;
wire x_8107;
wire x_8108;
wire x_8109;
wire x_8110;
wire x_8111;
wire x_8112;
wire x_8113;
wire x_8114;
wire x_8115;
wire x_8116;
wire x_8117;
wire x_8118;
wire x_8119;
wire x_8120;
wire x_8121;
wire x_8122;
wire x_8123;
wire x_8124;
wire x_8125;
wire x_8126;
wire x_8127;
wire x_8128;
wire x_8129;
wire x_8130;
wire x_8131;
wire x_8132;
wire x_8133;
wire x_8134;
wire x_8135;
wire x_8136;
wire x_8137;
wire x_8138;
wire x_8139;
wire x_8140;
wire x_8141;
wire x_8142;
wire x_8143;
wire x_8144;
wire x_8145;
wire x_8146;
wire x_8147;
wire x_8148;
wire x_8149;
wire x_8150;
wire x_8151;
wire x_8152;
wire x_8153;
wire x_8154;
wire x_8155;
wire x_8156;
wire x_8157;
wire x_8158;
wire x_8159;
wire x_8160;
wire x_8161;
wire x_8162;
wire x_8163;
wire x_8164;
wire x_8165;
wire x_8166;
wire x_8167;
wire x_8168;
wire x_8169;
wire x_8170;
wire x_8171;
wire x_8172;
wire x_8173;
wire x_8174;
wire x_8175;
wire x_8176;
wire x_8177;
wire x_8178;
wire x_8179;
wire x_8180;
wire x_8181;
wire x_8182;
wire x_8183;
wire x_8184;
wire x_8185;
wire x_8186;
wire x_8187;
wire x_8188;
wire x_8189;
wire x_8190;
wire x_8191;
wire x_8192;
wire x_8193;
wire x_8194;
wire x_8195;
wire x_8196;
wire x_8197;
wire x_8198;
wire x_8199;
wire x_8200;
wire x_8201;
wire x_8202;
wire x_8203;
wire x_8204;
wire x_8205;
wire x_8206;
wire x_8207;
wire x_8208;
wire x_8209;
wire x_8210;
wire x_8211;
wire x_8212;
wire x_8213;
wire x_8214;
wire x_8215;
wire x_8216;
wire x_8217;
wire x_8218;
wire x_8219;
wire x_8220;
wire x_8221;
wire x_8222;
wire x_8223;
wire x_8224;
wire x_8225;
wire x_8226;
wire x_8227;
wire x_8228;
wire x_8229;
wire x_8230;
wire x_8231;
wire x_8232;
wire x_8233;
wire x_8234;
wire x_8235;
wire x_8236;
wire x_8237;
wire x_8238;
wire x_8239;
wire x_8240;
wire x_8241;
wire x_8242;
wire x_8243;
wire x_8244;
wire x_8245;
wire x_8246;
wire x_8247;
wire x_8248;
wire x_8249;
wire x_8250;
wire x_8251;
wire x_8252;
wire x_8253;
wire x_8254;
wire x_8255;
wire x_8256;
wire x_8257;
wire x_8258;
wire x_8259;
wire x_8260;
wire x_8261;
wire x_8262;
wire x_8263;
wire x_8264;
wire x_8265;
wire x_8266;
wire x_8267;
wire x_8268;
wire x_8269;
wire x_8270;
wire x_8271;
wire x_8272;
wire x_8273;
wire x_8274;
wire x_8275;
wire x_8276;
wire x_8277;
wire x_8278;
wire x_8279;
wire x_8280;
wire x_8281;
wire x_8282;
wire x_8283;
wire x_8284;
wire x_8285;
wire x_8286;
wire x_8287;
wire x_8288;
wire x_8289;
wire x_8290;
wire x_8291;
wire x_8292;
wire x_8293;
wire x_8294;
wire x_8295;
wire x_8296;
wire x_8297;
wire x_8298;
wire x_8299;
wire x_8300;
wire x_8301;
wire x_8302;
wire x_8303;
wire x_8304;
wire x_8305;
wire x_8306;
wire x_8307;
wire x_8308;
wire x_8309;
wire x_8310;
wire x_8311;
wire x_8312;
wire x_8313;
wire x_8314;
wire x_8315;
wire x_8316;
wire x_8317;
wire x_8318;
wire x_8319;
wire x_8320;
wire x_8321;
wire x_8322;
wire x_8323;
wire x_8324;
wire x_8325;
wire x_8326;
wire x_8327;
wire x_8328;
wire x_8329;
wire x_8330;
wire x_8331;
wire x_8332;
wire x_8333;
wire x_8334;
wire x_8335;
wire x_8336;
wire x_8337;
wire x_8338;
wire x_8339;
wire x_8340;
wire x_8341;
wire x_8342;
wire x_8343;
wire x_8344;
wire x_8345;
wire x_8346;
wire x_8347;
wire x_8348;
wire x_8349;
wire x_8350;
wire x_8351;
wire x_8352;
wire x_8353;
wire x_8354;
wire x_8355;
wire x_8356;
wire x_8357;
wire x_8358;
wire x_8359;
wire x_8360;
wire x_8361;
wire x_8362;
wire x_8363;
wire x_8364;
wire x_8365;
wire x_8366;
wire x_8367;
wire x_8368;
wire x_8369;
wire x_8370;
wire x_8371;
wire x_8372;
wire x_8373;
wire x_8374;
wire x_8375;
wire x_8376;
wire x_8377;
wire x_8378;
wire x_8379;
wire x_8380;
wire x_8381;
wire x_8382;
wire x_8383;
wire x_8384;
wire x_8385;
wire x_8386;
wire x_8387;
wire x_8388;
wire x_8389;
wire x_8390;
wire x_8391;
wire x_8392;
wire x_8393;
wire x_8394;
wire x_8395;
wire x_8396;
wire x_8397;
wire x_8398;
wire x_8399;
wire x_8400;
wire x_8401;
wire x_8402;
wire x_8403;
wire x_8404;
wire x_8405;
wire x_8406;
wire x_8407;
wire x_8408;
wire x_8409;
wire x_8410;
wire x_8411;
wire x_8412;
wire x_8413;
wire x_8414;
wire x_8415;
wire x_8416;
wire x_8417;
wire x_8418;
wire x_8419;
wire x_8420;
wire x_8421;
wire x_8422;
wire x_8423;
wire x_8424;
wire x_8425;
wire x_8426;
wire x_8427;
wire x_8428;
wire x_8429;
wire x_8430;
wire x_8431;
wire x_8432;
wire x_8433;
wire x_8434;
wire x_8435;
wire x_8436;
wire x_8437;
wire x_8438;
wire x_8439;
wire x_8440;
wire x_8441;
wire x_8442;
wire x_8443;
wire x_8444;
wire x_8445;
wire x_8446;
wire x_8447;
wire x_8448;
wire x_8449;
wire x_8450;
wire x_8451;
wire x_8452;
wire x_8453;
wire x_8454;
wire x_8455;
wire x_8456;
wire x_8457;
wire x_8458;
wire x_8459;
wire x_8460;
wire x_8461;
wire x_8462;
wire x_8463;
wire x_8464;
wire x_8465;
wire x_8466;
wire x_8467;
wire x_8468;
wire x_8469;
wire x_8470;
wire x_8471;
wire x_8472;
wire x_8473;
wire x_8474;
wire x_8475;
wire x_8476;
wire x_8477;
wire x_8478;
wire x_8479;
wire x_8480;
wire x_8481;
wire x_8482;
wire x_8483;
wire x_8484;
wire x_8485;
wire x_8486;
wire x_8487;
wire x_8488;
wire x_8489;
wire x_8490;
wire x_8491;
wire x_8492;
wire x_8493;
wire x_8494;
wire x_8495;
wire x_8496;
wire x_8497;
wire x_8498;
wire x_8499;
wire x_8500;
wire x_8501;
wire x_8502;
wire x_8503;
wire x_8504;
wire x_8505;
wire x_8506;
wire x_8507;
wire x_8508;
wire x_8509;
wire x_8510;
wire x_8511;
wire x_8512;
wire x_8513;
wire x_8514;
wire x_8515;
wire x_8516;
wire x_8517;
wire x_8518;
wire x_8519;
wire x_8520;
wire x_8521;
wire x_8522;
wire x_8523;
wire x_8524;
wire x_8525;
wire x_8526;
wire x_8527;
wire x_8528;
wire x_8529;
wire x_8530;
wire x_8531;
wire x_8532;
wire x_8533;
wire x_8534;
wire x_8535;
wire x_8536;
wire x_8537;
wire x_8538;
wire x_8539;
wire x_8540;
wire x_8541;
wire x_8542;
wire x_8543;
wire x_8544;
wire x_8545;
wire x_8546;
wire x_8547;
wire x_8548;
wire x_8549;
wire x_8550;
wire x_8551;
wire x_8552;
wire x_8553;
wire x_8554;
wire x_8555;
wire x_8556;
wire x_8557;
wire x_8558;
wire x_8559;
wire x_8560;
wire x_8561;
wire x_8562;
wire x_8563;
wire x_8564;
wire x_8565;
wire x_8566;
wire x_8567;
wire x_8568;
wire x_8569;
wire x_8570;
wire x_8571;
wire x_8572;
wire x_8573;
wire x_8574;
wire x_8575;
wire x_8576;
wire x_8577;
wire x_8578;
wire x_8579;
wire x_8580;
wire x_8581;
wire x_8582;
wire x_8583;
wire x_8584;
wire x_8585;
wire x_8586;
wire x_8587;
wire x_8588;
wire x_8589;
wire x_8590;
wire x_8591;
wire x_8592;
wire x_8593;
wire x_8594;
wire x_8595;
wire x_8596;
wire x_8597;
wire x_8598;
wire x_8599;
wire x_8600;
wire x_8601;
wire x_8602;
wire x_8603;
wire x_8604;
wire x_8605;
wire x_8606;
wire x_8607;
wire x_8608;
wire x_8609;
wire x_8610;
wire x_8611;
wire x_8612;
wire x_8613;
wire x_8614;
wire x_8615;
wire x_8616;
wire x_8617;
wire x_8618;
wire x_8619;
wire x_8620;
wire x_8621;
wire x_8622;
wire x_8623;
wire x_8624;
wire x_8625;
wire x_8626;
wire x_8627;
wire x_8628;
wire x_8629;
wire x_8630;
wire x_8631;
wire x_8632;
wire x_8633;
wire x_8634;
wire x_8635;
wire x_8636;
wire x_8637;
wire x_8638;
wire x_8639;
wire x_8640;
wire x_8641;
wire x_8642;
wire x_8643;
wire x_8644;
wire x_8645;
wire x_8646;
wire x_8647;
wire x_8648;
wire x_8649;
wire x_8650;
wire x_8651;
wire x_8652;
wire x_8653;
wire x_8654;
wire x_8655;
wire x_8656;
wire x_8657;
wire x_8658;
wire x_8659;
wire x_8660;
wire x_8661;
wire x_8662;
wire x_8663;
wire x_8664;
wire x_8665;
wire x_8666;
wire x_8667;
wire x_8668;
wire x_8669;
wire x_8670;
wire x_8671;
wire x_8672;
wire x_8673;
wire x_8674;
wire x_8675;
wire x_8676;
wire x_8677;
wire x_8678;
wire x_8679;
wire x_8680;
wire x_8681;
wire x_8682;
wire x_8683;
wire x_8684;
wire x_8685;
wire x_8686;
wire x_8687;
wire x_8688;
wire x_8689;
wire x_8690;
wire x_8691;
wire x_8692;
wire x_8693;
wire x_8694;
wire x_8695;
wire x_8696;
wire x_8697;
wire x_8698;
wire x_8699;
wire x_8700;
wire x_8701;
wire x_8702;
wire x_8703;
wire x_8704;
wire x_8705;
wire x_8706;
wire x_8707;
wire x_8708;
wire x_8709;
wire x_8710;
wire x_8711;
wire x_8712;
wire x_8713;
wire x_8714;
wire x_8715;
wire x_8716;
wire x_8717;
wire x_8718;
wire x_8719;
wire x_8720;
wire x_8721;
wire x_8722;
wire x_8723;
wire x_8724;
wire x_8725;
wire x_8726;
wire x_8727;
wire x_8728;
wire x_8729;
wire x_8730;
wire x_8731;
wire x_8732;
wire x_8733;
wire x_8734;
wire x_8735;
wire x_8736;
wire x_8737;
wire x_8738;
wire x_8739;
wire x_8740;
wire x_8741;
wire x_8742;
wire x_8743;
wire x_8744;
wire x_8745;
wire x_8746;
wire x_8747;
wire x_8748;
wire x_8749;
wire x_8750;
wire x_8751;
wire x_8752;
wire x_8753;
wire x_8754;
wire x_8755;
wire x_8756;
wire x_8757;
wire x_8758;
wire x_8759;
wire x_8760;
wire x_8761;
wire x_8762;
wire x_8763;
wire x_8764;
wire x_8765;
wire x_8766;
wire x_8767;
wire x_8768;
wire x_8769;
wire x_8770;
wire x_8771;
wire x_8772;
wire x_8773;
wire x_8774;
wire x_8775;
wire x_8776;
wire x_8777;
wire x_8778;
wire x_8779;
wire x_8780;
wire x_8781;
wire x_8782;
wire x_8783;
wire x_8784;
wire x_8785;
wire x_8786;
wire x_8787;
wire x_8788;
wire x_8789;
wire x_8790;
wire x_8791;
wire x_8792;
wire x_8793;
wire x_8794;
wire x_8795;
wire x_8796;
wire x_8797;
wire x_8798;
wire x_8799;
wire x_8800;
wire x_8801;
wire x_8802;
wire x_8803;
wire x_8804;
wire x_8805;
wire x_8806;
wire x_8807;
wire x_8808;
wire x_8809;
wire x_8810;
wire x_8811;
wire x_8812;
wire x_8813;
wire x_8814;
wire x_8815;
wire x_8816;
wire x_8817;
wire x_8818;
wire x_8819;
wire x_8820;
wire x_8821;
wire x_8822;
wire x_8823;
wire x_8824;
wire x_8825;
wire x_8826;
wire x_8827;
wire x_8828;
wire x_8829;
wire x_8830;
wire x_8831;
wire x_8832;
wire x_8833;
wire x_8834;
wire x_8835;
wire x_8836;
wire x_8837;
wire x_8838;
wire x_8839;
wire x_8840;
wire x_8841;
wire x_8842;
wire x_8843;
wire x_8844;
wire x_8845;
wire x_8846;
wire x_8847;
wire x_8848;
wire x_8849;
wire x_8850;
wire x_8851;
wire x_8852;
wire x_8853;
wire x_8854;
wire x_8855;
wire x_8856;
wire x_8857;
wire x_8858;
wire x_8859;
wire x_8860;
wire x_8861;
wire x_8862;
wire x_8863;
wire x_8864;
wire x_8865;
wire x_8866;
wire x_8867;
wire x_8868;
wire x_8869;
wire x_8870;
wire x_8871;
wire x_8872;
wire x_8873;
wire x_8874;
wire x_8875;
wire x_8876;
wire x_8877;
wire x_8878;
wire x_8879;
wire x_8880;
wire x_8881;
wire x_8882;
wire x_8883;
wire x_8884;
wire x_8885;
wire x_8886;
wire x_8887;
wire x_8888;
wire x_8889;
wire x_8890;
wire x_8891;
wire x_8892;
wire x_8893;
wire x_8894;
wire x_8895;
wire x_8896;
wire x_8897;
wire x_8898;
wire x_8899;
wire x_8900;
wire x_8901;
wire x_8902;
wire x_8903;
wire x_8904;
wire x_8905;
wire x_8906;
wire x_8907;
wire x_8908;
wire x_8909;
wire x_8910;
wire x_8911;
wire x_8912;
wire x_8913;
wire x_8914;
wire x_8915;
wire x_8916;
wire x_8917;
wire x_8918;
wire x_8919;
wire x_8920;
wire x_8921;
wire x_8922;
wire x_8923;
wire x_8924;
wire x_8925;
wire x_8926;
wire x_8927;
wire x_8928;
wire x_8929;
wire x_8930;
wire x_8931;
wire x_8932;
wire x_8933;
wire x_8934;
wire x_8935;
wire x_8936;
wire x_8937;
wire x_8938;
wire x_8939;
wire x_8940;
wire x_8941;
wire x_8942;
wire x_8943;
wire x_8944;
wire x_8945;
wire x_8946;
wire x_8947;
wire x_8948;
wire x_8949;
wire x_8950;
wire x_8951;
wire x_8952;
wire x_8953;
wire x_8954;
wire x_8955;
wire x_8956;
wire x_8957;
wire x_8958;
wire x_8959;
wire x_8960;
wire x_8961;
wire x_8962;
wire x_8963;
wire x_8964;
wire x_8965;
wire x_8966;
wire x_8967;
wire x_8968;
wire x_8969;
wire x_8970;
wire x_8971;
wire x_8972;
wire x_8973;
wire x_8974;
wire x_8975;
wire x_8976;
wire x_8977;
wire x_8978;
wire x_8979;
wire x_8980;
wire x_8981;
wire x_8982;
wire x_8983;
wire x_8984;
wire x_8985;
wire x_8986;
wire x_8987;
wire x_8988;
wire x_8989;
wire x_8990;
wire x_8991;
wire x_8992;
wire x_8993;
wire x_8994;
wire x_8995;
wire x_8996;
wire x_8997;
wire x_8998;
wire x_8999;
wire x_9000;
wire x_9001;
wire x_9002;
wire x_9003;
wire x_9004;
wire x_9005;
wire x_9006;
wire x_9007;
wire x_9008;
wire x_9009;
wire x_9010;
wire x_9011;
wire x_9012;
wire x_9013;
wire x_9014;
wire x_9015;
wire x_9016;
wire x_9017;
wire x_9018;
wire x_9019;
wire x_9020;
wire x_9021;
wire x_9022;
wire x_9023;
wire x_9024;
wire x_9025;
wire x_9026;
wire x_9027;
wire x_9028;
wire x_9029;
wire x_9030;
wire x_9031;
wire x_9032;
wire x_9033;
wire x_9034;
wire x_9035;
wire x_9036;
wire x_9037;
wire x_9038;
wire x_9039;
wire x_9040;
wire x_9041;
wire x_9042;
wire x_9043;
wire x_9044;
wire x_9045;
wire x_9046;
wire x_9047;
wire x_9048;
wire x_9049;
wire x_9050;
wire x_9051;
wire x_9052;
wire x_9053;
wire x_9054;
wire x_9055;
wire x_9056;
wire x_9057;
wire x_9058;
wire x_9059;
wire x_9060;
wire x_9061;
wire x_9062;
wire x_9063;
wire x_9064;
wire x_9065;
wire x_9066;
wire x_9067;
wire x_9068;
wire x_9069;
wire x_9070;
wire x_9071;
wire x_9072;
wire x_9073;
wire x_9074;
wire x_9075;
wire x_9076;
wire x_9077;
wire x_9078;
wire x_9079;
wire x_9080;
wire x_9081;
wire x_9082;
wire x_9083;
wire x_9084;
wire x_9085;
wire x_9086;
wire x_9087;
wire x_9088;
wire x_9089;
wire x_9090;
wire x_9091;
wire x_9092;
wire x_9093;
wire x_9094;
wire x_9095;
wire x_9096;
wire x_9097;
wire x_9098;
wire x_9099;
wire x_9100;
wire x_9101;
wire x_9102;
wire x_9103;
wire x_9104;
wire x_9105;
wire x_9106;
wire x_9107;
wire x_9108;
wire x_9109;
wire x_9110;
wire x_9111;
wire x_9112;
wire x_9113;
wire x_9114;
wire x_9115;
wire x_9116;
wire x_9117;
wire x_9118;
wire x_9119;
wire x_9120;
wire x_9121;
wire x_9122;
wire x_9123;
wire x_9124;
wire x_9125;
wire x_9126;
wire x_9127;
wire x_9128;
wire x_9129;
wire x_9130;
wire x_9131;
wire x_9132;
wire x_9133;
wire x_9134;
wire x_9135;
wire x_9136;
wire x_9137;
wire x_9138;
wire x_9139;
wire x_9140;
wire x_9141;
wire x_9142;
wire x_9143;
wire x_9144;
wire x_9145;
wire x_9146;
wire x_9147;
wire x_9148;
wire x_9149;
wire x_9150;
wire x_9151;
wire x_9152;
wire x_9153;
wire x_9154;
wire x_9155;
wire x_9156;
wire x_9157;
wire x_9158;
wire x_9159;
wire x_9160;
wire x_9161;
wire x_9162;
wire x_9163;
wire x_9164;
wire x_9165;
wire x_9166;
wire x_9167;
wire x_9168;
wire x_9169;
wire x_9170;
wire x_9171;
wire x_9172;
wire x_9173;
wire x_9174;
wire x_9175;
wire x_9176;
wire x_9177;
wire x_9178;
wire x_9179;
wire x_9180;
wire x_9181;
wire x_9182;
wire x_9183;
wire x_9184;
wire x_9185;
wire x_9186;
wire x_9187;
wire x_9188;
wire x_9189;
wire x_9190;
wire x_9191;
wire x_9192;
wire x_9193;
wire x_9194;
wire x_9195;
wire x_9196;
wire x_9197;
wire x_9198;
wire x_9199;
wire x_9200;
wire x_9201;
wire x_9202;
wire x_9203;
wire x_9204;
wire x_9205;
wire x_9206;
wire x_9207;
wire x_9208;
wire x_9209;
wire x_9210;
wire x_9211;
wire x_9212;
wire x_9213;
wire x_9214;
wire x_9215;
wire x_9216;
wire x_9217;
wire x_9218;
wire x_9219;
wire x_9220;
wire x_9221;
wire x_9222;
wire x_9223;
wire x_9224;
wire x_9225;
wire x_9226;
wire x_9227;
wire x_9228;
wire x_9229;
wire x_9230;
wire x_9231;
wire x_9232;
wire x_9233;
wire x_9234;
wire x_9235;
wire x_9236;
wire x_9237;
wire x_9238;
wire x_9239;
wire x_9240;
wire x_9241;
wire x_9242;
wire x_9243;
wire x_9244;
wire x_9245;
wire x_9246;
wire x_9247;
wire x_9248;
wire x_9249;
wire x_9250;
wire x_9251;
wire x_9252;
wire x_9253;
wire x_9254;
wire x_9255;
wire x_9256;
wire x_9257;
wire x_9258;
wire x_9259;
wire x_9260;
wire x_9261;
wire x_9262;
wire x_9263;
wire x_9264;
wire x_9265;
wire x_9266;
wire x_9267;
wire x_9268;
wire x_9269;
wire x_9270;
wire x_9271;
wire x_9272;
wire x_9273;
wire x_9274;
wire x_9275;
wire x_9276;
wire x_9277;
wire x_9278;
wire x_9279;
wire x_9280;
wire x_9281;
wire x_9282;
wire x_9283;
wire x_9284;
wire x_9285;
wire x_9286;
wire x_9287;
wire x_9288;
wire x_9289;
wire x_9290;
wire x_9291;
wire x_9292;
wire x_9293;
wire x_9294;
wire x_9295;
wire x_9296;
wire x_9297;
wire x_9298;
wire x_9299;
wire x_9300;
wire x_9301;
wire x_9302;
wire x_9303;
wire x_9304;
wire x_9305;
wire x_9306;
wire x_9307;
wire x_9308;
wire x_9309;
wire x_9310;
wire x_9311;
wire x_9312;
wire x_9313;
wire x_9314;
wire x_9315;
wire x_9316;
wire x_9317;
wire x_9318;
wire x_9319;
wire x_9320;
wire x_9321;
wire x_9322;
wire x_9323;
wire x_9324;
wire x_9325;
wire x_9326;
wire x_9327;
wire x_9328;
wire x_9329;
wire x_9330;
wire x_9331;
wire x_9332;
wire x_9333;
wire x_9334;
wire x_9335;
wire x_9336;
wire x_9337;
wire x_9338;
wire x_9339;
wire x_9340;
wire x_9341;
wire x_9342;
wire x_9343;
wire x_9344;
wire x_9345;
wire x_9346;
wire x_9347;
wire x_9348;
wire x_9349;
wire x_9350;
wire x_9351;
wire x_9352;
wire x_9353;
wire x_9354;
wire x_9355;
wire x_9356;
wire x_9357;
wire x_9358;
wire x_9359;
wire x_9360;
wire x_9361;
wire x_9362;
wire x_9363;
wire x_9364;
wire x_9365;
wire x_9366;
wire x_9367;
wire x_9368;
wire x_9369;
wire x_9370;
wire x_9371;
wire x_9372;
wire x_9373;
wire x_9374;
wire x_9375;
wire x_9376;
wire x_9377;
wire x_9378;
wire x_9379;
wire x_9380;
wire x_9381;
wire x_9382;
wire x_9383;
wire x_9384;
wire x_9385;
wire x_9386;
wire x_9387;
wire x_9388;
wire x_9389;
wire x_9390;
wire x_9391;
wire x_9392;
wire x_9393;
wire x_9394;
wire x_9395;
wire x_9396;
wire x_9397;
wire x_9398;
wire x_9399;
wire x_9400;
wire x_9401;
wire x_9402;
wire x_9403;
wire x_9404;
wire x_9405;
wire x_9406;
wire x_9407;
wire x_9408;
wire x_9409;
wire x_9410;
wire x_9411;
wire x_9412;
wire x_9413;
wire x_9414;
wire x_9415;
wire x_9416;
wire x_9417;
wire x_9418;
wire x_9419;
wire x_9420;
wire x_9421;
wire x_9422;
wire x_9423;
wire x_9424;
wire x_9425;
wire x_9426;
wire x_9427;
wire x_9428;
wire x_9429;
wire x_9430;
wire x_9431;
wire x_9432;
wire x_9433;
wire x_9434;
wire x_9435;
wire x_9436;
wire x_9437;
wire x_9438;
wire x_9439;
wire x_9440;
wire x_9441;
wire x_9442;
wire x_9443;
wire x_9444;
wire x_9445;
wire x_9446;
wire x_9447;
wire x_9448;
wire x_9449;
wire x_9450;
wire x_9451;
wire x_9452;
wire x_9453;
wire x_9454;
wire x_9455;
wire x_9456;
wire x_9457;
wire x_9458;
wire x_9459;
wire x_9460;
wire x_9461;
wire x_9462;
wire x_9463;
wire x_9464;
wire x_9465;
wire x_9466;
wire x_9467;
wire x_9468;
wire x_9469;
wire x_9470;
wire x_9471;
wire x_9472;
wire x_9473;
wire x_9474;
wire x_9475;
wire x_9476;
wire x_9477;
wire x_9478;
wire x_9479;
wire x_9480;
wire x_9481;
wire x_9482;
wire x_9483;
wire x_9484;
wire x_9485;
wire x_9486;
wire x_9487;
wire x_9488;
wire x_9489;
wire x_9490;
wire x_9491;
wire x_9492;
wire x_9493;
wire x_9494;
wire x_9495;
wire x_9496;
wire x_9497;
wire x_9498;
wire x_9499;
wire x_9500;
wire x_9501;
wire x_9502;
wire x_9503;
wire x_9504;
wire x_9505;
wire x_9506;
wire x_9507;
wire x_9508;
wire x_9509;
wire x_9510;
wire x_9511;
wire x_9512;
wire x_9513;
wire x_9514;
wire x_9515;
wire x_9516;
wire x_9517;
wire x_9518;
wire x_9519;
wire x_9520;
wire x_9521;
wire x_9522;
wire x_9523;
wire x_9524;
wire x_9525;
wire x_9526;
wire x_9527;
wire x_9528;
wire x_9529;
wire x_9530;
wire x_9531;
wire x_9532;
wire x_9533;
wire x_9534;
wire x_9535;
wire x_9536;
wire x_9537;
wire x_9538;
wire x_9539;
wire x_9540;
wire x_9541;
wire x_9542;
wire x_9543;
wire x_9544;
wire x_9545;
wire x_9546;
wire x_9547;
wire x_9548;
wire x_9549;
wire x_9550;
wire x_9551;
wire x_9552;
wire x_9553;
wire x_9554;
wire x_9555;
wire x_9556;
wire x_9557;
wire x_9558;
wire x_9559;
wire x_9560;
wire x_9561;
wire x_9562;
wire x_9563;
wire x_9564;
wire x_9565;
wire x_9566;
wire x_9567;
wire x_9568;
wire x_9569;
wire x_9570;
wire x_9571;
wire x_9572;
wire x_9573;
wire x_9574;
wire x_9575;
wire x_9576;
wire x_9577;
wire x_9578;
wire x_9579;
wire x_9580;
wire x_9581;
wire x_9582;
wire x_9583;
wire x_9584;
wire x_9585;
wire x_9586;
wire x_9587;
wire x_9588;
wire x_9589;
wire x_9590;
wire x_9591;
wire x_9592;
wire x_9593;
wire x_9594;
wire x_9595;
wire x_9596;
wire x_9597;
wire x_9598;
wire x_9599;
wire x_9600;
wire x_9601;
wire x_9602;
wire x_9603;
wire x_9604;
wire x_9605;
wire x_9606;
wire x_9607;
wire x_9608;
wire x_9609;
wire x_9610;
wire x_9611;
wire x_9612;
wire x_9613;
wire x_9614;
wire x_9615;
wire x_9616;
wire x_9617;
wire x_9618;
wire x_9619;
wire x_9620;
wire x_9621;
wire x_9622;
wire x_9623;
wire x_9624;
wire x_9625;
wire x_9626;
wire x_9627;
wire x_9628;
wire x_9629;
wire x_9630;
wire x_9631;
wire x_9632;
wire x_9633;
wire x_9634;
wire x_9635;
wire x_9636;
wire x_9637;
wire x_9638;
wire x_9639;
wire x_9640;
wire x_9641;
wire x_9642;
wire x_9643;
wire x_9644;
wire x_9645;
wire x_9646;
wire x_9647;
wire x_9648;
wire x_9649;
wire x_9650;
wire x_9651;
wire x_9652;
wire x_9653;
wire x_9654;
wire x_9655;
wire x_9656;
wire x_9657;
wire x_9658;
wire x_9659;
wire x_9660;
wire x_9661;
wire x_9662;
wire x_9663;
wire x_9664;
wire x_9665;
wire x_9666;
wire x_9667;
wire x_9668;
wire x_9669;
wire x_9670;
wire x_9671;
wire x_9672;
wire x_9673;
wire x_9674;
wire x_9675;
wire x_9676;
wire x_9677;
wire x_9678;
wire x_9679;
wire x_9680;
wire x_9681;
wire x_9682;
wire x_9683;
wire x_9684;
wire x_9685;
wire x_9686;
wire x_9687;
wire x_9688;
wire x_9689;
wire x_9690;
wire x_9691;
wire x_9692;
wire x_9693;
wire x_9694;
wire x_9695;
wire x_9696;
wire x_9697;
wire x_9698;
wire x_9699;
wire x_9700;
wire x_9701;
wire x_9702;
wire x_9703;
wire x_9704;
wire x_9705;
wire x_9706;
wire x_9707;
wire x_9708;
wire x_9709;
wire x_9710;
wire x_9711;
wire x_9712;
wire x_9713;
wire x_9714;
wire x_9715;
wire x_9716;
wire x_9717;
wire x_9718;
wire x_9719;
wire x_9720;
wire x_9721;
wire x_9722;
wire x_9723;
wire x_9724;
wire x_9725;
wire x_9726;
wire x_9727;
wire x_9728;
wire x_9729;
wire x_9730;
wire x_9731;
wire x_9732;
wire x_9733;
wire x_9734;
wire x_9735;
wire x_9736;
wire x_9737;
wire x_9738;
wire x_9739;
wire x_9740;
wire x_9741;
wire x_9742;
wire x_9743;
wire x_9744;
wire x_9745;
wire x_9746;
wire x_9747;
wire x_9748;
wire x_9749;
wire x_9750;
wire x_9751;
wire x_9752;
wire x_9753;
wire x_9754;
wire x_9755;
wire x_9756;
wire x_9757;
wire x_9758;
wire x_9759;
wire x_9760;
wire x_9761;
wire x_9762;
wire x_9763;
wire x_9764;
wire x_9765;
wire x_9766;
wire x_9767;
wire x_9768;
wire x_9769;
wire x_9770;
wire x_9771;
wire x_9772;
wire x_9773;
wire x_9774;
wire x_9775;
wire x_9776;
wire x_9777;
wire x_9778;
wire x_9779;
wire x_9780;
wire x_9781;
wire x_9782;
wire x_9783;
wire x_9784;
wire x_9785;
wire x_9786;
wire x_9787;
wire x_9788;
wire x_9789;
wire x_9790;
wire x_9791;
wire x_9792;
wire x_9793;
wire x_9794;
wire x_9795;
wire x_9796;
wire x_9797;
wire x_9798;
wire x_9799;
wire x_9800;
wire x_9801;
wire x_9802;
wire x_9803;
wire x_9804;
wire x_9805;
wire x_9806;
wire x_9807;
wire x_9808;
wire x_9809;
wire x_9810;
wire x_9811;
wire x_9812;
wire x_9813;
wire x_9814;
wire x_9815;
wire x_9816;
wire x_9817;
wire x_9818;
wire x_9819;
wire x_9820;
wire x_9821;
wire x_9822;
wire x_9823;
wire x_9824;
wire x_9825;
wire x_9826;
wire x_9827;
wire x_9828;
wire x_9829;
wire x_9830;
wire x_9831;
wire x_9832;
wire x_9833;
wire x_9834;
wire x_9835;
wire x_9836;
wire x_9837;
wire x_9838;
wire x_9839;
wire x_9840;
wire x_9841;
wire x_9842;
wire x_9843;
wire x_9844;
wire x_9845;
wire x_9846;
wire x_9847;
wire x_9848;
wire x_9849;
wire x_9850;
wire x_9851;
wire x_9852;
wire x_9853;
wire x_9854;
wire x_9855;
wire x_9856;
wire x_9857;
wire x_9858;
wire x_9859;
wire x_9860;
wire x_9861;
wire x_9862;
wire x_9863;
wire x_9864;
wire x_9865;
wire x_9866;
wire x_9867;
wire x_9868;
wire x_9869;
wire x_9870;
wire x_9871;
wire x_9872;
wire x_9873;
wire x_9874;
wire x_9875;
wire x_9876;
wire x_9877;
wire x_9878;
wire x_9879;
wire x_9880;
wire x_9881;
wire x_9882;
wire x_9883;
wire x_9884;
wire x_9885;
wire x_9886;
wire x_9887;
wire x_9888;
wire x_9889;
wire x_9890;
wire x_9891;
wire x_9892;
wire x_9893;
wire x_9894;
wire x_9895;
wire x_9896;
wire x_9897;
wire x_9898;
wire x_9899;
wire x_9900;
wire x_9901;
wire x_9902;
wire x_9903;
wire x_9904;
wire x_9905;
wire x_9906;
wire x_9907;
wire x_9908;
wire x_9909;
wire x_9910;
wire x_9911;
wire x_9912;
wire x_9913;
wire x_9914;
wire x_9915;
wire x_9916;
wire x_9917;
wire x_9918;
wire x_9919;
wire x_9920;
wire x_9921;
wire x_9922;
wire x_9923;
wire x_9924;
wire x_9925;
wire x_9926;
wire x_9927;
wire x_9928;
wire x_9929;
wire x_9930;
wire x_9931;
wire x_9932;
wire x_9933;
wire x_9934;
wire x_9935;
wire x_9936;
wire x_9937;
wire x_9938;
wire x_9939;
wire x_9940;
wire x_9941;
wire x_9942;
wire x_9943;
wire x_9944;
wire x_9945;
wire x_9946;
wire x_9947;
wire x_9948;
wire x_9949;
wire x_9950;
wire x_9951;
wire x_9952;
wire x_9953;
wire x_9954;
wire x_9955;
wire x_9956;
wire x_9957;
wire x_9958;
wire x_9959;
wire x_9960;
wire x_9961;
wire x_9962;
wire x_9963;
wire x_9964;
wire x_9965;
wire x_9966;
wire x_9967;
wire x_9968;
wire x_9969;
wire x_9970;
wire x_9971;
wire x_9972;
wire x_9973;
wire x_9974;
wire x_9975;
wire x_9976;
wire x_9977;
wire x_9978;
wire x_9979;
wire x_9980;
wire x_9981;
wire x_9982;
wire x_9983;
wire x_9984;
wire x_9985;
wire x_9986;
wire x_9987;
wire x_9988;
wire x_9989;
wire x_9990;
wire x_9991;
wire x_9992;
wire x_9993;
wire x_9994;
wire x_9995;
wire x_9996;
wire x_9997;
wire x_9998;
wire x_9999;
wire x_10000;
wire x_10001;
wire x_10002;
wire x_10003;
wire x_10004;
wire x_10005;
wire x_10006;
wire x_10007;
wire x_10008;
wire x_10009;
wire x_10010;
wire x_10011;
wire x_10012;
wire x_10013;
wire x_10014;
wire x_10015;
wire x_10016;
wire x_10017;
wire x_10018;
wire x_10019;
wire x_10020;
wire x_10021;
wire x_10022;
wire x_10023;
wire x_10024;
wire x_10025;
wire x_10026;
wire x_10027;
wire x_10028;
wire x_10029;
wire x_10030;
wire x_10031;
wire x_10032;
wire x_10033;
wire x_10034;
wire x_10035;
wire x_10036;
wire x_10037;
wire x_10038;
wire x_10039;
wire x_10040;
wire x_10041;
wire x_10042;
wire x_10043;
wire x_10044;
wire x_10045;
wire x_10046;
wire x_10047;
wire x_10048;
wire x_10049;
wire x_10050;
wire x_10051;
wire x_10052;
wire x_10053;
wire x_10054;
wire x_10055;
wire x_10056;
wire x_10057;
wire x_10058;
wire x_10059;
wire x_10060;
wire x_10061;
wire x_10062;
wire x_10063;
wire x_10064;
wire x_10065;
wire x_10066;
wire x_10067;
wire x_10068;
wire x_10069;
wire x_10070;
wire x_10071;
wire x_10072;
wire x_10073;
wire x_10074;
wire x_10075;
wire x_10076;
wire x_10077;
wire x_10078;
wire x_10079;
wire x_10080;
wire x_10081;
wire x_10082;
wire x_10083;
wire x_10084;
wire x_10085;
wire x_10086;
wire x_10087;
wire x_10088;
wire x_10089;
wire x_10090;
wire x_10091;
wire x_10092;
wire x_10093;
wire x_10094;
wire x_10095;
wire x_10096;
wire x_10097;
wire x_10098;
wire x_10099;
wire x_10100;
wire x_10101;
wire x_10102;
wire x_10103;
wire x_10104;
wire x_10105;
wire x_10106;
wire x_10107;
wire x_10108;
wire x_10109;
wire x_10110;
wire x_10111;
wire x_10112;
wire x_10113;
wire x_10114;
wire x_10115;
wire x_10116;
wire x_10117;
wire x_10118;
wire x_10119;
wire x_10120;
wire x_10121;
wire x_10122;
wire x_10123;
wire x_10124;
wire x_10125;
wire x_10126;
wire x_10127;
wire x_10128;
wire x_10129;
wire x_10130;
wire x_10131;
wire x_10132;
wire x_10133;
wire x_10134;
wire x_10135;
wire x_10136;
wire x_10137;
wire x_10138;
wire x_10139;
wire x_10140;
wire x_10141;
wire x_10142;
wire x_10143;
wire x_10144;
wire x_10145;
wire x_10146;
wire x_10147;
wire x_10148;
wire x_10149;
wire x_10150;
wire x_10151;
wire x_10152;
wire x_10153;
wire x_10154;
wire x_10155;
wire x_10156;
wire x_10157;
wire x_10158;
wire x_10159;
wire x_10160;
wire x_10161;
wire x_10162;
wire x_10163;
wire x_10164;
wire x_10165;
wire x_10166;
wire x_10167;
wire x_10168;
wire x_10169;
wire x_10170;
wire x_10171;
wire x_10172;
wire x_10173;
wire x_10174;
wire x_10175;
wire x_10176;
wire x_10177;
wire x_10178;
wire x_10179;
wire x_10180;
wire x_10181;
wire x_10182;
wire x_10183;
wire x_10184;
wire x_10185;
wire x_10186;
wire x_10187;
wire x_10188;
wire x_10189;
wire x_10190;
wire x_10191;
wire x_10192;
wire x_10193;
wire x_10194;
wire x_10195;
wire x_10196;
wire x_10197;
wire x_10198;
wire x_10199;
wire x_10200;
wire x_10201;
wire x_10202;
wire x_10203;
wire x_10204;
wire x_10205;
wire x_10206;
wire x_10207;
wire x_10208;
wire x_10209;
wire x_10210;
wire x_10211;
wire x_10212;
wire x_10213;
wire x_10214;
wire x_10215;
wire x_10216;
wire x_10217;
wire x_10218;
wire x_10219;
wire x_10220;
wire x_10221;
wire x_10222;
wire x_10223;
wire x_10224;
wire x_10225;
wire x_10226;
wire x_10227;
wire x_10228;
wire x_10229;
wire x_10230;
wire x_10231;
wire x_10232;
wire x_10233;
wire x_10234;
wire x_10235;
wire x_10236;
wire x_10237;
wire x_10238;
wire x_10239;
wire x_10240;
wire x_10241;
wire x_10242;
wire x_10243;
wire x_10244;
wire x_10245;
wire x_10246;
wire x_10247;
wire x_10248;
wire x_10249;
wire x_10250;
wire x_10251;
wire x_10252;
wire x_10253;
wire x_10254;
wire x_10255;
wire x_10256;
wire x_10257;
wire x_10258;
wire x_10259;
wire x_10260;
wire x_10261;
wire x_10262;
wire x_10263;
wire x_10264;
wire x_10265;
wire x_10266;
wire x_10267;
wire x_10268;
wire x_10269;
wire x_10270;
wire x_10271;
wire x_10272;
wire x_10273;
wire x_10274;
wire x_10275;
wire x_10276;
wire x_10277;
wire x_10278;
wire x_10279;
wire x_10280;
wire x_10281;
wire x_10282;
wire x_10283;
wire x_10284;
wire x_10285;
wire x_10286;
wire x_10287;
wire x_10288;
wire x_10289;
wire x_10290;
wire x_10291;
wire x_10292;
wire x_10293;
wire x_10294;
wire x_10295;
wire x_10296;
wire x_10297;
wire x_10298;
wire x_10299;
wire x_10300;
wire x_10301;
wire x_10302;
wire x_10303;
wire x_10304;
wire x_10305;
wire x_10306;
wire x_10307;
wire x_10308;
wire x_10309;
wire x_10310;
wire x_10311;
wire x_10312;
wire x_10313;
wire x_10314;
wire x_10315;
wire x_10316;
wire x_10317;
wire x_10318;
wire x_10319;
wire x_10320;
wire x_10321;
wire x_10322;
wire x_10323;
wire x_10324;
wire x_10325;
wire x_10326;
wire x_10327;
wire x_10328;
wire x_10329;
wire x_10330;
wire x_10331;
wire x_10332;
wire x_10333;
wire x_10334;
wire x_10335;
wire x_10336;
wire x_10337;
wire x_10338;
wire x_10339;
wire x_10340;
wire x_10341;
wire x_10342;
wire x_10343;
wire x_10344;
wire x_10345;
wire x_10346;
wire x_10347;
wire x_10348;
wire x_10349;
wire x_10350;
wire x_10351;
wire x_10352;
wire x_10353;
wire x_10354;
wire x_10355;
wire x_10356;
wire x_10357;
wire x_10358;
wire x_10359;
wire x_10360;
wire x_10361;
wire x_10362;
wire x_10363;
wire x_10364;
wire x_10365;
wire x_10366;
wire x_10367;
wire x_10368;
wire x_10369;
wire x_10370;
wire x_10371;
wire x_10372;
wire x_10373;
wire x_10374;
wire x_10375;
wire x_10376;
wire x_10377;
wire x_10378;
wire x_10379;
wire x_10380;
wire x_10381;
wire x_10382;
wire x_10383;
wire x_10384;
wire x_10385;
wire x_10386;
wire x_10387;
wire x_10388;
wire x_10389;
wire x_10390;
wire x_10391;
wire x_10392;
wire x_10393;
wire x_10394;
wire x_10395;
wire x_10396;
wire x_10397;
wire x_10398;
wire x_10399;
wire x_10400;
wire x_10401;
wire x_10402;
wire x_10403;
wire x_10404;
wire x_10405;
wire x_10406;
wire x_10407;
wire x_10408;
wire x_10409;
wire x_10410;
wire x_10411;
wire x_10412;
wire x_10413;
wire x_10414;
wire x_10415;
wire x_10416;
wire x_10417;
wire x_10418;
wire x_10419;
wire x_10420;
wire x_10421;
wire x_10422;
wire x_10423;
wire x_10424;
wire x_10425;
wire x_10426;
wire x_10427;
wire x_10428;
wire x_10429;
wire x_10430;
wire x_10431;
wire x_10432;
wire x_10433;
wire x_10434;
wire x_10435;
wire x_10436;
wire x_10437;
wire x_10438;
wire x_10439;
wire x_10440;
wire x_10441;
wire x_10442;
wire x_10443;
wire x_10444;
wire x_10445;
wire x_10446;
wire x_10447;
wire x_10448;
wire x_10449;
wire x_10450;
wire x_10451;
wire x_10452;
wire x_10453;
wire x_10454;
wire x_10455;
wire x_10456;
wire x_10457;
wire x_10458;
wire x_10459;
wire x_10460;
wire x_10461;
wire x_10462;
wire x_10463;
wire x_10464;
wire x_10465;
wire x_10466;
wire x_10467;
wire x_10468;
wire x_10469;
wire x_10470;
wire x_10471;
wire x_10472;
wire x_10473;
wire x_10474;
wire x_10475;
wire x_10476;
wire x_10477;
wire x_10478;
wire x_10479;
wire x_10480;
wire x_10481;
wire x_10482;
wire x_10483;
wire x_10484;
wire x_10485;
wire x_10486;
wire x_10487;
wire x_10488;
wire x_10489;
wire x_10490;
wire x_10491;
wire x_10492;
wire x_10493;
wire x_10494;
wire x_10495;
wire x_10496;
wire x_10497;
wire x_10498;
wire x_10499;
wire x_10500;
wire x_10501;
wire x_10502;
wire x_10503;
wire x_10504;
wire x_10505;
wire x_10506;
wire x_10507;
wire x_10508;
wire x_10509;
wire x_10510;
wire x_10511;
wire x_10512;
wire x_10513;
wire x_10514;
wire x_10515;
wire x_10516;
wire x_10517;
wire x_10518;
wire x_10519;
wire x_10520;
wire x_10521;
wire x_10522;
wire x_10523;
wire x_10524;
wire x_10525;
wire x_10526;
wire x_10527;
wire x_10528;
wire x_10529;
wire x_10530;
wire x_10531;
wire x_10532;
wire x_10533;
wire x_10534;
wire x_10535;
wire x_10536;
wire x_10537;
wire x_10538;
wire x_10539;
wire x_10540;
wire x_10541;
wire x_10542;
wire x_10543;
wire x_10544;
wire x_10545;
wire x_10546;
wire x_10547;
wire x_10548;
wire x_10549;
wire x_10550;
wire x_10551;
wire x_10552;
wire x_10553;
wire x_10554;
wire x_10555;
wire x_10556;
wire x_10557;
wire x_10558;
wire x_10559;
wire x_10560;
wire x_10561;
wire x_10562;
wire x_10563;
wire x_10564;
wire x_10565;
wire x_10566;
wire x_10567;
wire x_10568;
wire x_10569;
wire x_10570;
wire x_10571;
wire x_10572;
wire x_10573;
wire x_10574;
wire x_10575;
wire x_10576;
wire x_10577;
wire x_10578;
wire x_10579;
wire x_10580;
wire x_10581;
wire x_10582;
wire x_10583;
wire x_10584;
wire x_10585;
wire x_10586;
wire x_10587;
wire x_10588;
wire x_10589;
wire x_10590;
wire x_10591;
wire x_10592;
wire x_10593;
wire x_10594;
wire x_10595;
wire x_10596;
wire x_10597;
wire x_10598;
wire x_10599;
wire x_10600;
wire x_10601;
wire x_10602;
wire x_10603;
wire x_10604;
wire x_10605;
wire x_10606;
wire x_10607;
wire x_10608;
wire x_10609;
wire x_10610;
wire x_10611;
wire x_10612;
wire x_10613;
wire x_10614;
wire x_10615;
wire x_10616;
wire x_10617;
wire x_10618;
wire x_10619;
wire x_10620;
wire x_10621;
wire x_10622;
wire x_10623;
wire x_10624;
wire x_10625;
wire x_10626;
wire x_10627;
wire x_10628;
wire x_10629;
wire x_10630;
wire x_10631;
wire x_10632;
wire x_10633;
wire x_10634;
wire x_10635;
wire x_10636;
wire x_10637;
wire x_10638;
wire x_10639;
wire x_10640;
wire x_10641;
wire x_10642;
wire x_10643;
wire x_10644;
wire x_10645;
wire x_10646;
wire x_10647;
wire x_10648;
wire x_10649;
wire x_10650;
wire x_10651;
wire x_10652;
wire x_10653;
wire x_10654;
wire x_10655;
wire x_10656;
wire x_10657;
wire x_10658;
wire x_10659;
wire x_10660;
wire x_10661;
wire x_10662;
wire x_10663;
wire x_10664;
wire x_10665;
wire x_10666;
wire x_10667;
wire x_10668;
wire x_10669;
wire x_10670;
wire x_10671;
wire x_10672;
wire x_10673;
wire x_10674;
wire x_10675;
wire x_10676;
wire x_10677;
wire x_10678;
wire x_10679;
wire x_10680;
wire x_10681;
wire x_10682;
wire x_10683;
wire x_10684;
wire x_10685;
wire x_10686;
wire x_10687;
wire x_10688;
wire x_10689;
wire x_10690;
wire x_10691;
wire x_10692;
wire x_10693;
wire x_10694;
wire x_10695;
wire x_10696;
wire x_10697;
wire x_10698;
wire x_10699;
wire x_10700;
wire x_10701;
wire x_10702;
wire x_10703;
wire x_10704;
wire x_10705;
wire x_10706;
wire x_10707;
wire x_10708;
wire x_10709;
wire x_10710;
wire x_10711;
wire x_10712;
wire x_10713;
wire x_10714;
wire x_10715;
wire x_10716;
wire x_10717;
wire x_10718;
wire x_10719;
wire x_10720;
wire x_10721;
wire x_10722;
wire x_10723;
wire x_10724;
wire x_10725;
wire x_10726;
wire x_10727;
wire x_10728;
wire x_10729;
wire x_10730;
wire x_10731;
wire x_10732;
wire x_10733;
wire x_10734;
wire x_10735;
wire x_10736;
wire x_10737;
wire x_10738;
wire x_10739;
wire x_10740;
wire x_10741;
wire x_10742;
wire x_10743;
wire x_10744;
wire x_10745;
wire x_10746;
wire x_10747;
wire x_10748;
wire x_10749;
wire x_10750;
wire x_10751;
wire x_10752;
wire x_10753;
wire x_10754;
wire x_10755;
wire x_10756;
wire x_10757;
wire x_10758;
wire x_10759;
wire x_10760;
wire x_10761;
wire x_10762;
wire x_10763;
wire x_10764;
wire x_10765;
wire x_10766;
wire x_10767;
wire x_10768;
wire x_10769;
wire x_10770;
wire x_10771;
wire x_10772;
wire x_10773;
wire x_10774;
wire x_10775;
wire x_10776;
wire x_10777;
wire x_10778;
wire x_10779;
wire x_10780;
wire x_10781;
wire x_10782;
wire x_10783;
wire x_10784;
wire x_10785;
wire x_10786;
wire x_10787;
wire x_10788;
wire x_10789;
wire x_10790;
wire x_10791;
wire x_10792;
wire x_10793;
wire x_10794;
wire x_10795;
wire x_10796;
wire x_10797;
wire x_10798;
wire x_10799;
wire x_10800;
wire x_10801;
wire x_10802;
wire x_10803;
wire x_10804;
wire x_10805;
wire x_10806;
wire x_10807;
wire x_10808;
wire x_10809;
wire x_10810;
wire x_10811;
wire x_10812;
wire x_10813;
wire x_10814;
wire x_10815;
wire x_10816;
wire x_10817;
wire x_10818;
wire x_10819;
wire x_10820;
wire x_10821;
wire x_10822;
wire x_10823;
wire x_10824;
wire x_10825;
wire x_10826;
wire x_10827;
wire x_10828;
wire x_10829;
wire x_10830;
wire x_10831;
wire x_10832;
wire x_10833;
wire x_10834;
wire x_10835;
wire x_10836;
wire x_10837;
wire x_10838;
wire x_10839;
wire x_10840;
wire x_10841;
wire x_10842;
wire x_10843;
wire x_10844;
wire x_10845;
wire x_10846;
wire x_10847;
wire x_10848;
wire x_10849;
wire x_10850;
wire x_10851;
wire x_10852;
wire x_10853;
wire x_10854;
wire x_10855;
wire x_10856;
wire x_10857;
wire x_10858;
wire x_10859;
wire x_10860;
wire x_10861;
wire x_10862;
wire x_10863;
wire x_10864;
wire x_10865;
wire x_10866;
wire x_10867;
wire x_10868;
wire x_10869;
wire x_10870;
wire x_10871;
wire x_10872;
wire x_10873;
wire x_10874;
wire x_10875;
wire x_10876;
wire x_10877;
wire x_10878;
wire x_10879;
wire x_10880;
wire x_10881;
wire x_10882;
wire x_10883;
wire x_10884;
wire x_10885;
wire x_10886;
wire x_10887;
wire x_10888;
wire x_10889;
wire x_10890;
wire x_10891;
wire x_10892;
wire x_10893;
wire x_10894;
wire x_10895;
wire x_10896;
wire x_10897;
wire x_10898;
wire x_10899;
wire x_10900;
wire x_10901;
wire x_10902;
wire x_10903;
wire x_10904;
wire x_10905;
wire x_10906;
wire x_10907;
wire x_10908;
wire x_10909;
wire x_10910;
wire x_10911;
wire x_10912;
wire x_10913;
wire x_10914;
wire x_10915;
wire x_10916;
wire x_10917;
wire x_10918;
wire x_10919;
wire x_10920;
wire x_10921;
wire x_10922;
wire x_10923;
wire x_10924;
wire x_10925;
wire x_10926;
wire x_10927;
wire x_10928;
wire x_10929;
wire x_10930;
wire x_10931;
wire x_10932;
wire x_10933;
wire x_10934;
wire x_10935;
wire x_10936;
wire x_10937;
wire x_10938;
wire x_10939;
wire x_10940;
wire x_10941;
wire x_10942;
wire x_10943;
wire x_10944;
wire x_10945;
wire x_10946;
wire x_10947;
wire x_10948;
wire x_10949;
wire x_10950;
wire x_10951;
wire x_10952;
wire x_10953;
wire x_10954;
wire x_10955;
wire x_10956;
wire x_10957;
wire x_10958;
wire x_10959;
wire x_10960;
wire x_10961;
wire x_10962;
wire x_10963;
wire x_10964;
wire x_10965;
wire x_10966;
wire x_10967;
wire x_10968;
wire x_10969;
wire x_10970;
wire x_10971;
wire x_10972;
wire x_10973;
wire x_10974;
wire x_10975;
wire x_10976;
wire x_10977;
wire x_10978;
wire x_10979;
wire x_10980;
wire x_10981;
wire x_10982;
wire x_10983;
wire x_10984;
wire x_10985;
wire x_10986;
wire x_10987;
wire x_10988;
wire x_10989;
wire x_10990;
wire x_10991;
wire x_10992;
wire x_10993;
wire x_10994;
wire x_10995;
wire x_10996;
wire x_10997;
wire x_10998;
wire x_10999;
wire x_11000;
wire x_11001;
wire x_11002;
wire x_11003;
wire x_11004;
wire x_11005;
wire x_11006;
wire x_11007;
wire x_11008;
wire x_11009;
wire x_11010;
wire x_11011;
wire x_11012;
wire x_11013;
wire x_11014;
wire x_11015;
wire x_11016;
wire x_11017;
wire x_11018;
wire x_11019;
wire x_11020;
wire x_11021;
wire x_11022;
wire x_11023;
wire x_11024;
wire x_11025;
wire x_11026;
wire x_11027;
wire x_11028;
wire x_11029;
wire x_11030;
wire x_11031;
wire x_11032;
wire x_11033;
wire x_11034;
wire x_11035;
wire x_11036;
wire x_11037;
wire x_11038;
wire x_11039;
wire x_11040;
wire x_11041;
wire x_11042;
wire x_11043;
wire x_11044;
wire x_11045;
wire x_11046;
wire x_11047;
wire x_11048;
wire x_11049;
wire x_11050;
wire x_11051;
wire x_11052;
wire x_11053;
wire x_11054;
wire x_11055;
wire x_11056;
wire x_11057;
wire x_11058;
wire x_11059;
wire x_11060;
wire x_11061;
wire x_11062;
wire x_11063;
wire x_11064;
wire x_11065;
wire x_11066;
wire x_11067;
wire x_11068;
wire x_11069;
wire x_11070;
wire x_11071;
wire x_11072;
wire x_11073;
wire x_11074;
wire x_11075;
wire x_11076;
wire x_11077;
wire x_11078;
wire x_11079;
wire x_11080;
wire x_11081;
wire x_11082;
wire x_11083;
wire x_11084;
wire x_11085;
wire x_11086;
wire x_11087;
wire x_11088;
wire x_11089;
wire x_11090;
wire x_11091;
wire x_11092;
wire x_11093;
wire x_11094;
wire x_11095;
wire x_11096;
wire x_11097;
wire x_11098;
wire x_11099;
wire x_11100;
wire x_11101;
wire x_11102;
wire x_11103;
wire x_11104;
wire x_11105;
wire x_11106;
wire x_11107;
wire x_11108;
wire x_11109;
wire x_11110;
wire x_11111;
wire x_11112;
wire x_11113;
wire x_11114;
wire x_11115;
wire x_11116;
wire x_11117;
wire x_11118;
wire x_11119;
wire x_11120;
wire x_11121;
wire x_11122;
wire x_11123;
wire x_11124;
wire x_11125;
wire x_11126;
wire x_11127;
wire x_11128;
wire x_11129;
wire x_11130;
wire x_11131;
wire x_11132;
wire x_11133;
wire x_11134;
wire x_11135;
wire x_11136;
wire x_11137;
wire x_11138;
wire x_11139;
wire x_11140;
wire x_11141;
wire x_11142;
wire x_11143;
wire x_11144;
wire x_11145;
wire x_11146;
wire x_11147;
wire x_11148;
wire x_11149;
wire x_11150;
wire x_11151;
wire x_11152;
wire x_11153;
wire x_11154;
wire x_11155;
wire x_11156;
wire x_11157;
wire x_11158;
wire x_11159;
wire x_11160;
wire x_11161;
wire x_11162;
wire x_11163;
wire x_11164;
wire x_11165;
wire x_11166;
wire x_11167;
wire x_11168;
wire x_11169;
wire x_11170;
wire x_11171;
wire x_11172;
wire x_11173;
wire x_11174;
wire x_11175;
wire x_11176;
wire x_11177;
wire x_11178;
wire x_11179;
wire x_11180;
wire x_11181;
wire x_11182;
wire x_11183;
wire x_11184;
wire x_11185;
wire x_11186;
wire x_11187;
wire x_11188;
wire x_11189;
wire x_11190;
wire x_11191;
wire x_11192;
wire x_11193;
wire x_11194;
wire x_11195;
wire x_11196;
wire x_11197;
wire x_11198;
wire x_11199;
wire x_11200;
wire x_11201;
wire x_11202;
wire x_11203;
wire x_11204;
wire x_11205;
wire x_11206;
wire x_11207;
wire x_11208;
wire x_11209;
wire x_11210;
wire x_11211;
wire x_11212;
wire x_11213;
wire x_11214;
wire x_11215;
wire x_11216;
wire x_11217;
wire x_11218;
wire x_11219;
wire x_11220;
wire x_11221;
wire x_11222;
wire x_11223;
wire x_11224;
wire x_11225;
wire x_11226;
wire x_11227;
wire x_11228;
wire x_11229;
wire x_11230;
wire x_11231;
wire x_11232;
wire x_11233;
wire x_11234;
wire x_11235;
wire x_11236;
wire x_11237;
wire x_11238;
wire x_11239;
wire x_11240;
wire x_11241;
wire x_11242;
wire x_11243;
wire x_11244;
wire x_11245;
wire x_11246;
wire x_11247;
wire x_11248;
wire x_11249;
wire x_11250;
wire x_11251;
wire x_11252;
wire x_11253;
wire x_11254;
wire x_11255;
wire x_11256;
wire x_11257;
wire x_11258;
wire x_11259;
wire x_11260;
wire x_11261;
wire x_11262;
wire x_11263;
wire x_11264;
wire x_11265;
wire x_11266;
wire x_11267;
wire x_11268;
wire x_11269;
wire x_11270;
wire x_11271;
wire x_11272;
wire x_11273;
wire x_11274;
wire x_11275;
wire x_11276;
wire x_11277;
wire x_11278;
wire x_11279;
wire x_11280;
wire x_11281;
wire x_11282;
wire x_11283;
wire x_11284;
wire x_11285;
wire x_11286;
wire x_11287;
wire x_11288;
wire x_11289;
wire x_11290;
wire x_11291;
wire x_11292;
wire x_11293;
wire x_11294;
wire x_11295;
wire x_11296;
wire x_11297;
wire x_11298;
wire x_11299;
wire x_11300;
wire x_11301;
wire x_11302;
wire x_11303;
wire x_11304;
wire x_11305;
wire x_11306;
wire x_11307;
wire x_11308;
wire x_11309;
wire x_11310;
wire x_11311;
wire x_11312;
wire x_11313;
wire x_11314;
wire x_11315;
wire x_11316;
wire x_11317;
wire x_11318;
wire x_11319;
wire x_11320;
wire x_11321;
wire x_11322;
wire x_11323;
wire x_11324;
wire x_11325;
wire x_11326;
wire x_11327;
wire x_11328;
wire x_11329;
wire x_11330;
wire x_11331;
wire x_11332;
wire x_11333;
wire x_11334;
wire x_11335;
wire x_11336;
wire x_11337;
wire x_11338;
wire x_11339;
wire x_11340;
wire x_11341;
wire x_11342;
wire x_11343;
wire x_11344;
wire x_11345;
wire x_11346;
wire x_11347;
wire x_11348;
wire x_11349;
wire x_11350;
wire x_11351;
wire x_11352;
wire x_11353;
wire x_11354;
wire x_11355;
wire x_11356;
wire x_11357;
wire x_11358;
wire x_11359;
wire x_11360;
wire x_11361;
wire x_11362;
wire x_11363;
wire x_11364;
wire x_11365;
wire x_11366;
wire x_11367;
wire x_11368;
wire x_11369;
wire x_11370;
wire x_11371;
wire x_11372;
wire x_11373;
wire x_11374;
wire x_11375;
wire x_11376;
wire x_11377;
wire x_11378;
wire x_11379;
wire x_11380;
wire x_11381;
wire x_11382;
wire x_11383;
wire x_11384;
wire x_11385;
wire x_11386;
wire x_11387;
wire x_11388;
wire x_11389;
wire x_11390;
wire x_11391;
wire x_11392;
wire x_11393;
wire x_11394;
wire x_11395;
wire x_11396;
wire x_11397;
wire x_11398;
wire x_11399;
wire x_11400;
wire x_11401;
wire x_11402;
wire x_11403;
wire x_11404;
wire x_11405;
wire x_11406;
wire x_11407;
wire x_11408;
wire x_11409;
wire x_11410;
wire x_11411;
wire x_11412;
wire x_11413;
wire x_11414;
wire x_11415;
wire x_11416;
wire x_11417;
wire x_11418;
wire x_11419;
wire x_11420;
wire x_11421;
wire x_11422;
wire x_11423;
wire x_11424;
wire x_11425;
wire x_11426;
wire x_11427;
wire x_11428;
wire x_11429;
wire x_11430;
wire x_11431;
wire x_11432;
wire x_11433;
wire x_11434;
wire x_11435;
wire x_11436;
wire x_11437;
wire x_11438;
wire x_11439;
wire x_11440;
wire x_11441;
wire x_11442;
wire x_11443;
wire x_11444;
wire x_11445;
wire x_11446;
wire x_11447;
wire x_11448;
wire x_11449;
wire x_11450;
wire x_11451;
wire x_11452;
wire x_11453;
wire x_11454;
wire x_11455;
wire x_11456;
wire x_11457;
wire x_11458;
wire x_11459;
wire x_11460;
wire x_11461;
wire x_11462;
wire x_11463;
wire x_11464;
wire x_11465;
wire x_11466;
wire x_11467;
wire x_11468;
wire x_11469;
wire x_11470;
wire x_11471;
wire x_11472;
wire x_11473;
wire x_11474;
wire x_11475;
wire x_11476;
wire x_11477;
wire x_11478;
wire x_11479;
wire x_11480;
wire x_11481;
wire x_11482;
wire x_11483;
wire x_11484;
wire x_11485;
wire x_11486;
wire x_11487;
wire x_11488;
wire x_11489;
wire x_11490;
wire x_11491;
wire x_11492;
wire x_11493;
wire x_11494;
wire x_11495;
wire x_11496;
wire x_11497;
wire x_11498;
wire x_11499;
wire x_11500;
wire x_11501;
wire x_11502;
wire x_11503;
wire x_11504;
wire x_11505;
wire x_11506;
wire x_11507;
wire x_11508;
wire x_11509;
wire x_11510;
wire x_11511;
wire x_11512;
wire x_11513;
wire x_11514;
wire x_11515;
wire x_11516;
wire x_11517;
wire x_11518;
wire x_11519;
wire x_11520;
wire x_11521;
wire x_11522;
wire x_11523;
wire x_11524;
wire x_11525;
wire x_11526;
wire x_11527;
wire x_11528;
wire x_11529;
wire x_11530;
wire x_11531;
wire x_11532;
wire x_11533;
wire x_11534;
wire x_11535;
wire x_11536;
wire x_11537;
wire x_11538;
wire x_11539;
wire x_11540;
wire x_11541;
wire x_11542;
wire x_11543;
wire x_11544;
wire x_11545;
wire x_11546;
wire x_11547;
wire x_11548;
wire x_11549;
wire x_11550;
wire x_11551;
wire x_11552;
wire x_11553;
wire x_11554;
wire x_11555;
wire x_11556;
wire x_11557;
wire x_11558;
wire x_11559;
wire x_11560;
wire x_11561;
wire x_11562;
wire x_11563;
wire x_11564;
wire x_11565;
wire x_11566;
wire x_11567;
wire x_11568;
wire x_11569;
wire x_11570;
wire x_11571;
wire x_11572;
wire x_11573;
wire x_11574;
wire x_11575;
wire x_11576;
wire x_11577;
wire x_11578;
wire x_11579;
wire x_11580;
wire x_11581;
wire x_11582;
wire x_11583;
wire x_11584;
wire x_11585;
wire x_11586;
wire x_11587;
wire x_11588;
wire x_11589;
wire x_11590;
wire x_11591;
wire x_11592;
wire x_11593;
wire x_11594;
wire x_11595;
wire x_11596;
wire x_11597;
wire x_11598;
wire x_11599;
wire x_11600;
wire x_11601;
wire x_11602;
wire x_11603;
wire x_11604;
wire x_11605;
wire x_11606;
wire x_11607;
wire x_11608;
wire x_11609;
wire x_11610;
wire x_11611;
wire x_11612;
wire x_11613;
wire x_11614;
wire x_11615;
wire x_11616;
wire x_11617;
wire x_11618;
wire x_11619;
wire x_11620;
wire x_11621;
wire x_11622;
wire x_11623;
wire x_11624;
wire x_11625;
wire x_11626;
wire x_11627;
wire x_11628;
wire x_11629;
wire x_11630;
wire x_11631;
wire x_11632;
wire x_11633;
wire x_11634;
wire x_11635;
wire x_11636;
wire x_11637;
wire x_11638;
wire x_11639;
wire x_11640;
wire x_11641;
wire x_11642;
wire x_11643;
wire x_11644;
wire x_11645;
wire x_11646;
wire x_11647;
wire x_11648;
wire x_11649;
wire x_11650;
wire x_11651;
wire x_11652;
wire x_11653;
wire x_11654;
wire x_11655;
wire x_11656;
wire x_11657;
wire x_11658;
wire x_11659;
wire x_11660;
wire x_11661;
wire x_11662;
wire x_11663;
wire x_11664;
wire x_11665;
wire x_11666;
wire x_11667;
wire x_11668;
wire x_11669;
wire x_11670;
wire x_11671;
wire x_11672;
wire x_11673;
wire x_11674;
wire x_11675;
wire x_11676;
wire x_11677;
wire x_11678;
wire x_11679;
wire x_11680;
wire x_11681;
wire x_11682;
wire x_11683;
wire x_11684;
wire x_11685;
wire x_11686;
wire x_11687;
wire x_11688;
wire x_11689;
wire x_11690;
wire x_11691;
wire x_11692;
wire x_11693;
wire x_11694;
wire x_11695;
wire x_11696;
wire x_11697;
wire x_11698;
wire x_11699;
wire x_11700;
wire x_11701;
wire x_11702;
wire x_11703;
wire x_11704;
wire x_11705;
wire x_11706;
wire x_11707;
wire x_11708;
wire x_11709;
wire x_11710;
wire x_11711;
wire x_11712;
wire x_11713;
wire x_11714;
wire x_11715;
wire x_11716;
wire x_11717;
wire x_11718;
wire x_11719;
wire x_11720;
wire x_11721;
wire x_11722;
wire x_11723;
wire x_11724;
wire x_11725;
wire x_11726;
wire x_11727;
wire x_11728;
wire x_11729;
wire x_11730;
wire x_11731;
wire x_11732;
wire x_11733;
wire x_11734;
wire x_11735;
wire x_11736;
wire x_11737;
wire x_11738;
wire x_11739;
wire x_11740;
wire x_11741;
wire x_11742;
wire x_11743;
wire x_11744;
wire x_11745;
wire x_11746;
wire x_11747;
wire x_11748;
wire x_11749;
wire x_11750;
wire x_11751;
wire x_11752;
wire x_11753;
wire x_11754;
wire x_11755;
wire x_11756;
wire x_11757;
wire x_11758;
wire x_11759;
wire x_11760;
wire x_11761;
wire x_11762;
wire x_11763;
wire x_11764;
wire x_11765;
wire x_11766;
wire x_11767;
wire x_11768;
wire x_11769;
wire x_11770;
wire x_11771;
wire x_11772;
wire x_11773;
wire x_11774;
wire x_11775;
wire x_11776;
wire x_11777;
wire x_11778;
wire x_11779;
wire x_11780;
wire x_11781;
wire x_11782;
wire x_11783;
wire x_11784;
wire x_11785;
wire x_11786;
wire x_11787;
wire x_11788;
wire x_11789;
wire x_11790;
wire x_11791;
wire x_11792;
wire x_11793;
wire x_11794;
wire x_11795;
wire x_11796;
wire x_11797;
wire x_11798;
wire x_11799;
wire x_11800;
wire x_11801;
wire x_11802;
wire x_11803;
wire x_11804;
wire x_11805;
wire x_11806;
wire x_11807;
wire x_11808;
wire x_11809;
wire x_11810;
wire x_11811;
wire x_11812;
wire x_11813;
wire x_11814;
wire x_11815;
wire x_11816;
wire x_11817;
wire x_11818;
wire x_11819;
wire x_11820;
wire x_11821;
wire x_11822;
wire x_11823;
wire x_11824;
wire x_11825;
wire x_11826;
wire x_11827;
wire x_11828;
wire x_11829;
wire x_11830;
wire x_11831;
wire x_11832;
wire x_11833;
wire x_11834;
wire x_11835;
wire x_11836;
wire x_11837;
wire x_11838;
wire x_11839;
wire x_11840;
wire x_11841;
wire x_11842;
wire x_11843;
wire x_11844;
wire x_11845;
wire x_11846;
wire x_11847;
wire x_11848;
wire x_11849;
wire x_11850;
wire x_11851;
wire x_11852;
wire x_11853;
wire x_11854;
wire x_11855;
wire x_11856;
wire x_11857;
wire x_11858;
wire x_11859;
wire x_11860;
wire x_11861;
wire x_11862;
wire x_11863;
wire x_11864;
wire x_11865;
wire x_11866;
wire x_11867;
wire x_11868;
wire x_11869;
wire x_11870;
wire x_11871;
wire x_11872;
wire x_11873;
wire x_11874;
wire x_11875;
wire x_11876;
wire x_11877;
wire x_11878;
wire x_11879;
wire x_11880;
wire x_11881;
wire x_11882;
wire x_11883;
wire x_11884;
wire x_11885;
wire x_11886;
wire x_11887;
wire x_11888;
wire x_11889;
wire x_11890;
wire x_11891;
wire x_11892;
wire x_11893;
wire x_11894;
wire x_11895;
wire x_11896;
wire x_11897;
wire x_11898;
wire x_11899;
wire x_11900;
wire x_11901;
wire x_11902;
wire x_11903;
wire x_11904;
wire x_11905;
wire x_11906;
wire x_11907;
wire x_11908;
wire x_11909;
wire x_11910;
wire x_11911;
wire x_11912;
wire x_11913;
wire x_11914;
wire x_11915;
wire x_11916;
wire x_11917;
wire x_11918;
wire x_11919;
wire x_11920;
wire x_11921;
wire x_11922;
wire x_11923;
wire x_11924;
wire x_11925;
wire x_11926;
wire x_11927;
wire x_11928;
wire x_11929;
wire x_11930;
wire x_11931;
wire x_11932;
wire x_11933;
wire x_11934;
wire x_11935;
wire x_11936;
wire x_11937;
wire x_11938;
wire x_11939;
wire x_11940;
wire x_11941;
wire x_11942;
wire x_11943;
wire x_11944;
wire x_11945;
wire x_11946;
wire x_11947;
wire x_11948;
wire x_11949;
wire x_11950;
wire x_11951;
wire x_11952;
wire x_11953;
wire x_11954;
wire x_11955;
wire x_11956;
wire x_11957;
wire x_11958;
wire x_11959;
wire x_11960;
wire x_11961;
wire x_11962;
wire x_11963;
wire x_11964;
wire x_11965;
wire x_11966;
wire x_11967;
wire x_11968;
wire x_11969;
wire x_11970;
wire x_11971;
wire x_11972;
wire x_11973;
wire x_11974;
wire x_11975;
wire x_11976;
wire x_11977;
wire x_11978;
wire x_11979;
wire x_11980;
wire x_11981;
wire x_11982;
wire x_11983;
wire x_11984;
wire x_11985;
wire x_11986;
wire x_11987;
wire x_11988;
wire x_11989;
wire x_11990;
wire x_11991;
wire x_11992;
wire x_11993;
wire x_11994;
wire x_11995;
wire x_11996;
wire x_11997;
wire x_11998;
wire x_11999;
wire x_12000;
wire x_12001;
wire x_12002;
wire x_12003;
wire x_12004;
wire x_12005;
wire x_12006;
wire x_12007;
wire x_12008;
wire x_12009;
wire x_12010;
wire x_12011;
wire x_12012;
wire x_12013;
wire x_12014;
wire x_12015;
wire x_12016;
wire x_12017;
wire x_12018;
wire x_12019;
wire x_12020;
wire x_12021;
wire x_12022;
wire x_12023;
wire x_12024;
wire x_12025;
wire x_12026;
wire x_12027;
wire x_12028;
wire x_12029;
wire x_12030;
wire x_12031;
wire x_12032;
wire x_12033;
wire x_12034;
wire x_12035;
wire x_12036;
wire x_12037;
wire x_12038;
wire x_12039;
wire x_12040;
wire x_12041;
wire x_12042;
wire x_12043;
wire x_12044;
wire x_12045;
wire x_12046;
wire x_12047;
wire x_12048;
wire x_12049;
wire x_12050;
wire x_12051;
wire x_12052;
wire x_12053;
wire x_12054;
wire x_12055;
wire x_12056;
wire x_12057;
wire x_12058;
wire x_12059;
wire x_12060;
wire x_12061;
wire x_12062;
wire x_12063;
wire x_12064;
wire x_12065;
wire x_12066;
wire x_12067;
wire x_12068;
wire x_12069;
wire x_12070;
wire x_12071;
wire x_12072;
wire x_12073;
wire x_12074;
wire x_12075;
wire x_12076;
wire x_12077;
wire x_12078;
wire x_12079;
wire x_12080;
wire x_12081;
wire x_12082;
wire x_12083;
wire x_12084;
wire x_12085;
wire x_12086;
wire x_12087;
wire x_12088;
wire x_12089;
wire x_12090;
wire x_12091;
wire x_12092;
wire x_12093;
wire x_12094;
wire x_12095;
wire x_12096;
wire x_12097;
wire x_12098;
wire x_12099;
wire x_12100;
wire x_12101;
wire x_12102;
wire x_12103;
wire x_12104;
wire x_12105;
wire x_12106;
wire x_12107;
wire x_12108;
wire x_12109;
wire x_12110;
wire x_12111;
wire x_12112;
wire x_12113;
wire x_12114;
wire x_12115;
wire x_12116;
wire x_12117;
wire x_12118;
wire x_12119;
wire x_12120;
wire x_12121;
wire x_12122;
wire x_12123;
wire x_12124;
wire x_12125;
wire x_12126;
wire x_12127;
wire x_12128;
wire x_12129;
wire x_12130;
wire x_12131;
wire x_12132;
wire x_12133;
wire x_12134;
wire x_12135;
wire x_12136;
wire x_12137;
wire x_12138;
wire x_12139;
wire x_12140;
wire x_12141;
wire x_12142;
wire x_12143;
wire x_12144;
wire x_12145;
wire x_12146;
wire x_12147;
wire x_12148;
wire x_12149;
wire x_12150;
wire x_12151;
wire x_12152;
wire x_12153;
wire x_12154;
wire x_12155;
wire x_12156;
wire x_12157;
wire x_12158;
wire x_12159;
wire x_12160;
wire x_12161;
wire x_12162;
wire x_12163;
wire x_12164;
wire x_12165;
wire x_12166;
wire x_12167;
wire x_12168;
wire x_12169;
wire x_12170;
wire x_12171;
wire x_12172;
wire x_12173;
wire x_12174;
wire x_12175;
wire x_12176;
wire x_12177;
wire x_12178;
wire x_12179;
wire x_12180;
wire x_12181;
wire x_12182;
wire x_12183;
wire x_12184;
wire x_12185;
wire x_12186;
wire x_12187;
wire x_12188;
wire x_12189;
wire x_12190;
wire x_12191;
wire x_12192;
wire x_12193;
wire x_12194;
wire x_12195;
wire x_12196;
wire x_12197;
wire x_12198;
wire x_12199;
wire x_12200;
wire x_12201;
wire x_12202;
wire x_12203;
wire x_12204;
wire x_12205;
wire x_12206;
wire x_12207;
wire x_12208;
wire x_12209;
wire x_12210;
wire x_12211;
wire x_12212;
wire x_12213;
wire x_12214;
wire x_12215;
wire x_12216;
wire x_12217;
wire x_12218;
wire x_12219;
wire x_12220;
wire x_12221;
wire x_12222;
wire x_12223;
wire x_12224;
wire x_12225;
wire x_12226;
wire x_12227;
wire x_12228;
wire x_12229;
wire x_12230;
wire x_12231;
wire x_12232;
wire x_12233;
wire x_12234;
wire x_12235;
wire x_12236;
wire x_12237;
wire x_12238;
wire x_12239;
wire x_12240;
wire x_12241;
wire x_12242;
wire x_12243;
wire x_12244;
wire x_12245;
wire x_12246;
wire x_12247;
wire x_12248;
wire x_12249;
wire x_12250;
wire x_12251;
wire x_12252;
wire x_12253;
wire x_12254;
wire x_12255;
wire x_12256;
wire x_12257;
wire x_12258;
wire x_12259;
wire x_12260;
wire x_12261;
wire x_12262;
wire x_12263;
wire x_12264;
wire x_12265;
wire x_12266;
wire x_12267;
wire x_12268;
wire x_12269;
wire x_12270;
wire x_12271;
wire x_12272;
wire x_12273;
wire x_12274;
wire x_12275;
wire x_12276;
wire x_12277;
wire x_12278;
wire x_12279;
wire x_12280;
wire x_12281;
wire x_12282;
wire x_12283;
wire x_12284;
wire x_12285;
wire x_12286;
wire x_12287;
wire x_12288;
wire x_12289;
wire x_12290;
wire x_12291;
wire x_12292;
wire x_12293;
wire x_12294;
wire x_12295;
wire x_12296;
wire x_12297;
wire x_12298;
wire x_12299;
wire x_12300;
wire x_12301;
wire x_12302;
wire x_12303;
wire x_12304;
wire x_12305;
wire x_12306;
wire x_12307;
wire x_12308;
wire x_12309;
wire x_12310;
wire x_12311;
wire x_12312;
wire x_12313;
wire x_12314;
wire x_12315;
wire x_12316;
wire x_12317;
wire x_12318;
wire x_12319;
wire x_12320;
wire x_12321;
wire x_12322;
wire x_12323;
wire x_12324;
wire x_12325;
wire x_12326;
wire x_12327;
wire x_12328;
wire x_12329;
wire x_12330;
wire x_12331;
wire x_12332;
wire x_12333;
wire x_12334;
wire x_12335;
wire x_12336;
wire x_12337;
wire x_12338;
wire x_12339;
wire x_12340;
wire x_12341;
wire x_12342;
wire x_12343;
wire x_12344;
wire x_12345;
wire x_12346;
wire x_12347;
wire x_12348;
wire x_12349;
wire x_12350;
wire x_12351;
wire x_12352;
wire x_12353;
wire x_12354;
wire x_12355;
wire x_12356;
wire x_12357;
wire x_12358;
wire x_12359;
wire x_12360;
wire x_12361;
wire x_12362;
wire x_12363;
wire x_12364;
wire x_12365;
wire x_12366;
wire x_12367;
wire x_12368;
wire x_12369;
wire x_12370;
wire x_12371;
wire x_12372;
wire x_12373;
wire x_12374;
wire x_12375;
wire x_12376;
wire x_12377;
wire x_12378;
wire x_12379;
wire x_12380;
wire x_12381;
wire x_12382;
wire x_12383;
wire x_12384;
wire x_12385;
wire x_12386;
wire x_12387;
wire x_12388;
wire x_12389;
wire x_12390;
wire x_12391;
wire x_12392;
wire x_12393;
wire x_12394;
wire x_12395;
wire x_12396;
wire x_12397;
wire x_12398;
wire x_12399;
wire x_12400;
wire x_12401;
wire x_12402;
wire x_12403;
wire x_12404;
wire x_12405;
wire x_12406;
wire x_12407;
wire x_12408;
wire x_12409;
wire x_12410;
wire x_12411;
wire x_12412;
wire x_12413;
wire x_12414;
wire x_12415;
wire x_12416;
wire x_12417;
wire x_12418;
wire x_12419;
wire x_12420;
wire x_12421;
wire x_12422;
wire x_12423;
wire x_12424;
wire x_12425;
wire x_12426;
wire x_12427;
wire x_12428;
wire x_12429;
wire x_12430;
wire x_12431;
wire x_12432;
wire x_12433;
wire x_12434;
wire x_12435;
wire x_12436;
wire x_12437;
wire x_12438;
wire x_12439;
wire x_12440;
wire x_12441;
wire x_12442;
wire x_12443;
wire x_12444;
wire x_12445;
wire x_12446;
wire x_12447;
wire x_12448;
wire x_12449;
wire x_12450;
wire x_12451;
wire x_12452;
wire x_12453;
wire x_12454;
wire x_12455;
wire x_12456;
wire x_12457;
wire x_12458;
wire x_12459;
wire x_12460;
wire x_12461;
wire x_12462;
wire x_12463;
wire x_12464;
wire x_12465;
wire x_12466;
wire x_12467;
wire x_12468;
wire x_12469;
wire x_12470;
wire x_12471;
wire x_12472;
wire x_12473;
wire x_12474;
wire x_12475;
wire x_12476;
wire x_12477;
wire x_12478;
wire x_12479;
wire x_12480;
wire x_12481;
wire x_12482;
wire x_12483;
wire x_12484;
wire x_12485;
wire x_12486;
wire x_12487;
wire x_12488;
wire x_12489;
wire x_12490;
wire x_12491;
wire x_12492;
wire x_12493;
wire x_12494;
wire x_12495;
wire x_12496;
wire x_12497;
wire x_12498;
wire x_12499;
wire x_12500;
wire x_12501;
wire x_12502;
wire x_12503;
wire x_12504;
wire x_12505;
wire x_12506;
wire x_12507;
wire x_12508;
wire x_12509;
wire x_12510;
wire x_12511;
wire x_12512;
wire x_12513;
wire x_12514;
wire x_12515;
wire x_12516;
wire x_12517;
wire x_12518;
wire x_12519;
wire x_12520;
wire x_12521;
wire x_12522;
wire x_12523;
wire x_12524;
wire x_12525;
wire x_12526;
wire x_12527;
wire x_12528;
wire x_12529;
wire x_12530;
wire x_12531;
wire x_12532;
wire x_12533;
wire x_12534;
wire x_12535;
wire x_12536;
wire x_12537;
wire x_12538;
wire x_12539;
wire x_12540;
wire x_12541;
wire x_12542;
wire x_12543;
wire x_12544;
wire x_12545;
wire x_12546;
wire x_12547;
wire x_12548;
wire x_12549;
wire x_12550;
wire x_12551;
wire x_12552;
wire x_12553;
wire x_12554;
wire x_12555;
wire x_12556;
wire x_12557;
wire x_12558;
wire x_12559;
wire x_12560;
wire x_12561;
wire x_12562;
wire x_12563;
wire x_12564;
wire x_12565;
wire x_12566;
wire x_12567;
wire x_12568;
wire x_12569;
wire x_12570;
wire x_12571;
wire x_12572;
wire x_12573;
wire x_12574;
wire x_12575;
wire x_12576;
wire x_12577;
wire x_12578;
wire x_12579;
wire x_12580;
wire x_12581;
wire x_12582;
wire x_12583;
wire x_12584;
wire x_12585;
wire x_12586;
wire x_12587;
wire x_12588;
wire x_12589;
wire x_12590;
wire x_12591;
wire x_12592;
wire x_12593;
wire x_12594;
wire x_12595;
wire x_12596;
wire x_12597;
wire x_12598;
wire x_12599;
wire x_12600;
wire x_12601;
wire x_12602;
wire x_12603;
wire x_12604;
wire x_12605;
wire x_12606;
wire x_12607;
wire x_12608;
wire x_12609;
wire x_12610;
wire x_12611;
wire x_12612;
wire x_12613;
wire x_12614;
wire x_12615;
wire x_12616;
wire x_12617;
wire x_12618;
wire x_12619;
wire x_12620;
wire x_12621;
wire x_12622;
wire x_12623;
wire x_12624;
wire x_12625;
wire x_12626;
wire x_12627;
wire x_12628;
wire x_12629;
wire x_12630;
wire x_12631;
wire x_12632;
wire x_12633;
wire x_12634;
wire x_12635;
wire x_12636;
wire x_12637;
wire x_12638;
wire x_12639;
wire x_12640;
wire x_12641;
wire x_12642;
wire x_12643;
wire x_12644;
wire x_12645;
wire x_12646;
wire x_12647;
wire x_12648;
wire x_12649;
wire x_12650;
wire x_12651;
wire x_12652;
wire x_12653;
wire x_12654;
wire x_12655;
wire x_12656;
wire x_12657;
wire x_12658;
wire x_12659;
wire x_12660;
wire x_12661;
wire x_12662;
wire x_12663;
wire x_12664;
wire x_12665;
wire x_12666;
wire x_12667;
wire x_12668;
wire x_12669;
wire x_12670;
wire x_12671;
wire x_12672;
wire x_12673;
wire x_12674;
wire x_12675;
wire x_12676;
wire x_12677;
wire x_12678;
wire x_12679;
wire x_12680;
wire x_12681;
wire x_12682;
wire x_12683;
wire x_12684;
wire x_12685;
wire x_12686;
wire x_12687;
wire x_12688;
wire x_12689;
wire x_12690;
wire x_12691;
wire x_12692;
wire x_12693;
wire x_12694;
wire x_12695;
wire x_12696;
wire x_12697;
wire x_12698;
wire x_12699;
wire x_12700;
wire x_12701;
wire x_12702;
wire x_12703;
wire x_12704;
wire x_12705;
wire x_12706;
wire x_12707;
wire x_12708;
wire x_12709;
wire x_12710;
wire x_12711;
wire x_12712;
wire x_12713;
wire x_12714;
wire x_12715;
wire x_12716;
wire x_12717;
wire x_12718;
wire x_12719;
wire x_12720;
wire x_12721;
wire x_12722;
wire x_12723;
wire x_12724;
wire x_12725;
wire x_12726;
wire x_12727;
wire x_12728;
wire x_12729;
wire x_12730;
wire x_12731;
wire x_12732;
wire x_12733;
wire x_12734;
wire x_12735;
wire x_12736;
wire x_12737;
wire x_12738;
wire x_12739;
wire x_12740;
wire x_12741;
wire x_12742;
wire x_12743;
wire x_12744;
wire x_12745;
wire x_12746;
wire x_12747;
wire x_12748;
wire x_12749;
wire x_12750;
wire x_12751;
wire x_12752;
wire x_12753;
wire x_12754;
wire x_12755;
wire x_12756;
wire x_12757;
wire x_12758;
wire x_12759;
wire x_12760;
wire x_12761;
wire x_12762;
wire x_12763;
wire x_12764;
wire x_12765;
wire x_12766;
wire x_12767;
wire x_12768;
wire x_12769;
wire x_12770;
wire x_12771;
wire x_12772;
wire x_12773;
wire x_12774;
wire x_12775;
wire x_12776;
wire x_12777;
wire x_12778;
wire x_12779;
wire x_12780;
wire x_12781;
wire x_12782;
wire x_12783;
wire x_12784;
wire x_12785;
wire x_12786;
wire x_12787;
wire x_12788;
wire x_12789;
wire x_12790;
wire x_12791;
wire x_12792;
wire x_12793;
wire x_12794;
wire x_12795;
wire x_12796;
wire x_12797;
wire x_12798;
wire x_12799;
wire x_12800;
wire x_12801;
wire x_12802;
wire x_12803;
wire x_12804;
wire x_12805;
wire x_12806;
wire x_12807;
wire x_12808;
wire x_12809;
wire x_12810;
wire x_12811;
wire x_12812;
wire x_12813;
wire x_12814;
wire x_12815;
wire x_12816;
wire x_12817;
wire x_12818;
wire x_12819;
wire x_12820;
wire x_12821;
wire x_12822;
wire x_12823;
wire x_12824;
wire x_12825;
wire x_12826;
wire x_12827;
wire x_12828;
wire x_12829;
wire x_12830;
wire x_12831;
wire x_12832;
wire x_12833;
wire x_12834;
wire x_12835;
wire x_12836;
wire x_12837;
wire x_12838;
wire x_12839;
wire x_12840;
wire x_12841;
wire x_12842;
wire x_12843;
wire x_12844;
wire x_12845;
wire x_12846;
wire x_12847;
wire x_12848;
wire x_12849;
wire x_12850;
wire x_12851;
wire x_12852;
wire x_12853;
wire x_12854;
wire x_12855;
wire x_12856;
wire x_12857;
wire x_12858;
wire x_12859;
wire x_12860;
wire x_12861;
wire x_12862;
wire x_12863;
wire x_12864;
wire x_12865;
wire x_12866;
wire x_12867;
wire x_12868;
wire x_12869;
wire x_12870;
wire x_12871;
wire x_12872;
wire x_12873;
wire x_12874;
wire x_12875;
wire x_12876;
wire x_12877;
wire x_12878;
wire x_12879;
wire x_12880;
wire x_12881;
wire x_12882;
wire x_12883;
wire x_12884;
wire x_12885;
wire x_12886;
wire x_12887;
wire x_12888;
wire x_12889;
wire x_12890;
wire x_12891;
wire x_12892;
wire x_12893;
wire x_12894;
wire x_12895;
wire x_12896;
wire x_12897;
wire x_12898;
wire x_12899;
wire x_12900;
wire x_12901;
wire x_12902;
wire x_12903;
wire x_12904;
wire x_12905;
wire x_12906;
wire x_12907;
wire x_12908;
wire x_12909;
wire x_12910;
wire x_12911;
wire x_12912;
wire x_12913;
wire x_12914;
wire x_12915;
wire x_12916;
wire x_12917;
wire x_12918;
wire x_12919;
wire x_12920;
wire x_12921;
wire x_12922;
wire x_12923;
wire x_12924;
wire x_12925;
wire x_12926;
wire x_12927;
wire x_12928;
wire x_12929;
wire x_12930;
wire x_12931;
wire x_12932;
wire x_12933;
wire x_12934;
wire x_12935;
wire x_12936;
wire x_12937;
wire x_12938;
wire x_12939;
wire x_12940;
wire x_12941;
wire x_12942;
wire x_12943;
wire x_12944;
wire x_12945;
wire x_12946;
wire x_12947;
wire x_12948;
wire x_12949;
wire x_12950;
wire x_12951;
wire x_12952;
wire x_12953;
wire x_12954;
wire x_12955;
wire x_12956;
wire x_12957;
wire x_12958;
wire x_12959;
wire x_12960;
wire x_12961;
wire x_12962;
wire x_12963;
wire x_12964;
wire x_12965;
wire x_12966;
wire x_12967;
wire x_12968;
wire x_12969;
wire x_12970;
wire x_12971;
wire x_12972;
wire x_12973;
wire x_12974;
wire x_12975;
wire x_12976;
wire x_12977;
wire x_12978;
wire x_12979;
wire x_12980;
wire x_12981;
wire x_12982;
wire x_12983;
wire x_12984;
wire x_12985;
wire x_12986;
wire x_12987;
wire x_12988;
wire x_12989;
wire x_12990;
wire x_12991;
wire x_12992;
wire x_12993;
wire x_12994;
wire x_12995;
wire x_12996;
wire x_12997;
wire x_12998;
wire x_12999;
wire x_13000;
wire x_13001;
wire x_13002;
wire x_13003;
wire x_13004;
wire x_13005;
wire x_13006;
wire x_13007;
wire x_13008;
wire x_13009;
wire x_13010;
wire x_13011;
wire x_13012;
wire x_13013;
wire x_13014;
wire x_13015;
wire x_13016;
wire x_13017;
wire x_13018;
wire x_13019;
wire x_13020;
wire x_13021;
wire x_13022;
wire x_13023;
wire x_13024;
wire x_13025;
wire x_13026;
wire x_13027;
wire x_13028;
wire x_13029;
wire x_13030;
wire x_13031;
wire x_13032;
wire x_13033;
wire x_13034;
wire x_13035;
wire x_13036;
wire x_13037;
wire x_13038;
wire x_13039;
wire x_13040;
wire x_13041;
wire x_13042;
wire x_13043;
wire x_13044;
wire x_13045;
wire x_13046;
wire x_13047;
wire x_13048;
wire x_13049;
wire x_13050;
wire x_13051;
wire x_13052;
wire x_13053;
wire x_13054;
wire x_13055;
wire x_13056;
wire x_13057;
wire x_13058;
wire x_13059;
wire x_13060;
wire x_13061;
wire x_13062;
wire x_13063;
wire x_13064;
wire x_13065;
wire x_13066;
wire x_13067;
wire x_13068;
wire x_13069;
wire x_13070;
wire x_13071;
wire x_13072;
wire x_13073;
wire x_13074;
wire x_13075;
wire x_13076;
wire x_13077;
wire x_13078;
wire x_13079;
wire x_13080;
wire x_13081;
wire x_13082;
wire x_13083;
wire x_13084;
wire x_13085;
wire x_13086;
wire x_13087;
wire x_13088;
wire x_13089;
wire x_13090;
wire x_13091;
wire x_13092;
wire x_13093;
wire x_13094;
wire x_13095;
wire x_13096;
wire x_13097;
wire x_13098;
wire x_13099;
wire x_13100;
wire x_13101;
wire x_13102;
wire x_13103;
wire x_13104;
wire x_13105;
wire x_13106;
wire x_13107;
wire x_13108;
wire x_13109;
wire x_13110;
wire x_13111;
wire x_13112;
wire x_13113;
wire x_13114;
wire x_13115;
wire x_13116;
wire x_13117;
wire x_13118;
wire x_13119;
wire x_13120;
wire x_13121;
wire x_13122;
wire x_13123;
wire x_13124;
wire x_13125;
wire x_13126;
wire x_13127;
wire x_13128;
wire x_13129;
wire x_13130;
wire x_13131;
wire x_13132;
wire x_13133;
wire x_13134;
wire x_13135;
wire x_13136;
wire x_13137;
wire x_13138;
wire x_13139;
wire x_13140;
wire x_13141;
wire x_13142;
wire x_13143;
wire x_13144;
wire x_13145;
wire x_13146;
wire x_13147;
wire x_13148;
wire x_13149;
wire x_13150;
wire x_13151;
wire x_13152;
wire x_13153;
wire x_13154;
wire x_13155;
wire x_13156;
wire x_13157;
wire x_13158;
wire x_13159;
wire x_13160;
wire x_13161;
wire x_13162;
wire x_13163;
wire x_13164;
wire x_13165;
wire x_13166;
wire x_13167;
wire x_13168;
wire x_13169;
wire x_13170;
wire x_13171;
wire x_13172;
wire x_13173;
wire x_13174;
wire x_13175;
wire x_13176;
wire x_13177;
wire x_13178;
wire x_13179;
wire x_13180;
wire x_13181;
wire x_13182;
wire x_13183;
wire x_13184;
wire x_13185;
wire x_13186;
wire x_13187;
wire x_13188;
wire x_13189;
wire x_13190;
wire x_13191;
wire x_13192;
wire x_13193;
wire x_13194;
wire x_13195;
wire x_13196;
wire x_13197;
wire x_13198;
wire x_13199;
wire x_13200;
wire x_13201;
wire x_13202;
wire x_13203;
wire x_13204;
wire x_13205;
wire x_13206;
wire x_13207;
wire x_13208;
wire x_13209;
wire x_13210;
wire x_13211;
wire x_13212;
wire x_13213;
wire x_13214;
wire x_13215;
wire x_13216;
wire x_13217;
wire x_13218;
wire x_13219;
wire x_13220;
wire x_13221;
wire x_13222;
wire x_13223;
wire x_13224;
wire x_13225;
wire x_13226;
wire x_13227;
wire x_13228;
wire x_13229;
wire x_13230;
wire x_13231;
wire x_13232;
wire x_13233;
wire x_13234;
wire x_13235;
wire x_13236;
wire x_13237;
wire x_13238;
wire x_13239;
wire x_13240;
wire x_13241;
wire x_13242;
wire x_13243;
wire x_13244;
wire x_13245;
wire x_13246;
wire x_13247;
wire x_13248;
wire x_13249;
wire x_13250;
wire x_13251;
wire x_13252;
wire x_13253;
wire x_13254;
wire x_13255;
wire x_13256;
wire x_13257;
wire x_13258;
wire x_13259;
wire x_13260;
wire x_13261;
wire x_13262;
wire x_13263;
wire x_13264;
wire x_13265;
wire x_13266;
wire x_13267;
wire x_13268;
wire x_13269;
wire x_13270;
wire x_13271;
wire x_13272;
wire x_13273;
wire x_13274;
wire x_13275;
wire x_13276;
wire x_13277;
wire x_13278;
wire x_13279;
wire x_13280;
wire x_13281;
wire x_13282;
wire x_13283;
wire x_13284;
wire x_13285;
wire x_13286;
wire x_13287;
wire x_13288;
wire x_13289;
wire x_13290;
wire x_13291;
wire x_13292;
wire x_13293;
wire x_13294;
wire x_13295;
wire x_13296;
wire x_13297;
wire x_13298;
wire x_13299;
wire x_13300;
wire x_13301;
wire x_13302;
wire x_13303;
wire x_13304;
wire x_13305;
wire x_13306;
wire x_13307;
wire x_13308;
wire x_13309;
wire x_13310;
wire x_13311;
wire x_13312;
wire x_13313;
wire x_13314;
wire x_13315;
wire x_13316;
wire x_13317;
wire x_13318;
wire x_13319;
wire x_13320;
wire x_13321;
wire x_13322;
wire x_13323;
wire x_13324;
wire x_13325;
wire x_13326;
wire x_13327;
wire x_13328;
wire x_13329;
wire x_13330;
wire x_13331;
wire x_13332;
wire x_13333;
wire x_13334;
wire x_13335;
wire x_13336;
wire x_13337;
wire x_13338;
wire x_13339;
wire x_13340;
wire x_13341;
wire x_13342;
wire x_13343;
wire x_13344;
wire x_13345;
wire x_13346;
wire x_13347;
wire x_13348;
wire x_13349;
wire x_13350;
wire x_13351;
wire x_13352;
wire x_13353;
wire x_13354;
wire x_13355;
wire x_13356;
wire x_13357;
wire x_13358;
wire x_13359;
wire x_13360;
wire x_13361;
wire x_13362;
wire x_13363;
wire x_13364;
wire x_13365;
wire x_13366;
wire x_13367;
wire x_13368;
wire x_13369;
wire x_13370;
wire x_13371;
wire x_13372;
wire x_13373;
wire x_13374;
wire x_13375;
wire x_13376;
wire x_13377;
wire x_13378;
wire x_13379;
wire x_13380;
wire x_13381;
wire x_13382;
wire x_13383;
wire x_13384;
wire x_13385;
wire x_13386;
wire x_13387;
wire x_13388;
wire x_13389;
wire x_13390;
wire x_13391;
wire x_13392;
wire x_13393;
wire x_13394;
wire x_13395;
wire x_13396;
wire x_13397;
wire x_13398;
wire x_13399;
wire x_13400;
wire x_13401;
wire x_13402;
wire x_13403;
wire x_13404;
wire x_13405;
wire x_13406;
wire x_13407;
wire x_13408;
wire x_13409;
wire x_13410;
wire x_13411;
wire x_13412;
wire x_13413;
wire x_13414;
wire x_13415;
wire x_13416;
wire x_13417;
wire x_13418;
wire x_13419;
wire x_13420;
wire x_13421;
wire x_13422;
wire x_13423;
wire x_13424;
wire x_13425;
wire x_13426;
wire x_13427;
wire x_13428;
wire x_13429;
wire x_13430;
wire x_13431;
wire x_13432;
wire x_13433;
wire x_13434;
wire x_13435;
wire x_13436;
wire x_13437;
wire x_13438;
wire x_13439;
wire x_13440;
wire x_13441;
wire x_13442;
wire x_13443;
wire x_13444;
wire x_13445;
wire x_13446;
wire x_13447;
wire x_13448;
wire x_13449;
wire x_13450;
wire x_13451;
wire x_13452;
wire x_13453;
wire x_13454;
wire x_13455;
wire x_13456;
wire x_13457;
wire x_13458;
wire x_13459;
wire x_13460;
wire x_13461;
wire x_13462;
wire x_13463;
wire x_13464;
wire x_13465;
wire x_13466;
wire x_13467;
wire x_13468;
wire x_13469;
wire x_13470;
wire x_13471;
wire x_13472;
wire x_13473;
wire x_13474;
wire x_13475;
wire x_13476;
wire x_13477;
wire x_13478;
wire x_13479;
wire x_13480;
wire x_13481;
wire x_13482;
wire x_13483;
wire x_13484;
wire x_13485;
wire x_13486;
wire x_13487;
wire x_13488;
wire x_13489;
wire x_13490;
wire x_13491;
wire x_13492;
wire x_13493;
wire x_13494;
wire x_13495;
wire x_13496;
wire x_13497;
wire x_13498;
wire x_13499;
wire x_13500;
wire x_13501;
wire x_13502;
wire x_13503;
wire x_13504;
wire x_13505;
wire x_13506;
wire x_13507;
wire x_13508;
wire x_13509;
wire x_13510;
wire x_13511;
wire x_13512;
wire x_13513;
wire x_13514;
wire x_13515;
wire x_13516;
wire x_13517;
wire x_13518;
wire x_13519;
wire x_13520;
wire x_13521;
wire x_13522;
wire x_13523;
wire x_13524;
wire x_13525;
wire x_13526;
wire x_13527;
wire x_13528;
wire x_13529;
wire x_13530;
wire x_13531;
wire x_13532;
wire x_13533;
wire x_13534;
wire x_13535;
wire x_13536;
wire x_13537;
wire x_13538;
wire x_13539;
wire x_13540;
wire x_13541;
wire x_13542;
wire x_13543;
wire x_13544;
wire x_13545;
wire x_13546;
wire x_13547;
wire x_13548;
wire x_13549;
wire x_13550;
wire x_13551;
wire x_13552;
wire x_13553;
wire x_13554;
wire x_13555;
wire x_13556;
wire x_13557;
wire x_13558;
wire x_13559;
wire x_13560;
wire x_13561;
wire x_13562;
wire x_13563;
wire x_13564;
wire x_13565;
wire x_13566;
wire x_13567;
wire x_13568;
wire x_13569;
wire x_13570;
wire x_13571;
wire x_13572;
wire x_13573;
wire x_13574;
wire x_13575;
wire x_13576;
wire x_13577;
wire x_13578;
wire x_13579;
wire x_13580;
wire x_13581;
wire x_13582;
wire x_13583;
wire x_13584;
wire x_13585;
wire x_13586;
wire x_13587;
wire x_13588;
wire x_13589;
wire x_13590;
wire x_13591;
wire x_13592;
wire x_13593;
wire x_13594;
wire x_13595;
wire x_13596;
wire x_13597;
wire x_13598;
wire x_13599;
wire x_13600;
wire x_13601;
wire x_13602;
wire x_13603;
wire x_13604;
wire x_13605;
wire x_13606;
wire x_13607;
wire x_13608;
wire x_13609;
wire x_13610;
wire x_13611;
wire x_13612;
wire x_13613;
wire x_13614;
wire x_13615;
wire x_13616;
wire x_13617;
wire x_13618;
wire x_13619;
wire x_13620;
wire x_13621;
wire x_13622;
wire x_13623;
wire x_13624;
wire x_13625;
wire x_13626;
wire x_13627;
wire x_13628;
wire x_13629;
wire x_13630;
wire x_13631;
wire x_13632;
wire x_13633;
wire x_13634;
wire x_13635;
wire x_13636;
wire x_13637;
wire x_13638;
wire x_13639;
wire x_13640;
wire x_13641;
wire x_13642;
wire x_13643;
wire x_13644;
wire x_13645;
wire x_13646;
wire x_13647;
wire x_13648;
wire x_13649;
wire x_13650;
wire x_13651;
wire x_13652;
wire x_13653;
wire x_13654;
wire x_13655;
wire x_13656;
wire x_13657;
wire x_13658;
wire x_13659;
wire x_13660;
wire x_13661;
wire x_13662;
wire x_13663;
wire x_13664;
wire x_13665;
wire x_13666;
wire x_13667;
wire x_13668;
wire x_13669;
wire x_13670;
wire x_13671;
wire x_13672;
wire x_13673;
wire x_13674;
wire x_13675;
wire x_13676;
wire x_13677;
wire x_13678;
wire x_13679;
wire x_13680;
wire x_13681;
wire x_13682;
wire x_13683;
wire x_13684;
wire x_13685;
wire x_13686;
wire x_13687;
wire x_13688;
wire x_13689;
wire x_13690;
wire x_13691;
wire x_13692;
wire x_13693;
wire x_13694;
wire x_13695;
wire x_13696;
wire x_13697;
wire x_13698;
wire x_13699;
wire x_13700;
wire x_13701;
wire x_13702;
wire x_13703;
wire x_13704;
wire x_13705;
wire x_13706;
wire x_13707;
wire x_13708;
wire x_13709;
wire x_13710;
wire x_13711;
wire x_13712;
wire x_13713;
wire x_13714;
wire x_13715;
wire x_13716;
wire x_13717;
wire x_13718;
wire x_13719;
wire x_13720;
wire x_13721;
wire x_13722;
wire x_13723;
wire x_13724;
wire x_13725;
wire x_13726;
wire x_13727;
wire x_13728;
wire x_13729;
wire x_13730;
wire x_13731;
wire x_13732;
wire x_13733;
wire x_13734;
wire x_13735;
wire x_13736;
wire x_13737;
wire x_13738;
wire x_13739;
wire x_13740;
wire x_13741;
wire x_13742;
wire x_13743;
wire x_13744;
wire x_13745;
wire x_13746;
wire x_13747;
wire x_13748;
wire x_13749;
wire x_13750;
wire x_13751;
wire x_13752;
wire x_13753;
wire x_13754;
wire x_13755;
wire x_13756;
wire x_13757;
wire x_13758;
wire x_13759;
wire x_13760;
wire x_13761;
wire x_13762;
wire x_13763;
wire x_13764;
wire x_13765;
wire x_13766;
wire x_13767;
wire x_13768;
wire x_13769;
wire x_13770;
wire x_13771;
wire x_13772;
wire x_13773;
wire x_13774;
wire x_13775;
wire x_13776;
wire x_13777;
wire x_13778;
wire x_13779;
wire x_13780;
wire x_13781;
wire x_13782;
wire x_13783;
wire x_13784;
wire x_13785;
wire x_13786;
wire x_13787;
wire x_13788;
wire x_13789;
wire x_13790;
wire x_13791;
wire x_13792;
wire x_13793;
wire x_13794;
wire x_13795;
wire x_13796;
wire x_13797;
wire x_13798;
wire x_13799;
wire x_13800;
wire x_13801;
wire x_13802;
wire x_13803;
wire x_13804;
wire x_13805;
wire x_13806;
wire x_13807;
wire x_13808;
wire x_13809;
wire x_13810;
wire x_13811;
wire x_13812;
wire x_13813;
wire x_13814;
wire x_13815;
wire x_13816;
wire x_13817;
wire x_13818;
wire x_13819;
wire x_13820;
wire x_13821;
wire x_13822;
wire x_13823;
wire x_13824;
wire x_13825;
wire x_13826;
wire x_13827;
wire x_13828;
wire x_13829;
wire x_13830;
wire x_13831;
wire x_13832;
wire x_13833;
wire x_13834;
wire x_13835;
wire x_13836;
wire x_13837;
wire x_13838;
wire x_13839;
wire x_13840;
wire x_13841;
wire x_13842;
wire x_13843;
wire x_13844;
wire x_13845;
wire x_13846;
wire x_13847;
wire x_13848;
wire x_13849;
wire x_13850;
wire x_13851;
wire x_13852;
wire x_13853;
wire x_13854;
wire x_13855;
wire x_13856;
wire x_13857;
wire x_13858;
wire x_13859;
wire x_13860;
wire x_13861;
wire x_13862;
wire x_13863;
wire x_13864;
wire x_13865;
wire x_13866;
wire x_13867;
wire x_13868;
wire x_13869;
wire x_13870;
wire x_13871;
wire x_13872;
wire x_13873;
wire x_13874;
wire x_13875;
wire x_13876;
wire x_13877;
wire x_13878;
wire x_13879;
wire x_13880;
wire x_13881;
wire x_13882;
wire x_13883;
wire x_13884;
wire x_13885;
wire x_13886;
wire x_13887;
wire x_13888;
wire x_13889;
wire x_13890;
wire x_13891;
wire x_13892;
wire x_13893;
wire x_13894;
wire x_13895;
wire x_13896;
wire x_13897;
wire x_13898;
wire x_13899;
wire x_13900;
wire x_13901;
wire x_13902;
wire x_13903;
wire x_13904;
wire x_13905;
wire x_13906;
wire x_13907;
wire x_13908;
wire x_13909;
wire x_13910;
wire x_13911;
wire x_13912;
wire x_13913;
wire x_13914;
wire x_13915;
wire x_13916;
wire x_13917;
wire x_13918;
wire x_13919;
wire x_13920;
wire x_13921;
wire x_13922;
wire x_13923;
wire x_13924;
wire x_13925;
wire x_13926;
wire x_13927;
wire x_13928;
wire x_13929;
wire x_13930;
wire x_13931;
wire x_13932;
wire x_13933;
wire x_13934;
wire x_13935;
wire x_13936;
wire x_13937;
wire x_13938;
wire x_13939;
wire x_13940;
wire x_13941;
wire x_13942;
wire x_13943;
wire x_13944;
wire x_13945;
wire x_13946;
wire x_13947;
wire x_13948;
wire x_13949;
wire x_13950;
wire x_13951;
wire x_13952;
wire x_13953;
wire x_13954;
wire x_13955;
wire x_13956;
wire x_13957;
wire x_13958;
wire x_13959;
wire x_13960;
wire x_13961;
wire x_13962;
wire x_13963;
wire x_13964;
wire x_13965;
wire x_13966;
wire x_13967;
wire x_13968;
wire x_13969;
wire x_13970;
wire x_13971;
wire x_13972;
wire x_13973;
wire x_13974;
wire x_13975;
wire x_13976;
wire x_13977;
wire x_13978;
wire x_13979;
wire x_13980;
wire x_13981;
wire x_13982;
wire x_13983;
wire x_13984;
wire x_13985;
wire x_13986;
wire x_13987;
wire x_13988;
wire x_13989;
wire x_13990;
wire x_13991;
wire x_13992;
wire x_13993;
wire x_13994;
wire x_13995;
wire x_13996;
wire x_13997;
wire x_13998;
wire x_13999;
wire x_14000;
wire x_14001;
wire x_14002;
wire x_14003;
wire x_14004;
wire x_14005;
wire x_14006;
wire x_14007;
wire x_14008;
wire x_14009;
wire x_14010;
wire x_14011;
wire x_14012;
wire x_14013;
wire x_14014;
wire x_14015;
wire x_14016;
wire x_14017;
wire x_14018;
wire x_14019;
wire x_14020;
wire x_14021;
wire x_14022;
wire x_14023;
wire x_14024;
wire x_14025;
wire x_14026;
wire x_14027;
wire x_14028;
wire x_14029;
wire x_14030;
wire x_14031;
wire x_14032;
wire x_14033;
wire x_14034;
wire x_14035;
wire x_14036;
wire x_14037;
wire x_14038;
wire x_14039;
wire x_14040;
wire x_14041;
wire x_14042;
wire x_14043;
wire x_14044;
wire x_14045;
wire x_14046;
wire x_14047;
wire x_14048;
wire x_14049;
wire x_14050;
wire x_14051;
wire x_14052;
wire x_14053;
wire x_14054;
wire x_14055;
wire x_14056;
wire x_14057;
wire x_14058;
wire x_14059;
wire x_14060;
wire x_14061;
wire x_14062;
wire x_14063;
wire x_14064;
wire x_14065;
wire x_14066;
wire x_14067;
wire x_14068;
wire x_14069;
wire x_14070;
wire x_14071;
wire x_14072;
wire x_14073;
wire x_14074;
wire x_14075;
wire x_14076;
wire x_14077;
wire x_14078;
wire x_14079;
wire x_14080;
wire x_14081;
wire x_14082;
wire x_14083;
wire x_14084;
wire x_14085;
wire x_14086;
wire x_14087;
wire x_14088;
wire x_14089;
wire x_14090;
wire x_14091;
wire x_14092;
wire x_14093;
wire x_14094;
wire x_14095;
wire x_14096;
wire x_14097;
wire x_14098;
wire x_14099;
wire x_14100;
wire x_14101;
wire x_14102;
wire x_14103;
wire x_14104;
wire x_14105;
wire x_14106;
wire x_14107;
wire x_14108;
wire x_14109;
wire x_14110;
wire x_14111;
wire x_14112;
wire x_14113;
wire x_14114;
wire x_14115;
wire x_14116;
wire x_14117;
wire x_14118;
wire x_14119;
wire x_14120;
wire x_14121;
wire x_14122;
wire x_14123;
wire x_14124;
wire x_14125;
wire x_14126;
wire x_14127;
wire x_14128;
wire x_14129;
wire x_14130;
wire x_14131;
wire x_14132;
wire x_14133;
wire x_14134;
wire x_14135;
wire x_14136;
wire x_14137;
wire x_14138;
wire x_14139;
wire x_14140;
wire x_14141;
wire x_14142;
wire x_14143;
wire x_14144;
wire x_14145;
wire x_14146;
wire x_14147;
wire x_14148;
wire x_14149;
wire x_14150;
wire x_14151;
wire x_14152;
wire x_14153;
wire x_14154;
wire x_14155;
wire x_14156;
wire x_14157;
wire x_14158;
wire x_14159;
wire x_14160;
wire x_14161;
wire x_14162;
wire x_14163;
wire x_14164;
wire x_14165;
wire x_14166;
wire x_14167;
wire x_14168;
wire x_14169;
wire x_14170;
wire x_14171;
wire x_14172;
wire x_14173;
wire x_14174;
wire x_14175;
wire x_14176;
wire x_14177;
wire x_14178;
wire x_14179;
wire x_14180;
wire x_14181;
wire x_14182;
wire x_14183;
wire x_14184;
wire x_14185;
wire x_14186;
wire x_14187;
wire x_14188;
wire x_14189;
wire x_14190;
wire x_14191;
wire x_14192;
wire x_14193;
wire x_14194;
wire x_14195;
wire x_14196;
wire x_14197;
wire x_14198;
wire x_14199;
wire x_14200;
wire x_14201;
wire x_14202;
wire x_14203;
wire x_14204;
wire x_14205;
wire x_14206;
wire x_14207;
wire x_14208;
wire x_14209;
wire x_14210;
wire x_14211;
wire x_14212;
wire x_14213;
wire x_14214;
wire x_14215;
wire x_14216;
wire x_14217;
wire x_14218;
wire x_14219;
wire x_14220;
wire x_14221;
wire x_14222;
wire x_14223;
wire x_14224;
wire x_14225;
wire x_14226;
wire x_14227;
wire x_14228;
wire x_14229;
wire x_14230;
wire x_14231;
wire x_14232;
wire x_14233;
wire x_14234;
wire x_14235;
wire x_14236;
wire x_14237;
wire x_14238;
wire x_14239;
wire x_14240;
wire x_14241;
wire x_14242;
wire x_14243;
wire x_14244;
wire x_14245;
wire x_14246;
wire x_14247;
wire x_14248;
wire x_14249;
wire x_14250;
wire x_14251;
wire x_14252;
wire x_14253;
wire x_14254;
wire x_14255;
wire x_14256;
wire x_14257;
wire x_14258;
wire x_14259;
wire x_14260;
wire x_14261;
wire x_14262;
wire x_14263;
wire x_14264;
wire x_14265;
wire x_14266;
wire x_14267;
wire x_14268;
wire x_14269;
wire x_14270;
wire x_14271;
wire x_14272;
wire x_14273;
wire x_14274;
wire x_14275;
wire x_14276;
wire x_14277;
wire x_14278;
wire x_14279;
wire x_14280;
wire x_14281;
wire x_14282;
wire x_14283;
wire x_14284;
wire x_14285;
wire x_14286;
wire x_14287;
wire x_14288;
wire x_14289;
wire x_14290;
wire x_14291;
wire x_14292;
wire x_14293;
wire x_14294;
wire x_14295;
wire x_14296;
wire x_14297;
wire x_14298;
wire x_14299;
wire x_14300;
wire x_14301;
wire x_14302;
wire x_14303;
wire x_14304;
wire x_14305;
wire x_14306;
wire x_14307;
wire x_14308;
wire x_14309;
wire x_14310;
wire x_14311;
wire x_14312;
wire x_14313;
wire x_14314;
wire x_14315;
wire x_14316;
wire x_14317;
wire x_14318;
wire x_14319;
wire x_14320;
wire x_14321;
wire x_14322;
wire x_14323;
wire x_14324;
wire x_14325;
wire x_14326;
wire x_14327;
wire x_14328;
wire x_14329;
wire x_14330;
wire x_14331;
wire x_14332;
wire x_14333;
wire x_14334;
wire x_14335;
wire x_14336;
wire x_14337;
wire x_14338;
wire x_14339;
wire x_14340;
wire x_14341;
wire x_14342;
wire x_14343;
wire x_14344;
wire x_14345;
wire x_14346;
wire x_14347;
wire x_14348;
wire x_14349;
wire x_14350;
wire x_14351;
wire x_14352;
wire x_14353;
wire x_14354;
wire x_14355;
wire x_14356;
wire x_14357;
wire x_14358;
wire x_14359;
wire x_14360;
wire x_14361;
wire x_14362;
wire x_14363;
wire x_14364;
wire x_14365;
wire x_14366;
wire x_14367;
wire x_14368;
wire x_14369;
wire x_14370;
wire x_14371;
wire x_14372;
wire x_14373;
wire x_14374;
wire x_14375;
wire x_14376;
wire x_14377;
wire x_14378;
wire x_14379;
wire x_14380;
wire x_14381;
wire x_14382;
wire x_14383;
wire x_14384;
wire x_14385;
wire x_14386;
wire x_14387;
wire x_14388;
wire x_14389;
wire x_14390;
wire x_14391;
wire x_14392;
wire x_14393;
wire x_14394;
wire x_14395;
wire x_14396;
wire x_14397;
wire x_14398;
wire x_14399;
wire x_14400;
wire x_14401;
wire x_14402;
wire x_14403;
wire x_14404;
wire x_14405;
wire x_14406;
wire x_14407;
wire x_14408;
wire x_14409;
wire x_14410;
wire x_14411;
wire x_14412;
wire x_14413;
wire x_14414;
wire x_14415;
wire x_14416;
wire x_14417;
wire x_14418;
wire x_14419;
wire x_14420;
wire x_14421;
wire x_14422;
wire x_14423;
wire x_14424;
wire x_14425;
wire x_14426;
wire x_14427;
wire x_14428;
wire x_14429;
wire x_14430;
wire x_14431;
wire x_14432;
wire x_14433;
wire x_14434;
wire x_14435;
wire x_14436;
wire x_14437;
wire x_14438;
wire x_14439;
wire x_14440;
wire x_14441;
wire x_14442;
wire x_14443;
wire x_14444;
wire x_14445;
wire x_14446;
wire x_14447;
wire x_14448;
wire x_14449;
wire x_14450;
wire x_14451;
wire x_14452;
wire x_14453;
wire x_14454;
wire x_14455;
wire x_14456;
wire x_14457;
wire x_14458;
wire x_14459;
wire x_14460;
wire x_14461;
wire x_14462;
wire x_14463;
wire x_14464;
wire x_14465;
wire x_14466;
wire x_14467;
wire x_14468;
wire x_14469;
wire x_14470;
wire x_14471;
wire x_14472;
wire x_14473;
wire x_14474;
wire x_14475;
wire x_14476;
wire x_14477;
wire x_14478;
wire x_14479;
wire x_14480;
wire x_14481;
wire x_14482;
wire x_14483;
wire x_14484;
wire x_14485;
wire x_14486;
wire x_14487;
wire x_14488;
wire x_14489;
wire x_14490;
wire x_14491;
wire x_14492;
wire x_14493;
wire x_14494;
wire x_14495;
wire x_14496;
wire x_14497;
wire x_14498;
wire x_14499;
wire x_14500;
wire x_14501;
wire x_14502;
wire x_14503;
wire x_14504;
wire x_14505;
wire x_14506;
wire x_14507;
wire x_14508;
wire x_14509;
wire x_14510;
wire x_14511;
wire x_14512;
wire x_14513;
wire x_14514;
wire x_14515;
wire x_14516;
wire x_14517;
wire x_14518;
wire x_14519;
wire x_14520;
wire x_14521;
wire x_14522;
wire x_14523;
wire x_14524;
wire x_14525;
wire x_14526;
wire x_14527;
wire x_14528;
wire x_14529;
wire x_14530;
wire x_14531;
wire x_14532;
wire x_14533;
wire x_14534;
wire x_14535;
wire x_14536;
wire x_14537;
wire x_14538;
wire x_14539;
wire x_14540;
wire x_14541;
wire x_14542;
wire x_14543;
wire x_14544;
wire x_14545;
wire x_14546;
wire x_14547;
wire x_14548;
wire x_14549;
wire x_14550;
wire x_14551;
wire x_14552;
wire x_14553;
wire x_14554;
wire x_14555;
wire x_14556;
wire x_14557;
wire x_14558;
wire x_14559;
wire x_14560;
wire x_14561;
wire x_14562;
wire x_14563;
wire x_14564;
wire x_14565;
wire x_14566;
wire x_14567;
wire x_14568;
wire x_14569;
wire x_14570;
wire x_14571;
wire x_14572;
wire x_14573;
wire x_14574;
wire x_14575;
wire x_14576;
wire x_14577;
wire x_14578;
wire x_14579;
wire x_14580;
wire x_14581;
wire x_14582;
wire x_14583;
wire x_14584;
wire x_14585;
wire x_14586;
wire x_14587;
wire x_14588;
wire x_14589;
wire x_14590;
wire x_14591;
wire x_14592;
wire x_14593;
wire x_14594;
wire x_14595;
wire x_14596;
wire x_14597;
wire x_14598;
wire x_14599;
wire x_14600;
wire x_14601;
wire x_14602;
wire x_14603;
wire x_14604;
wire x_14605;
wire x_14606;
wire x_14607;
wire x_14608;
wire x_14609;
wire x_14610;
wire x_14611;
wire x_14612;
wire x_14613;
wire x_14614;
wire x_14615;
wire x_14616;
wire x_14617;
wire x_14618;
wire x_14619;
wire x_14620;
wire x_14621;
wire x_14622;
wire x_14623;
wire x_14624;
wire x_14625;
wire x_14626;
wire x_14627;
wire x_14628;
wire x_14629;
wire x_14630;
wire x_14631;
wire x_14632;
wire x_14633;
wire x_14634;
wire x_14635;
wire x_14636;
wire x_14637;
wire x_14638;
wire x_14639;
wire x_14640;
wire x_14641;
wire x_14642;
wire x_14643;
wire x_14644;
wire x_14645;
wire x_14646;
wire x_14647;
wire x_14648;
wire x_14649;
wire x_14650;
wire x_14651;
wire x_14652;
wire x_14653;
wire x_14654;
wire x_14655;
wire x_14656;
wire x_14657;
wire x_14658;
wire x_14659;
wire x_14660;
wire x_14661;
wire x_14662;
wire x_14663;
wire x_14664;
wire x_14665;
wire x_14666;
wire x_14667;
wire x_14668;
wire x_14669;
wire x_14670;
wire x_14671;
wire x_14672;
wire x_14673;
wire x_14674;
wire x_14675;
wire x_14676;
wire x_14677;
wire x_14678;
wire x_14679;
wire x_14680;
wire x_14681;
wire x_14682;
wire x_14683;
wire x_14684;
wire x_14685;
wire x_14686;
wire x_14687;
wire x_14688;
wire x_14689;
wire x_14690;
wire x_14691;
wire x_14692;
wire x_14693;
wire x_14694;
wire x_14695;
wire x_14696;
wire x_14697;
wire x_14698;
wire x_14699;
wire x_14700;
wire x_14701;
wire x_14702;
wire x_14703;
wire x_14704;
wire x_14705;
wire x_14706;
wire x_14707;
wire x_14708;
wire x_14709;
wire x_14710;
wire x_14711;
wire x_14712;
wire x_14713;
wire x_14714;
wire x_14715;
wire x_14716;
wire x_14717;
wire x_14718;
wire x_14719;
wire x_14720;
wire x_14721;
wire x_14722;
wire x_14723;
wire x_14724;
wire x_14725;
wire x_14726;
wire x_14727;
wire x_14728;
wire x_14729;
wire x_14730;
wire x_14731;
wire x_14732;
wire x_14733;
wire x_14734;
wire x_14735;
wire x_14736;
wire x_14737;
wire x_14738;
wire x_14739;
wire x_14740;
wire x_14741;
wire x_14742;
wire x_14743;
wire x_14744;
wire x_14745;
wire x_14746;
wire x_14747;
wire x_14748;
wire x_14749;
wire x_14750;
wire x_14751;
wire x_14752;
wire x_14753;
wire x_14754;
wire x_14755;
wire x_14756;
wire x_14757;
wire x_14758;
wire x_14759;
wire x_14760;
wire x_14761;
wire x_14762;
wire x_14763;
wire x_14764;
wire x_14765;
wire x_14766;
wire x_14767;
wire x_14768;
wire x_14769;
wire x_14770;
wire x_14771;
wire x_14772;
wire x_14773;
wire x_14774;
wire x_14775;
wire x_14776;
wire x_14777;
wire x_14778;
wire x_14779;
wire x_14780;
wire x_14781;
wire x_14782;
wire x_14783;
wire x_14784;
wire x_14785;
wire x_14786;
wire x_14787;
wire x_14788;
wire x_14789;
wire x_14790;
wire x_14791;
wire x_14792;
wire x_14793;
wire x_14794;
wire x_14795;
wire x_14796;
wire x_14797;
wire x_14798;
wire x_14799;
wire x_14800;
wire x_14801;
wire x_14802;
wire x_14803;
wire x_14804;
wire x_14805;
wire x_14806;
wire x_14807;
wire x_14808;
wire x_14809;
wire x_14810;
wire x_14811;
wire x_14812;
wire x_14813;
wire x_14814;
wire x_14815;
wire x_14816;
wire x_14817;
wire x_14818;
wire x_14819;
wire x_14820;
wire x_14821;
wire x_14822;
wire x_14823;
wire x_14824;
wire x_14825;
wire x_14826;
wire x_14827;
wire x_14828;
wire x_14829;
wire x_14830;
wire x_14831;
wire x_14832;
wire x_14833;
wire x_14834;
wire x_14835;
wire x_14836;
wire x_14837;
wire x_14838;
wire x_14839;
wire x_14840;
wire x_14841;
wire x_14842;
wire x_14843;
wire x_14844;
wire x_14845;
wire x_14846;
wire x_14847;
wire x_14848;
wire x_14849;
wire x_14850;
wire x_14851;
wire x_14852;
wire x_14853;
wire x_14854;
wire x_14855;
wire x_14856;
wire x_14857;
wire x_14858;
wire x_14859;
wire x_14860;
wire x_14861;
wire x_14862;
wire x_14863;
wire x_14864;
wire x_14865;
wire x_14866;
wire x_14867;
wire x_14868;
wire x_14869;
wire x_14870;
wire x_14871;
wire x_14872;
wire x_14873;
wire x_14874;
wire x_14875;
wire x_14876;
wire x_14877;
wire x_14878;
wire x_14879;
wire x_14880;
wire x_14881;
wire x_14882;
wire x_14883;
wire x_14884;
wire x_14885;
wire x_14886;
wire x_14887;
wire x_14888;
wire x_14889;
wire x_14890;
wire x_14891;
wire x_14892;
wire x_14893;
wire x_14894;
wire x_14895;
wire x_14896;
wire x_14897;
wire x_14898;
wire x_14899;
wire x_14900;
wire x_14901;
wire x_14902;
wire x_14903;
wire x_14904;
wire x_14905;
wire x_14906;
wire x_14907;
wire x_14908;
wire x_14909;
wire x_14910;
wire x_14911;
wire x_14912;
wire x_14913;
wire x_14914;
wire x_14915;
wire x_14916;
wire x_14917;
wire x_14918;
wire x_14919;
wire x_14920;
wire x_14921;
wire x_14922;
wire x_14923;
wire x_14924;
wire x_14925;
wire x_14926;
wire x_14927;
wire x_14928;
wire x_14929;
wire x_14930;
wire x_14931;
wire x_14932;
wire x_14933;
wire x_14934;
wire x_14935;
wire x_14936;
wire x_14937;
wire x_14938;
wire x_14939;
wire x_14940;
wire x_14941;
wire x_14942;
wire x_14943;
wire x_14944;
wire x_14945;
wire x_14946;
wire x_14947;
wire x_14948;
wire x_14949;
wire x_14950;
wire x_14951;
wire x_14952;
wire x_14953;
wire x_14954;
wire x_14955;
wire x_14956;
wire x_14957;
wire x_14958;
wire x_14959;
wire x_14960;
wire x_14961;
wire x_14962;
wire x_14963;
wire x_14964;
wire x_14965;
wire x_14966;
wire x_14967;
wire x_14968;
wire x_14969;
wire x_14970;
wire x_14971;
wire x_14972;
wire x_14973;
wire x_14974;
wire x_14975;
wire x_14976;
wire x_14977;
wire x_14978;
wire x_14979;
wire x_14980;
wire x_14981;
wire x_14982;
wire x_14983;
wire x_14984;
wire x_14985;
wire x_14986;
wire x_14987;
wire x_14988;
wire x_14989;
wire x_14990;
wire x_14991;
wire x_14992;
wire x_14993;
wire x_14994;
wire x_14995;
wire x_14996;
wire x_14997;
wire x_14998;
wire x_14999;
wire x_15000;
wire x_15001;
wire x_15002;
wire x_15003;
wire x_15004;
wire x_15005;
wire x_15006;
wire x_15007;
wire x_15008;
wire x_15009;
wire x_15010;
wire x_15011;
wire x_15012;
wire x_15013;
wire x_15014;
wire x_15015;
wire x_15016;
wire x_15017;
wire x_15018;
wire x_15019;
wire x_15020;
wire x_15021;
wire x_15022;
wire x_15023;
wire x_15024;
wire x_15025;
wire x_15026;
wire x_15027;
wire x_15028;
wire x_15029;
wire x_15030;
wire x_15031;
wire x_15032;
wire x_15033;
wire x_15034;
wire x_15035;
wire x_15036;
wire x_15037;
wire x_15038;
wire x_15039;
wire x_15040;
wire x_15041;
wire x_15042;
wire x_15043;
wire x_15044;
wire x_15045;
wire x_15046;
wire x_15047;
wire x_15048;
wire x_15049;
wire x_15050;
wire x_15051;
wire x_15052;
wire x_15053;
wire x_15054;
wire x_15055;
wire x_15056;
wire x_15057;
wire x_15058;
wire x_15059;
wire x_15060;
wire x_15061;
wire x_15062;
wire x_15063;
wire x_15064;
wire x_15065;
wire x_15066;
wire x_15067;
wire x_15068;
wire x_15069;
wire x_15070;
wire x_15071;
wire x_15072;
wire x_15073;
wire x_15074;
wire x_15075;
wire x_15076;
wire x_15077;
wire x_15078;
wire x_15079;
wire x_15080;
wire x_15081;
wire x_15082;
wire x_15083;
wire x_15084;
wire x_15085;
wire x_15086;
wire x_15087;
wire x_15088;
wire x_15089;
wire x_15090;
wire x_15091;
wire x_15092;
wire x_15093;
wire x_15094;
wire x_15095;
wire x_15096;
wire x_15097;
wire x_15098;
wire x_15099;
wire x_15100;
wire x_15101;
wire x_15102;
wire x_15103;
wire x_15104;
wire x_15105;
wire x_15106;
wire x_15107;
wire x_15108;
wire x_15109;
wire x_15110;
wire x_15111;
wire x_15112;
wire x_15113;
wire x_15114;
wire x_15115;
wire x_15116;
wire x_15117;
wire x_15118;
wire x_15119;
wire x_15120;
wire x_15121;
wire x_15122;
wire x_15123;
wire x_15124;
wire x_15125;
wire x_15126;
wire x_15127;
wire x_15128;
wire x_15129;
wire x_15130;
wire x_15131;
wire x_15132;
wire x_15133;
wire x_15134;
wire x_15135;
wire x_15136;
wire x_15137;
wire x_15138;
wire x_15139;
wire x_15140;
wire x_15141;
wire x_15142;
wire x_15143;
wire x_15144;
wire x_15145;
wire x_15146;
wire x_15147;
wire x_15148;
wire x_15149;
wire x_15150;
wire x_15151;
wire x_15152;
wire x_15153;
wire x_15154;
wire x_15155;
wire x_15156;
wire x_15157;
wire x_15158;
wire x_15159;
wire x_15160;
wire x_15161;
wire x_15162;
wire x_15163;
wire x_15164;
wire x_15165;
wire x_15166;
wire x_15167;
wire x_15168;
wire x_15169;
wire x_15170;
wire x_15171;
wire x_15172;
wire x_15173;
wire x_15174;
wire x_15175;
wire x_15176;
wire x_15177;
wire x_15178;
wire x_15179;
wire x_15180;
wire x_15181;
wire x_15182;
wire x_15183;
wire x_15184;
wire x_15185;
wire x_15186;
wire x_15187;
wire x_15188;
wire x_15189;
wire x_15190;
wire x_15191;
wire x_15192;
wire x_15193;
wire x_15194;
wire x_15195;
wire x_15196;
wire x_15197;
wire x_15198;
wire x_15199;
wire x_15200;
wire x_15201;
wire x_15202;
wire x_15203;
wire x_15204;
wire x_15205;
wire x_15206;
wire x_15207;
wire x_15208;
wire x_15209;
wire x_15210;
wire x_15211;
wire x_15212;
wire x_15213;
wire x_15214;
wire x_15215;
wire x_15216;
wire x_15217;
wire x_15218;
wire x_15219;
wire x_15220;
wire x_15221;
wire x_15222;
wire x_15223;
wire x_15224;
wire x_15225;
wire x_15226;
wire x_15227;
wire x_15228;
wire x_15229;
wire x_15230;
wire x_15231;
wire x_15232;
wire x_15233;
wire x_15234;
wire x_15235;
wire x_15236;
wire x_15237;
wire x_15238;
wire x_15239;
wire x_15240;
wire x_15241;
wire x_15242;
wire x_15243;
wire x_15244;
wire x_15245;
wire x_15246;
wire x_15247;
wire x_15248;
wire x_15249;
wire x_15250;
wire x_15251;
wire x_15252;
wire x_15253;
wire x_15254;
wire x_15255;
wire x_15256;
wire x_15257;
wire x_15258;
wire x_15259;
wire x_15260;
wire x_15261;
wire x_15262;
wire x_15263;
wire x_15264;
wire x_15265;
wire x_15266;
wire x_15267;
wire x_15268;
wire x_15269;
wire x_15270;
wire x_15271;
wire x_15272;
wire x_15273;
wire x_15274;
wire x_15275;
wire x_15276;
wire x_15277;
wire x_15278;
wire x_15279;
wire x_15280;
wire x_15281;
wire x_15282;
wire x_15283;
wire x_15284;
wire x_15285;
wire x_15286;
wire x_15287;
wire x_15288;
wire x_15289;
wire x_15290;
wire x_15291;
wire x_15292;
wire x_15293;
wire x_15294;
wire x_15295;
wire x_15296;
wire x_15297;
wire x_15298;
wire x_15299;
wire x_15300;
wire x_15301;
wire x_15302;
wire x_15303;
wire x_15304;
wire x_15305;
wire x_15306;
wire x_15307;
wire x_15308;
wire x_15309;
wire x_15310;
wire x_15311;
wire x_15312;
wire x_15313;
wire x_15314;
wire x_15315;
wire x_15316;
wire x_15317;
wire x_15318;
wire x_15319;
wire x_15320;
wire x_15321;
wire x_15322;
wire x_15323;
wire x_15324;
wire x_15325;
wire x_15326;
wire x_15327;
wire x_15328;
wire x_15329;
wire x_15330;
wire x_15331;
wire x_15332;
wire x_15333;
wire x_15334;
wire x_15335;
wire x_15336;
wire x_15337;
wire x_15338;
wire x_15339;
wire x_15340;
wire x_15341;
wire x_15342;
wire x_15343;
wire x_15344;
wire x_15345;
wire x_15346;
wire x_15347;
wire x_15348;
wire x_15349;
wire x_15350;
wire x_15351;
wire x_15352;
wire x_15353;
wire x_15354;
wire x_15355;
wire x_15356;
wire x_15357;
wire x_15358;
wire x_15359;
wire x_15360;
wire x_15361;
wire x_15362;
wire x_15363;
wire x_15364;
wire x_15365;
wire x_15366;
wire x_15367;
wire x_15368;
wire x_15369;
wire x_15370;
wire x_15371;
wire x_15372;
wire x_15373;
wire x_15374;
wire x_15375;
wire x_15376;
wire x_15377;
wire x_15378;
wire x_15379;
wire x_15380;
wire x_15381;
wire x_15382;
wire x_15383;
wire x_15384;
wire x_15385;
wire x_15386;
wire x_15387;
wire x_15388;
wire x_15389;
wire x_15390;
wire x_15391;
wire x_15392;
wire x_15393;
wire x_15394;
wire x_15395;
wire x_15396;
wire x_15397;
wire x_15398;
wire x_15399;
wire x_15400;
wire x_15401;
wire x_15402;
wire x_15403;
wire x_15404;
wire x_15405;
wire x_15406;
wire x_15407;
wire x_15408;
wire x_15409;
wire x_15410;
wire x_15411;
wire x_15412;
wire x_15413;
wire x_15414;
wire x_15415;
wire x_15416;
wire x_15417;
wire x_15418;
wire x_15419;
wire x_15420;
wire x_15421;
wire x_15422;
wire x_15423;
wire x_15424;
wire x_15425;
wire x_15426;
wire x_15427;
wire x_15428;
wire x_15429;
wire x_15430;
wire x_15431;
wire x_15432;
wire x_15433;
wire x_15434;
wire x_15435;
wire x_15436;
wire x_15437;
wire x_15438;
wire x_15439;
wire x_15440;
wire x_15441;
wire x_15442;
wire x_15443;
wire x_15444;
wire x_15445;
wire x_15446;
wire x_15447;
wire x_15448;
wire x_15449;
wire x_15450;
wire x_15451;
wire x_15452;
wire x_15453;
wire x_15454;
wire x_15455;
wire x_15456;
wire x_15457;
wire x_15458;
wire x_15459;
wire x_15460;
wire x_15461;
wire x_15462;
wire x_15463;
wire x_15464;
wire x_15465;
wire x_15466;
wire x_15467;
wire x_15468;
wire x_15469;
wire x_15470;
wire x_15471;
wire x_15472;
wire x_15473;
wire x_15474;
wire x_15475;
wire x_15476;
wire x_15477;
wire x_15478;
wire x_15479;
wire x_15480;
wire x_15481;
wire x_15482;
wire x_15483;
wire x_15484;
wire x_15485;
wire x_15486;
wire x_15487;
wire x_15488;
wire x_15489;
wire x_15490;
wire x_15491;
wire x_15492;
wire x_15493;
wire x_15494;
wire x_15495;
wire x_15496;
wire x_15497;
wire x_15498;
wire x_15499;
wire x_15500;
wire x_15501;
wire x_15502;
wire x_15503;
wire x_15504;
wire x_15505;
wire x_15506;
wire x_15507;
wire x_15508;
wire x_15509;
wire x_15510;
wire x_15511;
wire x_15512;
wire x_15513;
wire x_15514;
wire x_15515;
wire x_15516;
wire x_15517;
wire x_15518;
wire x_15519;
wire x_15520;
wire x_15521;
wire x_15522;
wire x_15523;
wire x_15524;
wire x_15525;
wire x_15526;
wire x_15527;
wire x_15528;
wire x_15529;
wire x_15530;
wire x_15531;
wire x_15532;
wire x_15533;
wire x_15534;
wire x_15535;
wire x_15536;
wire x_15537;
wire x_15538;
wire x_15539;
wire x_15540;
wire x_15541;
wire x_15542;
wire x_15543;
wire x_15544;
wire x_15545;
wire x_15546;
wire x_15547;
wire x_15548;
wire x_15549;
wire x_15550;
wire x_15551;
wire x_15552;
wire x_15553;
wire x_15554;
wire x_15555;
wire x_15556;
wire x_15557;
wire x_15558;
wire x_15559;
wire x_15560;
wire x_15561;
wire x_15562;
wire x_15563;
wire x_15564;
wire x_15565;
wire x_15566;
wire x_15567;
wire x_15568;
wire x_15569;
wire x_15570;
wire x_15571;
wire x_15572;
wire x_15573;
wire x_15574;
wire x_15575;
wire x_15576;
wire x_15577;
wire x_15578;
wire x_15579;
wire x_15580;
wire x_15581;
wire x_15582;
wire x_15583;
wire x_15584;
wire x_15585;
wire x_15586;
wire x_15587;
wire x_15588;
wire x_15589;
wire x_15590;
wire x_15591;
wire x_15592;
wire x_15593;
wire x_15594;
wire x_15595;
wire x_15596;
wire x_15597;
wire x_15598;
wire x_15599;
wire x_15600;
wire x_15601;
wire x_15602;
wire x_15603;
wire x_15604;
wire x_15605;
wire x_15606;
wire x_15607;
wire x_15608;
wire x_15609;
wire x_15610;
wire x_15611;
wire x_15612;
wire x_15613;
wire x_15614;
wire x_15615;
wire x_15616;
wire x_15617;
wire x_15618;
wire x_15619;
wire x_15620;
wire x_15621;
wire x_15622;
wire x_15623;
wire x_15624;
wire x_15625;
wire x_15626;
wire x_15627;
wire x_15628;
wire x_15629;
wire x_15630;
wire x_15631;
wire x_15632;
wire x_15633;
wire x_15634;
wire x_15635;
wire x_15636;
wire x_15637;
wire x_15638;
wire x_15639;
wire x_15640;
wire x_15641;
wire x_15642;
wire x_15643;
wire x_15644;
wire x_15645;
wire x_15646;
wire x_15647;
wire x_15648;
wire x_15649;
wire x_15650;
wire x_15651;
wire x_15652;
wire x_15653;
wire x_15654;
wire x_15655;
wire x_15656;
wire x_15657;
wire x_15658;
wire x_15659;
wire x_15660;
wire x_15661;
wire x_15662;
wire x_15663;
wire x_15664;
wire x_15665;
wire x_15666;
wire x_15667;
wire x_15668;
wire x_15669;
wire x_15670;
wire x_15671;
wire x_15672;
wire x_15673;
wire x_15674;
wire x_15675;
wire x_15676;
wire x_15677;
wire x_15678;
wire x_15679;
wire x_15680;
wire x_15681;
wire x_15682;
wire x_15683;
wire x_15684;
wire x_15685;
wire x_15686;
wire x_15687;
wire x_15688;
wire x_15689;
wire x_15690;
wire x_15691;
wire x_15692;
wire x_15693;
wire x_15694;
wire x_15695;
wire x_15696;
wire x_15697;
wire x_15698;
wire x_15699;
wire x_15700;
wire x_15701;
wire x_15702;
wire x_15703;
wire x_15704;
wire x_15705;
wire x_15706;
wire x_15707;
wire x_15708;
wire x_15709;
wire x_15710;
wire x_15711;
wire x_15712;
wire x_15713;
wire x_15714;
wire x_15715;
wire x_15716;
wire x_15717;
wire x_15718;
wire x_15719;
wire x_15720;
wire x_15721;
wire x_15722;
wire x_15723;
wire x_15724;
wire x_15725;
wire x_15726;
wire x_15727;
wire x_15728;
wire x_15729;
wire x_15730;
wire x_15731;
wire x_15732;
wire x_15733;
wire x_15734;
wire x_15735;
wire x_15736;
wire x_15737;
wire x_15738;
wire x_15739;
wire x_15740;
wire x_15741;
wire x_15742;
wire x_15743;
wire x_15744;
wire x_15745;
wire x_15746;
wire x_15747;
wire x_15748;
wire x_15749;
wire x_15750;
wire x_15751;
wire x_15752;
wire x_15753;
wire x_15754;
wire x_15755;
wire x_15756;
wire x_15757;
wire x_15758;
wire x_15759;
wire x_15760;
wire x_15761;
wire x_15762;
wire x_15763;
wire x_15764;
wire x_15765;
wire x_15766;
wire x_15767;
wire x_15768;
wire x_15769;
wire x_15770;
wire x_15771;
wire x_15772;
wire x_15773;
wire x_15774;
wire x_15775;
wire x_15776;
wire x_15777;
wire x_15778;
wire x_15779;
wire x_15780;
wire x_15781;
wire x_15782;
wire x_15783;
wire x_15784;
wire x_15785;
wire x_15786;
wire x_15787;
wire x_15788;
wire x_15789;
wire x_15790;
wire x_15791;
wire x_15792;
wire x_15793;
wire x_15794;
wire x_15795;
wire x_15796;
wire x_15797;
wire x_15798;
wire x_15799;
wire x_15800;
wire x_15801;
wire x_15802;
wire x_15803;
wire x_15804;
wire x_15805;
wire x_15806;
wire x_15807;
wire x_15808;
wire x_15809;
wire x_15810;
wire x_15811;
wire x_15812;
wire x_15813;
wire x_15814;
wire x_15815;
wire x_15816;
wire x_15817;
wire x_15818;
wire x_15819;
wire x_15820;
wire x_15821;
wire x_15822;
wire x_15823;
wire x_15824;
wire x_15825;
wire x_15826;
wire x_15827;
wire x_15828;
wire x_15829;
wire x_15830;
wire x_15831;
wire x_15832;
wire x_15833;
wire x_15834;
wire x_15835;
wire x_15836;
wire x_15837;
wire x_15838;
wire x_15839;
wire x_15840;
wire x_15841;
wire x_15842;
wire x_15843;
wire x_15844;
wire x_15845;
wire x_15846;
wire x_15847;
wire x_15848;
wire x_15849;
wire x_15850;
wire x_15851;
wire x_15852;
wire x_15853;
wire x_15854;
wire x_15855;
wire x_15856;
wire x_15857;
wire x_15858;
wire x_15859;
wire x_15860;
wire x_15861;
wire x_15862;
wire x_15863;
wire x_15864;
wire x_15865;
wire x_15866;
wire x_15867;
wire x_15868;
wire x_15869;
wire x_15870;
wire x_15871;
wire x_15872;
wire x_15873;
wire x_15874;
wire x_15875;
wire x_15876;
wire x_15877;
wire x_15878;
wire x_15879;
wire x_15880;
wire x_15881;
wire x_15882;
wire x_15883;
wire x_15884;
wire x_15885;
wire x_15886;
wire x_15887;
wire x_15888;
wire x_15889;
wire x_15890;
wire x_15891;
wire x_15892;
wire x_15893;
wire x_15894;
wire x_15895;
wire x_15896;
wire x_15897;
wire x_15898;
wire x_15899;
wire x_15900;
wire x_15901;
wire x_15902;
wire x_15903;
wire x_15904;
wire x_15905;
wire x_15906;
wire x_15907;
wire x_15908;
wire x_15909;
wire x_15910;
wire x_15911;
wire x_15912;
wire x_15913;
wire x_15914;
wire x_15915;
wire x_15916;
wire x_15917;
wire x_15918;
wire x_15919;
wire x_15920;
wire x_15921;
wire x_15922;
wire x_15923;
wire x_15924;
wire x_15925;
wire x_15926;
wire x_15927;
wire x_15928;
wire x_15929;
wire x_15930;
wire x_15931;
wire x_15932;
wire x_15933;
wire x_15934;
wire x_15935;
wire x_15936;
wire x_15937;
wire x_15938;
wire x_15939;
wire x_15940;
wire x_15941;
wire x_15942;
wire x_15943;
wire x_15944;
wire x_15945;
wire x_15946;
wire x_15947;
wire x_15948;
wire x_15949;
wire x_15950;
wire x_15951;
wire x_15952;
wire x_15953;
wire x_15954;
wire x_15955;
wire x_15956;
wire x_15957;
wire x_15958;
wire x_15959;
wire x_15960;
wire x_15961;
wire x_15962;
wire x_15963;
wire x_15964;
wire x_15965;
wire x_15966;
wire x_15967;
wire x_15968;
wire x_15969;
wire x_15970;
wire x_15971;
wire x_15972;
wire x_15973;
wire x_15974;
wire x_15975;
wire x_15976;
wire x_15977;
wire x_15978;
wire x_15979;
wire x_15980;
wire x_15981;
wire x_15982;
wire x_15983;
wire x_15984;
wire x_15985;
wire x_15986;
wire x_15987;
wire x_15988;
wire x_15989;
wire x_15990;
wire x_15991;
wire x_15992;
wire x_15993;
wire x_15994;
wire x_15995;
wire x_15996;
wire x_15997;
wire x_15998;
wire x_15999;
wire x_16000;
wire x_16001;
wire x_16002;
wire x_16003;
wire x_16004;
wire x_16005;
wire x_16006;
wire x_16007;
wire x_16008;
wire x_16009;
wire x_16010;
wire x_16011;
wire x_16012;
wire x_16013;
wire x_16014;
wire x_16015;
wire x_16016;
wire x_16017;
wire x_16018;
wire x_16019;
wire x_16020;
wire x_16021;
wire x_16022;
wire x_16023;
wire x_16024;
wire x_16025;
wire x_16026;
wire x_16027;
wire x_16028;
wire x_16029;
wire x_16030;
wire x_16031;
wire x_16032;
wire x_16033;
wire x_16034;
wire x_16035;
wire x_16036;
wire x_16037;
wire x_16038;
wire x_16039;
wire x_16040;
wire x_16041;
wire x_16042;
wire x_16043;
wire x_16044;
wire x_16045;
wire x_16046;
wire x_16047;
wire x_16048;
wire x_16049;
wire x_16050;
wire x_16051;
wire x_16052;
wire x_16053;
wire x_16054;
wire x_16055;
wire x_16056;
wire x_16057;
wire x_16058;
wire x_16059;
wire x_16060;
wire x_16061;
wire x_16062;
wire x_16063;
wire x_16064;
wire x_16065;
wire x_16066;
wire x_16067;
wire x_16068;
wire x_16069;
wire x_16070;
wire x_16071;
wire x_16072;
wire x_16073;
wire x_16074;
wire x_16075;
wire x_16076;
wire x_16077;
wire x_16078;
wire x_16079;
wire x_16080;
wire x_16081;
wire x_16082;
wire x_16083;
wire x_16084;
wire x_16085;
wire x_16086;
wire x_16087;
wire x_16088;
wire x_16089;
wire x_16090;
wire x_16091;
wire x_16092;
wire x_16093;
wire x_16094;
wire x_16095;
wire x_16096;
wire x_16097;
wire x_16098;
wire x_16099;
wire x_16100;
wire x_16101;
wire x_16102;
wire x_16103;
wire x_16104;
wire x_16105;
wire x_16106;
wire x_16107;
wire x_16108;
wire x_16109;
wire x_16110;
wire x_16111;
wire x_16112;
wire x_16113;
wire x_16114;
wire x_16115;
wire x_16116;
wire x_16117;
wire x_16118;
wire x_16119;
wire x_16120;
wire x_16121;
wire x_16122;
wire x_16123;
wire x_16124;
wire x_16125;
wire x_16126;
wire x_16127;
wire x_16128;
wire x_16129;
wire x_16130;
wire x_16131;
wire x_16132;
wire x_16133;
wire x_16134;
wire x_16135;
wire x_16136;
wire x_16137;
wire x_16138;
wire x_16139;
wire x_16140;
wire x_16141;
wire x_16142;
wire x_16143;
wire x_16144;
wire x_16145;
wire x_16146;
wire x_16147;
wire x_16148;
wire x_16149;
wire x_16150;
wire x_16151;
wire x_16152;
wire x_16153;
wire x_16154;
wire x_16155;
wire x_16156;
wire x_16157;
wire x_16158;
wire x_16159;
wire x_16160;
wire x_16161;
wire x_16162;
wire x_16163;
wire x_16164;
wire x_16165;
wire x_16166;
wire x_16167;
wire x_16168;
wire x_16169;
wire x_16170;
wire x_16171;
wire x_16172;
wire x_16173;
wire x_16174;
wire x_16175;
wire x_16176;
wire x_16177;
wire x_16178;
wire x_16179;
wire x_16180;
wire x_16181;
wire x_16182;
wire x_16183;
wire x_16184;
wire x_16185;
wire x_16186;
wire x_16187;
wire x_16188;
wire x_16189;
wire x_16190;
wire x_16191;
wire x_16192;
wire x_16193;
wire x_16194;
wire x_16195;
wire x_16196;
wire x_16197;
wire x_16198;
wire x_16199;
wire x_16200;
wire x_16201;
wire x_16202;
wire x_16203;
wire x_16204;
wire x_16205;
wire x_16206;
wire x_16207;
wire x_16208;
wire x_16209;
wire x_16210;
wire x_16211;
wire x_16212;
wire x_16213;
wire x_16214;
wire x_16215;
wire x_16216;
wire x_16217;
wire x_16218;
wire x_16219;
wire x_16220;
wire x_16221;
wire x_16222;
wire x_16223;
wire x_16224;
wire x_16225;
wire x_16226;
wire x_16227;
wire x_16228;
wire x_16229;
wire x_16230;
wire x_16231;
wire x_16232;
wire x_16233;
wire x_16234;
wire x_16235;
wire x_16236;
wire x_16237;
wire x_16238;
wire x_16239;
wire x_16240;
wire x_16241;
wire x_16242;
wire x_16243;
wire x_16244;
wire x_16245;
wire x_16246;
wire x_16247;
wire x_16248;
wire x_16249;
wire x_16250;
wire x_16251;
wire x_16252;
wire x_16253;
wire x_16254;
wire x_16255;
wire x_16256;
wire x_16257;
wire x_16258;
wire x_16259;
wire x_16260;
wire x_16261;
wire x_16262;
wire x_16263;
wire x_16264;
wire x_16265;
wire x_16266;
wire x_16267;
wire x_16268;
wire x_16269;
wire x_16270;
wire x_16271;
wire x_16272;
wire x_16273;
wire x_16274;
wire x_16275;
wire x_16276;
wire x_16277;
wire x_16278;
wire x_16279;
wire x_16280;
wire x_16281;
wire x_16282;
wire x_16283;
wire x_16284;
wire x_16285;
wire x_16286;
wire x_16287;
wire x_16288;
wire x_16289;
wire x_16290;
wire x_16291;
wire x_16292;
wire x_16293;
wire x_16294;
wire x_16295;
wire x_16296;
wire x_16297;
wire x_16298;
wire x_16299;
wire x_16300;
wire x_16301;
wire x_16302;
wire x_16303;
wire x_16304;
wire x_16305;
wire x_16306;
wire x_16307;
wire x_16308;
wire x_16309;
wire x_16310;
wire x_16311;
wire x_16312;
wire x_16313;
wire x_16314;
wire x_16315;
wire x_16316;
wire x_16317;
wire x_16318;
wire x_16319;
wire x_16320;
wire x_16321;
wire x_16322;
wire x_16323;
wire x_16324;
wire x_16325;
wire x_16326;
wire x_16327;
wire x_16328;
wire x_16329;
wire x_16330;
wire x_16331;
wire x_16332;
wire x_16333;
wire x_16334;
wire x_16335;
wire x_16336;
wire x_16337;
wire x_16338;
wire x_16339;
wire x_16340;
wire x_16341;
wire x_16342;
wire x_16343;
wire x_16344;
wire x_16345;
wire x_16346;
wire x_16347;
wire x_16348;
wire x_16349;
wire x_16350;
wire x_16351;
wire x_16352;
wire x_16353;
wire x_16354;
wire x_16355;
wire x_16356;
wire x_16357;
wire x_16358;
wire x_16359;
wire x_16360;
wire x_16361;
wire x_16362;
wire x_16363;
wire x_16364;
wire x_16365;
wire x_16366;
wire x_16367;
wire x_16368;
wire x_16369;
wire x_16370;
wire x_16371;
wire x_16372;
wire x_16373;
wire x_16374;
wire x_16375;
wire x_16376;
wire x_16377;
wire x_16378;
wire x_16379;
wire x_16380;
wire x_16381;
wire x_16382;
wire x_16383;
wire x_16384;
wire x_16385;
wire x_16386;
wire x_16387;
wire x_16388;
wire x_16389;
wire x_16390;
wire x_16391;
wire x_16392;
wire x_16393;
wire x_16394;
wire x_16395;
wire x_16396;
wire x_16397;
wire x_16398;
wire x_16399;
wire x_16400;
wire x_16401;
wire x_16402;
wire x_16403;
wire x_16404;
wire x_16405;
wire x_16406;
wire x_16407;
wire x_16408;
wire x_16409;
wire x_16410;
wire x_16411;
wire x_16412;
wire x_16413;
wire x_16414;
wire x_16415;
wire x_16416;
wire x_16417;
wire x_16418;
wire x_16419;
wire x_16420;
wire x_16421;
wire x_16422;
wire x_16423;
wire x_16424;
wire x_16425;
wire x_16426;
wire x_16427;
wire x_16428;
wire x_16429;
wire x_16430;
wire x_16431;
wire x_16432;
wire x_16433;
wire x_16434;
wire x_16435;
wire x_16436;
wire x_16437;
wire x_16438;
wire x_16439;
wire x_16440;
wire x_16441;
wire x_16442;
wire x_16443;
wire x_16444;
wire x_16445;
wire x_16446;
wire x_16447;
wire x_16448;
wire x_16449;
wire x_16450;
wire x_16451;
wire x_16452;
wire x_16453;
wire x_16454;
wire x_16455;
wire x_16456;
wire x_16457;
wire x_16458;
wire x_16459;
wire x_16460;
wire x_16461;
wire x_16462;
wire x_16463;
wire x_16464;
wire x_16465;
wire x_16466;
wire x_16467;
wire x_16468;
wire x_16469;
wire x_16470;
wire x_16471;
wire x_16472;
wire x_16473;
wire x_16474;
wire x_16475;
wire x_16476;
wire x_16477;
wire x_16478;
wire x_16479;
wire x_16480;
wire x_16481;
wire x_16482;
wire x_16483;
wire x_16484;
wire x_16485;
wire x_16486;
wire x_16487;
wire x_16488;
wire x_16489;
wire x_16490;
wire x_16491;
wire x_16492;
wire x_16493;
wire x_16494;
wire x_16495;
wire x_16496;
wire x_16497;
wire x_16498;
wire x_16499;
wire x_16500;
wire x_16501;
wire x_16502;
wire x_16503;
wire x_16504;
wire x_16505;
wire x_16506;
wire x_16507;
wire x_16508;
wire x_16509;
wire x_16510;
wire x_16511;
wire x_16512;
wire x_16513;
wire x_16514;
wire x_16515;
wire x_16516;
wire x_16517;
wire x_16518;
wire x_16519;
wire x_16520;
wire x_16521;
wire x_16522;
wire x_16523;
wire x_16524;
wire x_16525;
wire x_16526;
wire x_16527;
wire x_16528;
wire x_16529;
wire x_16530;
wire x_16531;
wire x_16532;
wire x_16533;
wire x_16534;
wire x_16535;
wire x_16536;
wire x_16537;
wire x_16538;
wire x_16539;
wire x_16540;
wire x_16541;
wire x_16542;
wire x_16543;
wire x_16544;
wire x_16545;
wire x_16546;
wire x_16547;
wire x_16548;
wire x_16549;
wire x_16550;
wire x_16551;
wire x_16552;
wire x_16553;
wire x_16554;
wire x_16555;
wire x_16556;
wire x_16557;
wire x_16558;
wire x_16559;
wire x_16560;
wire x_16561;
wire x_16562;
wire x_16563;
wire x_16564;
wire x_16565;
wire x_16566;
wire x_16567;
wire x_16568;
wire x_16569;
wire x_16570;
wire x_16571;
wire x_16572;
wire x_16573;
wire x_16574;
wire x_16575;
wire x_16576;
wire x_16577;
wire x_16578;
wire x_16579;
wire x_16580;
wire x_16581;
wire x_16582;
wire x_16583;
wire x_16584;
wire x_16585;
wire x_16586;
wire x_16587;
wire x_16588;
wire x_16589;
wire x_16590;
wire x_16591;
wire x_16592;
wire x_16593;
wire x_16594;
wire x_16595;
wire x_16596;
wire x_16597;
wire x_16598;
wire x_16599;
wire x_16600;
wire x_16601;
wire x_16602;
wire x_16603;
wire x_16604;
wire x_16605;
wire x_16606;
wire x_16607;
wire x_16608;
wire x_16609;
wire x_16610;
wire x_16611;
wire x_16612;
wire x_16613;
wire x_16614;
wire x_16615;
wire x_16616;
wire x_16617;
wire x_16618;
wire x_16619;
wire x_16620;
wire x_16621;
wire x_16622;
wire x_16623;
wire x_16624;
wire x_16625;
wire x_16626;
wire x_16627;
wire x_16628;
wire x_16629;
wire x_16630;
wire x_16631;
wire x_16632;
wire x_16633;
wire x_16634;
wire x_16635;
wire x_16636;
wire x_16637;
wire x_16638;
wire x_16639;
wire x_16640;
wire x_16641;
wire x_16642;
wire x_16643;
wire x_16644;
wire x_16645;
wire x_16646;
wire x_16647;
wire x_16648;
wire x_16649;
wire x_16650;
wire x_16651;
wire x_16652;
wire x_16653;
wire x_16654;
wire x_16655;
wire x_16656;
wire x_16657;
wire x_16658;
wire x_16659;
wire x_16660;
wire x_16661;
wire x_16662;
wire x_16663;
wire x_16664;
wire x_16665;
wire x_16666;
wire x_16667;
wire x_16668;
wire x_16669;
wire x_16670;
wire x_16671;
wire x_16672;
wire x_16673;
wire x_16674;
wire x_16675;
wire x_16676;
wire x_16677;
wire x_16678;
wire x_16679;
wire x_16680;
wire x_16681;
wire x_16682;
wire x_16683;
wire x_16684;
wire x_16685;
wire x_16686;
wire x_16687;
wire x_16688;
wire x_16689;
wire x_16690;
wire x_16691;
wire x_16692;
wire x_16693;
wire x_16694;
wire x_16695;
wire x_16696;
wire x_16697;
wire x_16698;
wire x_16699;
wire x_16700;
wire x_16701;
wire x_16702;
wire x_16703;
wire x_16704;
wire x_16705;
wire x_16706;
wire x_16707;
wire x_16708;
wire x_16709;
wire x_16710;
wire x_16711;
wire x_16712;
wire x_16713;
wire x_16714;
wire x_16715;
wire x_16716;
wire x_16717;
wire x_16718;
wire x_16719;
wire x_16720;
wire x_16721;
wire x_16722;
wire x_16723;
wire x_16724;
wire x_16725;
wire x_16726;
wire x_16727;
wire x_16728;
wire x_16729;
wire x_16730;
wire x_16731;
wire x_16732;
wire x_16733;
wire x_16734;
wire x_16735;
wire x_16736;
wire x_16737;
wire x_16738;
wire x_16739;
wire x_16740;
wire x_16741;
wire x_16742;
wire x_16743;
wire x_16744;
wire x_16745;
wire x_16746;
wire x_16747;
wire x_16748;
wire x_16749;
wire x_16750;
wire x_16751;
wire x_16752;
wire x_16753;
wire x_16754;
wire x_16755;
wire x_16756;
wire x_16757;
wire x_16758;
wire x_16759;
wire x_16760;
wire x_16761;
wire x_16762;
wire x_16763;
wire x_16764;
wire x_16765;
wire x_16766;
wire x_16767;
wire x_16768;
wire x_16769;
wire x_16770;
wire x_16771;
wire x_16772;
wire x_16773;
wire x_16774;
wire x_16775;
wire x_16776;
wire x_16777;
wire x_16778;
wire x_16779;
wire x_16780;
wire x_16781;
wire x_16782;
wire x_16783;
wire x_16784;
wire x_16785;
wire x_16786;
wire x_16787;
wire x_16788;
wire x_16789;
wire x_16790;
wire x_16791;
wire x_16792;
wire x_16793;
wire x_16794;
wire x_16795;
wire x_16796;
wire x_16797;
wire x_16798;
wire x_16799;
wire x_16800;
wire x_16801;
wire x_16802;
wire x_16803;
wire x_16804;
wire x_16805;
wire x_16806;
wire x_16807;
wire x_16808;
wire x_16809;
wire x_16810;
wire x_16811;
wire x_16812;
wire x_16813;
wire x_16814;
wire x_16815;
wire x_16816;
wire x_16817;
wire x_16818;
wire x_16819;
wire x_16820;
wire x_16821;
wire x_16822;
wire x_16823;
wire x_16824;
wire x_16825;
wire x_16826;
wire x_16827;
wire x_16828;
wire x_16829;
wire x_16830;
wire x_16831;
wire x_16832;
wire x_16833;
wire x_16834;
wire x_16835;
wire x_16836;
wire x_16837;
wire x_16838;
wire x_16839;
wire x_16840;
wire x_16841;
wire x_16842;
wire x_16843;
wire x_16844;
wire x_16845;
wire x_16846;
wire x_16847;
wire x_16848;
wire x_16849;
wire x_16850;
wire x_16851;
wire x_16852;
wire x_16853;
wire x_16854;
wire x_16855;
wire x_16856;
wire x_16857;
wire x_16858;
wire x_16859;
wire x_16860;
wire x_16861;
wire x_16862;
wire x_16863;
wire x_16864;
wire x_16865;
wire x_16866;
wire x_16867;
wire x_16868;
wire x_16869;
wire x_16870;
wire x_16871;
wire x_16872;
wire x_16873;
wire x_16874;
wire x_16875;
wire x_16876;
wire x_16877;
wire x_16878;
wire x_16879;
wire x_16880;
wire x_16881;
wire x_16882;
wire x_16883;
wire x_16884;
wire x_16885;
wire x_16886;
wire x_16887;
wire x_16888;
wire x_16889;
wire x_16890;
wire x_16891;
wire x_16892;
wire x_16893;
wire x_16894;
wire x_16895;
wire x_16896;
wire x_16897;
wire x_16898;
wire x_16899;
wire x_16900;
wire x_16901;
wire x_16902;
wire x_16903;
wire x_16904;
wire x_16905;
wire x_16906;
wire x_16907;
wire x_16908;
wire x_16909;
wire x_16910;
wire x_16911;
wire x_16912;
wire x_16913;
wire x_16914;
wire x_16915;
wire x_16916;
wire x_16917;
wire x_16918;
wire x_16919;
wire x_16920;
wire x_16921;
wire x_16922;
wire x_16923;
wire x_16924;
wire x_16925;
wire x_16926;
wire x_16927;
wire x_16928;
wire x_16929;
wire x_16930;
wire x_16931;
wire x_16932;
wire x_16933;
wire x_16934;
wire x_16935;
wire x_16936;
wire x_16937;
wire x_16938;
wire x_16939;
wire x_16940;
wire x_16941;
wire x_16942;
wire x_16943;
wire x_16944;
wire x_16945;
wire x_16946;
wire x_16947;
wire x_16948;
wire x_16949;
wire x_16950;
wire x_16951;
wire x_16952;
wire x_16953;
wire x_16954;
wire x_16955;
wire x_16956;
wire x_16957;
wire x_16958;
wire x_16959;
wire x_16960;
wire x_16961;
wire x_16962;
wire x_16963;
wire x_16964;
wire x_16965;
wire x_16966;
wire x_16967;
wire x_16968;
wire x_16969;
wire x_16970;
wire x_16971;
wire x_16972;
wire x_16973;
wire x_16974;
wire x_16975;
wire x_16976;
wire x_16977;
wire x_16978;
wire x_16979;
wire x_16980;
wire x_16981;
wire x_16982;
wire x_16983;
wire x_16984;
wire x_16985;
wire x_16986;
wire x_16987;
wire x_16988;
wire x_16989;
wire x_16990;
wire x_16991;
wire x_16992;
wire x_16993;
wire x_16994;
wire x_16995;
wire x_16996;
wire x_16997;
wire x_16998;
wire x_16999;
wire x_17000;
wire x_17001;
wire x_17002;
wire x_17003;
wire x_17004;
wire x_17005;
wire x_17006;
wire x_17007;
wire x_17008;
wire x_17009;
wire x_17010;
wire x_17011;
wire x_17012;
wire x_17013;
wire x_17014;
wire x_17015;
wire x_17016;
wire x_17017;
wire x_17018;
wire x_17019;
wire x_17020;
wire x_17021;
wire x_17022;
wire x_17023;
wire x_17024;
wire x_17025;
wire x_17026;
wire x_17027;
wire x_17028;
wire x_17029;
wire x_17030;
wire x_17031;
wire x_17032;
wire x_17033;
wire x_17034;
wire x_17035;
wire x_17036;
wire x_17037;
wire x_17038;
wire x_17039;
wire x_17040;
wire x_17041;
wire x_17042;
wire x_17043;
wire x_17044;
wire x_17045;
wire x_17046;
wire x_17047;
wire x_17048;
wire x_17049;
wire x_17050;
wire x_17051;
wire x_17052;
wire x_17053;
wire x_17054;
wire x_17055;
wire x_17056;
wire x_17057;
wire x_17058;
wire x_17059;
wire x_17060;
wire x_17061;
wire x_17062;
wire x_17063;
wire x_17064;
wire x_17065;
wire x_17066;
wire x_17067;
wire x_17068;
wire x_17069;
wire x_17070;
wire x_17071;
wire x_17072;
wire x_17073;
wire x_17074;
wire x_17075;
wire x_17076;
wire x_17077;
wire x_17078;
wire x_17079;
wire x_17080;
wire x_17081;
wire x_17082;
wire x_17083;
wire x_17084;
wire x_17085;
wire x_17086;
wire x_17087;
wire x_17088;
wire x_17089;
wire x_17090;
wire x_17091;
wire x_17092;
wire x_17093;
wire x_17094;
wire x_17095;
wire x_17096;
wire x_17097;
wire x_17098;
wire x_17099;
wire x_17100;
wire x_17101;
wire x_17102;
wire x_17103;
wire x_17104;
wire x_17105;
wire x_17106;
wire x_17107;
wire x_17108;
wire x_17109;
wire x_17110;
wire x_17111;
wire x_17112;
wire x_17113;
wire x_17114;
wire x_17115;
wire x_17116;
wire x_17117;
wire x_17118;
wire x_17119;
wire x_17120;
wire x_17121;
wire x_17122;
wire x_17123;
wire x_17124;
wire x_17125;
wire x_17126;
wire x_17127;
wire x_17128;
wire x_17129;
wire x_17130;
wire x_17131;
wire x_17132;
wire x_17133;
wire x_17134;
wire x_17135;
wire x_17136;
wire x_17137;
wire x_17138;
wire x_17139;
wire x_17140;
wire x_17141;
wire x_17142;
wire x_17143;
wire x_17144;
wire x_17145;
wire x_17146;
wire x_17147;
wire x_17148;
wire x_17149;
wire x_17150;
wire x_17151;
wire x_17152;
wire x_17153;
wire x_17154;
wire x_17155;
wire x_17156;
wire x_17157;
wire x_17158;
wire x_17159;
wire x_17160;
wire x_17161;
wire x_17162;
wire x_17163;
wire x_17164;
wire x_17165;
wire x_17166;
wire x_17167;
wire x_17168;
wire x_17169;
wire x_17170;
wire x_17171;
wire x_17172;
wire x_17173;
wire x_17174;
wire x_17175;
wire x_17176;
wire x_17177;
wire x_17178;
wire x_17179;
wire x_17180;
wire x_17181;
wire x_17182;
wire x_17183;
wire x_17184;
wire x_17185;
wire x_17186;
wire x_17187;
wire x_17188;
wire x_17189;
wire x_17190;
wire x_17191;
wire x_17192;
wire x_17193;
wire x_17194;
wire x_17195;
wire x_17196;
wire x_17197;
wire x_17198;
wire x_17199;
wire x_17200;
wire x_17201;
wire x_17202;
wire x_17203;
wire x_17204;
wire x_17205;
wire x_17206;
wire x_17207;
wire x_17208;
wire x_17209;
wire x_17210;
wire x_17211;
wire x_17212;
wire x_17213;
wire x_17214;
wire x_17215;
wire x_17216;
wire x_17217;
wire x_17218;
wire x_17219;
wire x_17220;
wire x_17221;
wire x_17222;
wire x_17223;
wire x_17224;
wire x_17225;
wire x_17226;
wire x_17227;
wire x_17228;
wire x_17229;
wire x_17230;
wire x_17231;
wire x_17232;
wire x_17233;
wire x_17234;
wire x_17235;
wire x_17236;
wire x_17237;
wire x_17238;
wire x_17239;
wire x_17240;
wire x_17241;
wire x_17242;
wire x_17243;
wire x_17244;
wire x_17245;
wire x_17246;
wire x_17247;
wire x_17248;
wire x_17249;
wire x_17250;
wire x_17251;
wire x_17252;
wire x_17253;
wire x_17254;
wire x_17255;
wire x_17256;
wire x_17257;
wire x_17258;
wire x_17259;
wire x_17260;
wire x_17261;
wire x_17262;
wire x_17263;
wire x_17264;
wire x_17265;
wire x_17266;
wire x_17267;
wire x_17268;
wire x_17269;
wire x_17270;
wire x_17271;
wire x_17272;
wire x_17273;
wire x_17274;
wire x_17275;
wire x_17276;
wire x_17277;
wire x_17278;
wire x_17279;
wire x_17280;
wire x_17281;
wire x_17282;
wire x_17283;
wire x_17284;
wire x_17285;
wire x_17286;
wire x_17287;
wire x_17288;
wire x_17289;
wire x_17290;
wire x_17291;
wire x_17292;
wire x_17293;
wire x_17294;
wire x_17295;
wire x_17296;
wire x_17297;
wire x_17298;
wire x_17299;
wire x_17300;
wire x_17301;
wire x_17302;
wire x_17303;
wire x_17304;
wire x_17305;
wire x_17306;
wire x_17307;
wire x_17308;
wire x_17309;
wire x_17310;
wire x_17311;
wire x_17312;
wire x_17313;
wire x_17314;
wire x_17315;
wire x_17316;
wire x_17317;
wire x_17318;
wire x_17319;
wire x_17320;
wire x_17321;
wire x_17322;
wire x_17323;
wire x_17324;
wire x_17325;
wire x_17326;
wire x_17327;
wire x_17328;
wire x_17329;
wire x_17330;
wire x_17331;
wire x_17332;
wire x_17333;
wire x_17334;
wire x_17335;
wire x_17336;
wire x_17337;
wire x_17338;
wire x_17339;
wire x_17340;
wire x_17341;
wire x_17342;
wire x_17343;
wire x_17344;
wire x_17345;
wire x_17346;
wire x_17347;
wire x_17348;
wire x_17349;
wire x_17350;
wire x_17351;
wire x_17352;
wire x_17353;
wire x_17354;
wire x_17355;
wire x_17356;
wire x_17357;
wire x_17358;
wire x_17359;
wire x_17360;
wire x_17361;
wire x_17362;
wire x_17363;
wire x_17364;
wire x_17365;
wire x_17366;
wire x_17367;
wire x_17368;
wire x_17369;
wire x_17370;
wire x_17371;
wire x_17372;
wire x_17373;
wire x_17374;
wire x_17375;
wire x_17376;
wire x_17377;
wire x_17378;
wire x_17379;
wire x_17380;
wire x_17381;
wire x_17382;
wire x_17383;
wire x_17384;
wire x_17385;
wire x_17386;
wire x_17387;
wire x_17388;
wire x_17389;
wire x_17390;
wire x_17391;
wire x_17392;
wire x_17393;
wire x_17394;
wire x_17395;
wire x_17396;
wire x_17397;
wire x_17398;
wire x_17399;
wire x_17400;
wire x_17401;
wire x_17402;
wire x_17403;
wire x_17404;
wire x_17405;
wire x_17406;
wire x_17407;
wire x_17408;
wire x_17409;
wire x_17410;
wire x_17411;
wire x_17412;
wire x_17413;
wire x_17414;
wire x_17415;
wire x_17416;
wire x_17417;
wire x_17418;
wire x_17419;
wire x_17420;
wire x_17421;
wire x_17422;
wire x_17423;
wire x_17424;
wire x_17425;
wire x_17426;
wire x_17427;
wire x_17428;
wire x_17429;
wire x_17430;
wire x_17431;
wire x_17432;
wire x_17433;
wire x_17434;
wire x_17435;
wire x_17436;
wire x_17437;
wire x_17438;
wire x_17439;
wire x_17440;
wire x_17441;
wire x_17442;
wire x_17443;
wire x_17444;
wire x_17445;
wire x_17446;
wire x_17447;
wire x_17448;
wire x_17449;
wire x_17450;
wire x_17451;
wire x_17452;
wire x_17453;
wire x_17454;
wire x_17455;
wire x_17456;
wire x_17457;
wire x_17458;
wire x_17459;
wire x_17460;
wire x_17461;
wire x_17462;
wire x_17463;
wire x_17464;
wire x_17465;
wire x_17466;
wire x_17467;
wire x_17468;
wire x_17469;
wire x_17470;
wire x_17471;
wire x_17472;
wire x_17473;
wire x_17474;
wire x_17475;
wire x_17476;
wire x_17477;
wire x_17478;
wire x_17479;
wire x_17480;
wire x_17481;
wire x_17482;
wire x_17483;
wire x_17484;
wire x_17485;
wire x_17486;
wire x_17487;
wire x_17488;
wire x_17489;
wire x_17490;
wire x_17491;
wire x_17492;
wire x_17493;
wire x_17494;
wire x_17495;
wire x_17496;
wire x_17497;
wire x_17498;
wire x_17499;
wire x_17500;
wire x_17501;
wire x_17502;
wire x_17503;
wire x_17504;
wire x_17505;
wire x_17506;
wire x_17507;
wire x_17508;
wire x_17509;
wire x_17510;
wire x_17511;
wire x_17512;
wire x_17513;
wire x_17514;
wire x_17515;
wire x_17516;
wire x_17517;
wire x_17518;
wire x_17519;
wire x_17520;
wire x_17521;
wire x_17522;
wire x_17523;
wire x_17524;
wire x_17525;
wire x_17526;
wire x_17527;
wire x_17528;
wire x_17529;
wire x_17530;
wire x_17531;
wire x_17532;
wire x_17533;
wire x_17534;
wire x_17535;
wire x_17536;
wire x_17537;
wire x_17538;
wire x_17539;
wire x_17540;
wire x_17541;
wire x_17542;
wire x_17543;
wire x_17544;
wire x_17545;
wire x_17546;
wire x_17547;
wire x_17548;
wire x_17549;
wire x_17550;
wire x_17551;
wire x_17552;
wire x_17553;
wire x_17554;
wire x_17555;
wire x_17556;
wire x_17557;
wire x_17558;
wire x_17559;
wire x_17560;
wire x_17561;
wire x_17562;
wire x_17563;
wire x_17564;
wire x_17565;
wire x_17566;
wire x_17567;
wire x_17568;
wire x_17569;
wire x_17570;
wire x_17571;
wire x_17572;
wire x_17573;
wire x_17574;
wire x_17575;
wire x_17576;
wire x_17577;
wire x_17578;
wire x_17579;
wire x_17580;
wire x_17581;
wire x_17582;
wire x_17583;
wire x_17584;
wire x_17585;
wire x_17586;
wire x_17587;
wire x_17588;
wire x_17589;
wire x_17590;
wire x_17591;
wire x_17592;
wire x_17593;
wire x_17594;
wire x_17595;
wire x_17596;
wire x_17597;
wire x_17598;
wire x_17599;
wire x_17600;
wire x_17601;
wire x_17602;
wire x_17603;
wire x_17604;
wire x_17605;
wire x_17606;
wire x_17607;
wire x_17608;
wire x_17609;
wire x_17610;
wire x_17611;
wire x_17612;
wire x_17613;
wire x_17614;
wire x_17615;
wire x_17616;
wire x_17617;
wire x_17618;
wire x_17619;
wire x_17620;
wire x_17621;
wire x_17622;
wire x_17623;
wire x_17624;
wire x_17625;
wire x_17626;
wire x_17627;
wire x_17628;
wire x_17629;
wire x_17630;
wire x_17631;
wire x_17632;
wire x_17633;
wire x_17634;
wire x_17635;
wire x_17636;
wire x_17637;
wire x_17638;
wire x_17639;
wire x_17640;
wire x_17641;
wire x_17642;
wire x_17643;
wire x_17644;
wire x_17645;
wire x_17646;
wire x_17647;
wire x_17648;
wire x_17649;
wire x_17650;
wire x_17651;
wire x_17652;
wire x_17653;
wire x_17654;
wire x_17655;
wire x_17656;
wire x_17657;
wire x_17658;
wire x_17659;
wire x_17660;
wire x_17661;
wire x_17662;
wire x_17663;
wire x_17664;
wire x_17665;
wire x_17666;
wire x_17667;
wire x_17668;
wire x_17669;
wire x_17670;
wire x_17671;
wire x_17672;
wire x_17673;
wire x_17674;
wire x_17675;
wire x_17676;
wire x_17677;
wire x_17678;
wire x_17679;
wire x_17680;
wire x_17681;
wire x_17682;
wire x_17683;
wire x_17684;
wire x_17685;
wire x_17686;
wire x_17687;
wire x_17688;
wire x_17689;
wire x_17690;
wire x_17691;
wire x_17692;
wire x_17693;
wire x_17694;
wire x_17695;
wire x_17696;
wire x_17697;
wire x_17698;
wire x_17699;
wire x_17700;
wire x_17701;
wire x_17702;
wire x_17703;
wire x_17704;
wire x_17705;
wire x_17706;
wire x_17707;
wire x_17708;
wire x_17709;
wire x_17710;
wire x_17711;
wire x_17712;
wire x_17713;
wire x_17714;
wire x_17715;
wire x_17716;
wire x_17717;
wire x_17718;
wire x_17719;
wire x_17720;
wire x_17721;
wire x_17722;
wire x_17723;
wire x_17724;
wire x_17725;
wire x_17726;
wire x_17727;
wire x_17728;
wire x_17729;
wire x_17730;
wire x_17731;
wire x_17732;
wire x_17733;
wire x_17734;
wire x_17735;
wire x_17736;
wire x_17737;
wire x_17738;
wire x_17739;
wire x_17740;
wire x_17741;
wire x_17742;
wire x_17743;
wire x_17744;
wire x_17745;
wire x_17746;
wire x_17747;
wire x_17748;
wire x_17749;
wire x_17750;
wire x_17751;
wire x_17752;
wire x_17753;
wire x_17754;
wire x_17755;
wire x_17756;
wire x_17757;
wire x_17758;
wire x_17759;
wire x_17760;
wire x_17761;
wire x_17762;
wire x_17763;
wire x_17764;
wire x_17765;
wire x_17766;
wire x_17767;
wire x_17768;
wire x_17769;
wire x_17770;
wire x_17771;
wire x_17772;
wire x_17773;
wire x_17774;
wire x_17775;
wire x_17776;
wire x_17777;
wire x_17778;
wire x_17779;
wire x_17780;
wire x_17781;
wire x_17782;
wire x_17783;
wire x_17784;
wire x_17785;
wire x_17786;
wire x_17787;
wire x_17788;
wire x_17789;
wire x_17790;
wire x_17791;
wire x_17792;
wire x_17793;
wire x_17794;
wire x_17795;
wire x_17796;
wire x_17797;
wire x_17798;
wire x_17799;
wire x_17800;
wire x_17801;
wire x_17802;
wire x_17803;
wire x_17804;
wire x_17805;
wire x_17806;
wire x_17807;
wire x_17808;
wire x_17809;
wire x_17810;
wire x_17811;
wire x_17812;
wire x_17813;
wire x_17814;
wire x_17815;
wire x_17816;
wire x_17817;
wire x_17818;
wire x_17819;
wire x_17820;
wire x_17821;
wire x_17822;
wire x_17823;
wire x_17824;
wire x_17825;
wire x_17826;
wire x_17827;
wire x_17828;
wire x_17829;
wire x_17830;
wire x_17831;
wire x_17832;
wire x_17833;
wire x_17834;
wire x_17835;
wire x_17836;
wire x_17837;
wire x_17838;
wire x_17839;
wire x_17840;
wire x_17841;
wire x_17842;
wire x_17843;
wire x_17844;
wire x_17845;
wire x_17846;
wire x_17847;
wire x_17848;
wire x_17849;
wire x_17850;
wire x_17851;
wire x_17852;
wire x_17853;
wire x_17854;
wire x_17855;
wire x_17856;
wire x_17857;
wire x_17858;
wire x_17859;
wire x_17860;
wire x_17861;
wire x_17862;
wire x_17863;
wire x_17864;
wire x_17865;
wire x_17866;
wire x_17867;
wire x_17868;
wire x_17869;
wire x_17870;
wire x_17871;
wire x_17872;
wire x_17873;
wire x_17874;
wire x_17875;
wire x_17876;
wire x_17877;
wire x_17878;
wire x_17879;
wire x_17880;
wire x_17881;
wire x_17882;
wire x_17883;
wire x_17884;
wire x_17885;
wire x_17886;
wire x_17887;
wire x_17888;
wire x_17889;
wire x_17890;
wire x_17891;
wire x_17892;
wire x_17893;
wire x_17894;
wire x_17895;
wire x_17896;
wire x_17897;
wire x_17898;
wire x_17899;
wire x_17900;
wire x_17901;
wire x_17902;
wire x_17903;
wire x_17904;
wire x_17905;
wire x_17906;
wire x_17907;
wire x_17908;
wire x_17909;
wire x_17910;
wire x_17911;
wire x_17912;
wire x_17913;
wire x_17914;
wire x_17915;
wire x_17916;
wire x_17917;
wire x_17918;
wire x_17919;
wire x_17920;
wire x_17921;
wire x_17922;
wire x_17923;
wire x_17924;
wire x_17925;
wire x_17926;
wire x_17927;
wire x_17928;
wire x_17929;
wire x_17930;
wire x_17931;
wire x_17932;
wire x_17933;
wire x_17934;
wire x_17935;
wire x_17936;
wire x_17937;
wire x_17938;
wire x_17939;
wire x_17940;
wire x_17941;
wire x_17942;
wire x_17943;
wire x_17944;
wire x_17945;
wire x_17946;
wire x_17947;
wire x_17948;
wire x_17949;
wire x_17950;
wire x_17951;
wire x_17952;
wire x_17953;
wire x_17954;
wire x_17955;
wire x_17956;
wire x_17957;
wire x_17958;
wire x_17959;
wire x_17960;
wire x_17961;
wire x_17962;
wire x_17963;
wire x_17964;
wire x_17965;
wire x_17966;
wire x_17967;
wire x_17968;
wire x_17969;
wire x_17970;
wire x_17971;
wire x_17972;
wire x_17973;
wire x_17974;
wire x_17975;
wire x_17976;
wire x_17977;
wire x_17978;
wire x_17979;
wire x_17980;
wire x_17981;
wire x_17982;
wire x_17983;
wire x_17984;
wire x_17985;
wire x_17986;
wire x_17987;
wire x_17988;
wire x_17989;
wire x_17990;
wire x_17991;
wire x_17992;
wire x_17993;
wire x_17994;
wire x_17995;
wire x_17996;
wire x_17997;
wire x_17998;
wire x_17999;
wire x_18000;
wire x_18001;
wire x_18002;
wire x_18003;
wire x_18004;
wire x_18005;
wire x_18006;
wire x_18007;
wire x_18008;
wire x_18009;
wire x_18010;
wire x_18011;
wire x_18012;
wire x_18013;
wire x_18014;
wire x_18015;
wire x_18016;
wire x_18017;
wire x_18018;
wire x_18019;
wire x_18020;
wire x_18021;
wire x_18022;
wire x_18023;
wire x_18024;
wire x_18025;
wire x_18026;
wire x_18027;
wire x_18028;
wire x_18029;
wire x_18030;
wire x_18031;
wire x_18032;
wire x_18033;
wire x_18034;
wire x_18035;
wire x_18036;
wire x_18037;
wire x_18038;
wire x_18039;
wire x_18040;
wire x_18041;
wire x_18042;
wire x_18043;
wire x_18044;
wire x_18045;
wire x_18046;
wire x_18047;
wire x_18048;
wire x_18049;
wire x_18050;
wire x_18051;
wire x_18052;
wire x_18053;
wire x_18054;
wire x_18055;
wire x_18056;
wire x_18057;
wire x_18058;
wire x_18059;
wire x_18060;
wire x_18061;
wire x_18062;
wire x_18063;
wire x_18064;
wire x_18065;
wire x_18066;
wire x_18067;
wire x_18068;
wire x_18069;
wire x_18070;
wire x_18071;
wire x_18072;
wire x_18073;
wire x_18074;
wire x_18075;
wire x_18076;
wire x_18077;
wire x_18078;
wire x_18079;
wire x_18080;
wire x_18081;
wire x_18082;
wire x_18083;
wire x_18084;
wire x_18085;
wire x_18086;
wire x_18087;
wire x_18088;
wire x_18089;
wire x_18090;
wire x_18091;
wire x_18092;
wire x_18093;
wire x_18094;
wire x_18095;
wire x_18096;
wire x_18097;
wire x_18098;
wire x_18099;
wire x_18100;
wire x_18101;
wire x_18102;
wire x_18103;
wire x_18104;
wire x_18105;
wire x_18106;
wire x_18107;
wire x_18108;
wire x_18109;
wire x_18110;
wire x_18111;
wire x_18112;
wire x_18113;
wire x_18114;
wire x_18115;
wire x_18116;
wire x_18117;
wire x_18118;
wire x_18119;
wire x_18120;
wire x_18121;
wire x_18122;
wire x_18123;
wire x_18124;
wire x_18125;
wire x_18126;
wire x_18127;
wire x_18128;
wire x_18129;
wire x_18130;
wire x_18131;
wire x_18132;
wire x_18133;
wire x_18134;
wire x_18135;
wire x_18136;
wire x_18137;
wire x_18138;
wire x_18139;
wire x_18140;
wire x_18141;
wire x_18142;
wire x_18143;
wire x_18144;
wire x_18145;
wire x_18146;
wire x_18147;
wire x_18148;
wire x_18149;
wire x_18150;
wire x_18151;
wire x_18152;
wire x_18153;
wire x_18154;
wire x_18155;
wire x_18156;
wire x_18157;
wire x_18158;
wire x_18159;
wire x_18160;
wire x_18161;
wire x_18162;
wire x_18163;
wire x_18164;
wire x_18165;
wire x_18166;
wire x_18167;
wire x_18168;
wire x_18169;
wire x_18170;
wire x_18171;
wire x_18172;
wire x_18173;
wire x_18174;
wire x_18175;
wire x_18176;
wire x_18177;
wire x_18178;
wire x_18179;
wire x_18180;
wire x_18181;
wire x_18182;
wire x_18183;
wire x_18184;
wire x_18185;
wire x_18186;
wire x_18187;
wire x_18188;
wire x_18189;
wire x_18190;
wire x_18191;
wire x_18192;
wire x_18193;
wire x_18194;
wire x_18195;
wire x_18196;
wire x_18197;
wire x_18198;
wire x_18199;
wire x_18200;
wire x_18201;
wire x_18202;
wire x_18203;
wire x_18204;
wire x_18205;
wire x_18206;
wire x_18207;
wire x_18208;
wire x_18209;
wire x_18210;
wire x_18211;
wire x_18212;
wire x_18213;
wire x_18214;
wire x_18215;
wire x_18216;
wire x_18217;
wire x_18218;
wire x_18219;
wire x_18220;
wire x_18221;
wire x_18222;
wire x_18223;
wire x_18224;
wire x_18225;
wire x_18226;
wire x_18227;
wire x_18228;
wire x_18229;
wire x_18230;
wire x_18231;
wire x_18232;
wire x_18233;
wire x_18234;
wire x_18235;
wire x_18236;
wire x_18237;
wire x_18238;
wire x_18239;
wire x_18240;
wire x_18241;
wire x_18242;
wire x_18243;
wire x_18244;
wire x_18245;
wire x_18246;
wire x_18247;
wire x_18248;
wire x_18249;
wire x_18250;
wire x_18251;
wire x_18252;
wire x_18253;
wire x_18254;
wire x_18255;
wire x_18256;
wire x_18257;
wire x_18258;
wire x_18259;
wire x_18260;
wire x_18261;
wire x_18262;
wire x_18263;
wire x_18264;
wire x_18265;
wire x_18266;
wire x_18267;
wire x_18268;
wire x_18269;
wire x_18270;
wire x_18271;
wire x_18272;
wire x_18273;
wire x_18274;
wire x_18275;
wire x_18276;
wire x_18277;
wire x_18278;
wire x_18279;
wire x_18280;
wire x_18281;
wire x_18282;
wire x_18283;
wire x_18284;
wire x_18285;
wire x_18286;
wire x_18287;
wire x_18288;
wire x_18289;
wire x_18290;
wire x_18291;
wire x_18292;
wire x_18293;
wire x_18294;
wire x_18295;
wire x_18296;
wire x_18297;
wire x_18298;
wire x_18299;
wire x_18300;
wire x_18301;
wire x_18302;
wire x_18303;
wire x_18304;
wire x_18305;
wire x_18306;
wire x_18307;
wire x_18308;
wire x_18309;
wire x_18310;
wire x_18311;
wire x_18312;
wire x_18313;
wire x_18314;
wire x_18315;
wire x_18316;
wire x_18317;
wire x_18318;
wire x_18319;
wire x_18320;
wire x_18321;
wire x_18322;
wire x_18323;
wire x_18324;
wire x_18325;
wire x_18326;
wire x_18327;
wire x_18328;
wire x_18329;
wire x_18330;
wire x_18331;
wire x_18332;
wire x_18333;
wire x_18334;
wire x_18335;
wire x_18336;
wire x_18337;
wire x_18338;
wire x_18339;
wire x_18340;
wire x_18341;
wire x_18342;
wire x_18343;
wire x_18344;
wire x_18345;
wire x_18346;
wire x_18347;
wire x_18348;
wire x_18349;
wire x_18350;
wire x_18351;
wire x_18352;
wire x_18353;
wire x_18354;
wire x_18355;
wire x_18356;
wire x_18357;
wire x_18358;
wire x_18359;
wire x_18360;
wire x_18361;
wire x_18362;
wire x_18363;
wire x_18364;
wire x_18365;
wire x_18366;
wire x_18367;
wire x_18368;
wire x_18369;
wire x_18370;
wire x_18371;
wire x_18372;
wire x_18373;
wire x_18374;
wire x_18375;
wire x_18376;
wire x_18377;
wire x_18378;
wire x_18379;
wire x_18380;
wire x_18381;
wire x_18382;
wire x_18383;
wire x_18384;
wire x_18385;
wire x_18386;
wire x_18387;
wire x_18388;
wire x_18389;
wire x_18390;
wire x_18391;
wire x_18392;
wire x_18393;
wire x_18394;
wire x_18395;
wire x_18396;
wire x_18397;
wire x_18398;
wire x_18399;
wire x_18400;
wire x_18401;
wire x_18402;
wire x_18403;
wire x_18404;
wire x_18405;
wire x_18406;
wire x_18407;
wire x_18408;
wire x_18409;
wire x_18410;
wire x_18411;
wire x_18412;
wire x_18413;
wire x_18414;
wire x_18415;
wire x_18416;
wire x_18417;
wire x_18418;
wire x_18419;
wire x_18420;
wire x_18421;
wire x_18422;
wire x_18423;
wire x_18424;
wire x_18425;
wire x_18426;
wire x_18427;
wire x_18428;
wire x_18429;
wire x_18430;
wire x_18431;
wire x_18432;
wire x_18433;
wire x_18434;
wire x_18435;
wire x_18436;
wire x_18437;
wire x_18438;
wire x_18439;
wire x_18440;
wire x_18441;
wire x_18442;
wire x_18443;
wire x_18444;
wire x_18445;
wire x_18446;
wire x_18447;
wire x_18448;
wire x_18449;
wire x_18450;
wire x_18451;
wire x_18452;
wire x_18453;
wire x_18454;
wire x_18455;
wire x_18456;
wire x_18457;
wire x_18458;
wire x_18459;
wire x_18460;
wire x_18461;
wire x_18462;
wire x_18463;
wire x_18464;
wire x_18465;
wire x_18466;
wire x_18467;
wire x_18468;
wire x_18469;
wire x_18470;
wire x_18471;
wire x_18472;
wire x_18473;
wire x_18474;
wire x_18475;
wire x_18476;
wire x_18477;
wire x_18478;
wire x_18479;
wire x_18480;
wire x_18481;
wire x_18482;
wire x_18483;
wire x_18484;
wire x_18485;
wire x_18486;
wire x_18487;
wire x_18488;
wire x_18489;
wire x_18490;
wire x_18491;
wire x_18492;
wire x_18493;
wire x_18494;
wire x_18495;
wire x_18496;
wire x_18497;
wire x_18498;
wire x_18499;
wire x_18500;
wire x_18501;
wire x_18502;
wire x_18503;
wire x_18504;
wire x_18505;
wire x_18506;
wire x_18507;
wire x_18508;
wire x_18509;
wire x_18510;
wire x_18511;
wire x_18512;
wire x_18513;
wire x_18514;
wire x_18515;
wire x_18516;
wire x_18517;
wire x_18518;
wire x_18519;
wire x_18520;
wire x_18521;
wire x_18522;
wire x_18523;
wire x_18524;
wire x_18525;
wire x_18526;
wire x_18527;
wire x_18528;
wire x_18529;
wire x_18530;
wire x_18531;
wire x_18532;
wire x_18533;
wire x_18534;
wire x_18535;
wire x_18536;
wire x_18537;
wire x_18538;
wire x_18539;
wire x_18540;
wire x_18541;
wire x_18542;
wire x_18543;
wire x_18544;
wire x_18545;
wire x_18546;
wire x_18547;
wire x_18548;
wire x_18549;
wire x_18550;
wire x_18551;
wire x_18552;
wire x_18553;
wire x_18554;
wire x_18555;
wire x_18556;
wire x_18557;
wire x_18558;
wire x_18559;
wire x_18560;
wire x_18561;
wire x_18562;
wire x_18563;
wire x_18564;
wire x_18565;
wire x_18566;
wire x_18567;
wire x_18568;
wire x_18569;
wire x_18570;
wire x_18571;
wire x_18572;
wire x_18573;
wire x_18574;
wire x_18575;
wire x_18576;
wire x_18577;
wire x_18578;
wire x_18579;
wire x_18580;
wire x_18581;
wire x_18582;
wire x_18583;
wire x_18584;
wire x_18585;
wire x_18586;
wire x_18587;
wire x_18588;
wire x_18589;
wire x_18590;
wire x_18591;
wire x_18592;
wire x_18593;
wire x_18594;
wire x_18595;
wire x_18596;
wire x_18597;
wire x_18598;
wire x_18599;
wire x_18600;
wire x_18601;
wire x_18602;
wire x_18603;
wire x_18604;
wire x_18605;
wire x_18606;
wire x_18607;
wire x_18608;
wire x_18609;
wire x_18610;
wire x_18611;
wire x_18612;
wire x_18613;
wire x_18614;
wire x_18615;
wire x_18616;
wire x_18617;
wire x_18618;
wire x_18619;
wire x_18620;
wire x_18621;
wire x_18622;
wire x_18623;
wire x_18624;
wire x_18625;
wire x_18626;
wire x_18627;
wire x_18628;
wire x_18629;
wire x_18630;
wire x_18631;
wire x_18632;
wire x_18633;
wire x_18634;
wire x_18635;
wire x_18636;
wire x_18637;
wire x_18638;
wire x_18639;
wire x_18640;
wire x_18641;
wire x_18642;
wire x_18643;
wire x_18644;
wire x_18645;
wire x_18646;
wire x_18647;
wire x_18648;
wire x_18649;
wire x_18650;
wire x_18651;
wire x_18652;
wire x_18653;
wire x_18654;
wire x_18655;
wire x_18656;
wire x_18657;
wire x_18658;
wire x_18659;
wire x_18660;
wire x_18661;
wire x_18662;
wire x_18663;
wire x_18664;
wire x_18665;
wire x_18666;
wire x_18667;
wire x_18668;
wire x_18669;
wire x_18670;
wire x_18671;
wire x_18672;
wire x_18673;
wire x_18674;
wire x_18675;
wire x_18676;
wire x_18677;
wire x_18678;
wire x_18679;
wire x_18680;
wire x_18681;
wire x_18682;
wire x_18683;
wire x_18684;
wire x_18685;
wire x_18686;
wire x_18687;
wire x_18688;
wire x_18689;
wire x_18690;
wire x_18691;
wire x_18692;
wire x_18693;
wire x_18694;
wire x_18695;
wire x_18696;
wire x_18697;
wire x_18698;
wire x_18699;
wire x_18700;
wire x_18701;
wire x_18702;
wire x_18703;
wire x_18704;
wire x_18705;
wire x_18706;
wire x_18707;
wire x_18708;
wire x_18709;
wire x_18710;
wire x_18711;
wire x_18712;
wire x_18713;
wire x_18714;
wire x_18715;
wire x_18716;
wire x_18717;
wire x_18718;
wire x_18719;
wire x_18720;
wire x_18721;
wire x_18722;
wire x_18723;
wire x_18724;
wire x_18725;
wire x_18726;
wire x_18727;
wire x_18728;
wire x_18729;
wire x_18730;
wire x_18731;
wire x_18732;
wire x_18733;
wire x_18734;
wire x_18735;
wire x_18736;
wire x_18737;
wire x_18738;
wire x_18739;
wire x_18740;
wire x_18741;
wire x_18742;
wire x_18743;
wire x_18744;
wire x_18745;
wire x_18746;
wire x_18747;
wire x_18748;
wire x_18749;
wire x_18750;
wire x_18751;
wire x_18752;
wire x_18753;
wire x_18754;
wire x_18755;
wire x_18756;
wire x_18757;
wire x_18758;
wire x_18759;
wire x_18760;
wire x_18761;
wire x_18762;
wire x_18763;
wire x_18764;
wire x_18765;
wire x_18766;
wire x_18767;
wire x_18768;
wire x_18769;
wire x_18770;
wire x_18771;
wire x_18772;
wire x_18773;
wire x_18774;
wire x_18775;
wire x_18776;
wire x_18777;
wire x_18778;
wire x_18779;
wire x_18780;
wire x_18781;
wire x_18782;
wire x_18783;
wire x_18784;
wire x_18785;
wire x_18786;
wire x_18787;
wire x_18788;
wire x_18789;
wire x_18790;
wire x_18791;
wire x_18792;
wire x_18793;
wire x_18794;
wire x_18795;
wire x_18796;
wire x_18797;
wire x_18798;
wire x_18799;
wire x_18800;
wire x_18801;
wire x_18802;
wire x_18803;
wire x_18804;
wire x_18805;
wire x_18806;
wire x_18807;
wire x_18808;
wire x_18809;
wire x_18810;
wire x_18811;
wire x_18812;
wire x_18813;
wire x_18814;
wire x_18815;
wire x_18816;
wire x_18817;
wire x_18818;
wire x_18819;
wire x_18820;
wire x_18821;
wire x_18822;
wire x_18823;
wire x_18824;
wire x_18825;
wire x_18826;
wire x_18827;
wire x_18828;
wire x_18829;
wire x_18830;
wire x_18831;
wire x_18832;
wire x_18833;
wire x_18834;
wire x_18835;
wire x_18836;
wire x_18837;
wire x_18838;
wire x_18839;
wire x_18840;
wire x_18841;
wire x_18842;
wire x_18843;
wire x_18844;
wire x_18845;
wire x_18846;
wire x_18847;
wire x_18848;
wire x_18849;
wire x_18850;
wire x_18851;
wire x_18852;
wire x_18853;
wire x_18854;
wire x_18855;
wire x_18856;
wire x_18857;
wire x_18858;
wire x_18859;
wire x_18860;
wire x_18861;
wire x_18862;
wire x_18863;
wire x_18864;
wire x_18865;
wire x_18866;
wire x_18867;
wire x_18868;
wire x_18869;
wire x_18870;
wire x_18871;
wire x_18872;
wire x_18873;
wire x_18874;
wire x_18875;
wire x_18876;
wire x_18877;
wire x_18878;
wire x_18879;
wire x_18880;
wire x_18881;
wire x_18882;
wire x_18883;
wire x_18884;
wire x_18885;
wire x_18886;
wire x_18887;
wire x_18888;
wire x_18889;
wire x_18890;
wire x_18891;
wire x_18892;
wire x_18893;
wire x_18894;
wire x_18895;
wire x_18896;
wire x_18897;
wire x_18898;
wire x_18899;
wire x_18900;
wire x_18901;
wire x_18902;
wire x_18903;
wire x_18904;
wire x_18905;
wire x_18906;
wire x_18907;
wire x_18908;
wire x_18909;
wire x_18910;
wire x_18911;
wire x_18912;
wire x_18913;
wire x_18914;
wire x_18915;
wire x_18916;
wire x_18917;
wire x_18918;
wire x_18919;
wire x_18920;
wire x_18921;
wire x_18922;
wire x_18923;
wire x_18924;
wire x_18925;
wire x_18926;
wire x_18927;
wire x_18928;
wire x_18929;
wire x_18930;
wire x_18931;
wire x_18932;
wire x_18933;
wire x_18934;
wire x_18935;
wire x_18936;
wire x_18937;
wire x_18938;
wire x_18939;
wire x_18940;
wire x_18941;
wire x_18942;
wire x_18943;
wire x_18944;
wire x_18945;
wire x_18946;
wire x_18947;
wire x_18948;
wire x_18949;
wire x_18950;
wire x_18951;
wire x_18952;
wire x_18953;
wire x_18954;
wire x_18955;
wire x_18956;
wire x_18957;
wire x_18958;
wire x_18959;
wire x_18960;
wire x_18961;
wire x_18962;
wire x_18963;
wire x_18964;
wire x_18965;
wire x_18966;
wire x_18967;
wire x_18968;
wire x_18969;
wire x_18970;
wire x_18971;
wire x_18972;
wire x_18973;
wire x_18974;
wire x_18975;
wire x_18976;
wire x_18977;
wire x_18978;
wire x_18979;
wire x_18980;
wire x_18981;
wire x_18982;
wire x_18983;
wire x_18984;
wire x_18985;
wire x_18986;
wire x_18987;
wire x_18988;
wire x_18989;
wire x_18990;
wire x_18991;
wire x_18992;
wire x_18993;
wire x_18994;
wire x_18995;
wire x_18996;
wire x_18997;
wire x_18998;
wire x_18999;
wire x_19000;
wire x_19001;
wire x_19002;
wire x_19003;
wire x_19004;
wire x_19005;
wire x_19006;
wire x_19007;
wire x_19008;
wire x_19009;
wire x_19010;
wire x_19011;
wire x_19012;
wire x_19013;
wire x_19014;
wire x_19015;
wire x_19016;
wire x_19017;
wire x_19018;
wire x_19019;
wire x_19020;
wire x_19021;
wire x_19022;
wire x_19023;
wire x_19024;
wire x_19025;
wire x_19026;
wire x_19027;
wire x_19028;
wire x_19029;
wire x_19030;
wire x_19031;
wire x_19032;
wire x_19033;
wire x_19034;
wire x_19035;
wire x_19036;
wire x_19037;
wire x_19038;
wire x_19039;
wire x_19040;
wire x_19041;
wire x_19042;
wire x_19043;
wire x_19044;
wire x_19045;
wire x_19046;
wire x_19047;
wire x_19048;
wire x_19049;
wire x_19050;
wire x_19051;
wire x_19052;
wire x_19053;
wire x_19054;
wire x_19055;
wire x_19056;
wire x_19057;
wire x_19058;
wire x_19059;
wire x_19060;
wire x_19061;
wire x_19062;
wire x_19063;
wire x_19064;
wire x_19065;
wire x_19066;
wire x_19067;
wire x_19068;
wire x_19069;
wire x_19070;
wire x_19071;
wire x_19072;
wire x_19073;
wire x_19074;
wire x_19075;
wire x_19076;
wire x_19077;
wire x_19078;
wire x_19079;
wire x_19080;
wire x_19081;
wire x_19082;
wire x_19083;
wire x_19084;
wire x_19085;
wire x_19086;
wire x_19087;
wire x_19088;
wire x_19089;
wire x_19090;
wire x_19091;
wire x_19092;
wire x_19093;
wire x_19094;
wire x_19095;
wire x_19096;
wire x_19097;
wire x_19098;
wire x_19099;
wire x_19100;
wire x_19101;
wire x_19102;
wire x_19103;
wire x_19104;
wire x_19105;
wire x_19106;
wire x_19107;
wire x_19108;
wire x_19109;
wire x_19110;
wire x_19111;
wire x_19112;
wire x_19113;
wire x_19114;
wire x_19115;
wire x_19116;
wire x_19117;
wire x_19118;
wire x_19119;
wire x_19120;
wire x_19121;
wire x_19122;
wire x_19123;
wire x_19124;
wire x_19125;
wire x_19126;
wire x_19127;
wire x_19128;
wire x_19129;
wire x_19130;
wire x_19131;
wire x_19132;
wire x_19133;
wire x_19134;
wire x_19135;
wire x_19136;
wire x_19137;
wire x_19138;
wire x_19139;
wire x_19140;
wire x_19141;
wire x_19142;
wire x_19143;
wire x_19144;
wire x_19145;
wire x_19146;
wire x_19147;
wire x_19148;
wire x_19149;
wire x_19150;
wire x_19151;
wire x_19152;
wire x_19153;
wire x_19154;
wire x_19155;
wire x_19156;
wire x_19157;
wire x_19158;
wire x_19159;
wire x_19160;
wire x_19161;
wire x_19162;
wire x_19163;
wire x_19164;
wire x_19165;
wire x_19166;
wire x_19167;
wire x_19168;
wire x_19169;
wire x_19170;
wire x_19171;
wire x_19172;
wire x_19173;
wire x_19174;
wire x_19175;
wire x_19176;
wire x_19177;
wire x_19178;
wire x_19179;
wire x_19180;
wire x_19181;
wire x_19182;
wire x_19183;
wire x_19184;
wire x_19185;
wire x_19186;
wire x_19187;
wire x_19188;
wire x_19189;
wire x_19190;
wire x_19191;
wire x_19192;
wire x_19193;
wire x_19194;
wire x_19195;
wire x_19196;
wire x_19197;
wire x_19198;
wire x_19199;
wire x_19200;
wire x_19201;
wire x_19202;
wire x_19203;
wire x_19204;
wire x_19205;
wire x_19206;
wire x_19207;
wire x_19208;
wire x_19209;
wire x_19210;
wire x_19211;
wire x_19212;
wire x_19213;
wire x_19214;
wire x_19215;
wire x_19216;
wire x_19217;
wire x_19218;
wire x_19219;
wire x_19220;
wire x_19221;
wire x_19222;
wire x_19223;
wire x_19224;
wire x_19225;
wire x_19226;
wire x_19227;
wire x_19228;
wire x_19229;
wire x_19230;
wire x_19231;
wire x_19232;
wire x_19233;
wire x_19234;
wire x_19235;
wire x_19236;
wire x_19237;
wire x_19238;
wire x_19239;
wire x_19240;
wire x_19241;
wire x_19242;
wire x_19243;
wire x_19244;
wire x_19245;
wire x_19246;
wire x_19247;
wire x_19248;
wire x_19249;
wire x_19250;
wire x_19251;
wire x_19252;
wire x_19253;
wire x_19254;
wire x_19255;
wire x_19256;
wire x_19257;
wire x_19258;
wire x_19259;
wire x_19260;
wire x_19261;
wire x_19262;
wire x_19263;
wire x_19264;
wire x_19265;
wire x_19266;
wire x_19267;
wire x_19268;
wire x_19269;
wire x_19270;
wire x_19271;
wire x_19272;
wire x_19273;
wire x_19274;
wire x_19275;
wire x_19276;
wire x_19277;
wire x_19278;
wire x_19279;
wire x_19280;
wire x_19281;
wire x_19282;
wire x_19283;
wire x_19284;
wire x_19285;
wire x_19286;
wire x_19287;
wire x_19288;
wire x_19289;
wire x_19290;
wire x_19291;
wire x_19292;
wire x_19293;
wire x_19294;
wire x_19295;
wire x_19296;
wire x_19297;
wire x_19298;
wire x_19299;
wire x_19300;
wire x_19301;
wire x_19302;
wire x_19303;
wire x_19304;
wire x_19305;
wire x_19306;
wire x_19307;
wire x_19308;
wire x_19309;
wire x_19310;
wire x_19311;
wire x_19312;
wire x_19313;
wire x_19314;
wire x_19315;
wire x_19316;
wire x_19317;
wire x_19318;
wire x_19319;
wire x_19320;
wire x_19321;
wire x_19322;
wire x_19323;
wire x_19324;
wire x_19325;
wire x_19326;
wire x_19327;
wire x_19328;
wire x_19329;
wire x_19330;
wire x_19331;
wire x_19332;
wire x_19333;
wire x_19334;
wire x_19335;
wire x_19336;
wire x_19337;
wire x_19338;
wire x_19339;
wire x_19340;
wire x_19341;
wire x_19342;
wire x_19343;
wire x_19344;
wire x_19345;
wire x_19346;
wire x_19347;
wire x_19348;
wire x_19349;
wire x_19350;
wire x_19351;
wire x_19352;
wire x_19353;
wire x_19354;
wire x_19355;
wire x_19356;
wire x_19357;
wire x_19358;
wire x_19359;
wire x_19360;
wire x_19361;
wire x_19362;
wire x_19363;
wire x_19364;
wire x_19365;
wire x_19366;
wire x_19367;
wire x_19368;
wire x_19369;
wire x_19370;
wire x_19371;
wire x_19372;
wire x_19373;
wire x_19374;
wire x_19375;
wire x_19376;
wire x_19377;
wire x_19378;
wire x_19379;
wire x_19380;
wire x_19381;
wire x_19382;
wire x_19383;
wire x_19384;
wire x_19385;
wire x_19386;
wire x_19387;
wire x_19388;
wire x_19389;
wire x_19390;
wire x_19391;
wire x_19392;
wire x_19393;
wire x_19394;
wire x_19395;
wire x_19396;
wire x_19397;
wire x_19398;
wire x_19399;
wire x_19400;
wire x_19401;
wire x_19402;
wire x_19403;
wire x_19404;
wire x_19405;
wire x_19406;
wire x_19407;
wire x_19408;
wire x_19409;
wire x_19410;
wire x_19411;
wire x_19412;
wire x_19413;
wire x_19414;
wire x_19415;
wire x_19416;
wire x_19417;
wire x_19418;
wire x_19419;
wire x_19420;
wire x_19421;
wire x_19422;
wire x_19423;
wire x_19424;
wire x_19425;
wire x_19426;
wire x_19427;
wire x_19428;
wire x_19429;
wire x_19430;
wire x_19431;
wire x_19432;
wire x_19433;
wire x_19434;
wire x_19435;
wire x_19436;
wire x_19437;
wire x_19438;
wire x_19439;
wire x_19440;
wire x_19441;
wire x_19442;
wire x_19443;
wire x_19444;
wire x_19445;
wire x_19446;
wire x_19447;
wire x_19448;
wire x_19449;
wire x_19450;
wire x_19451;
wire x_19452;
wire x_19453;
wire x_19454;
wire x_19455;
wire x_19456;
wire x_19457;
wire x_19458;
wire x_19459;
wire x_19460;
wire x_19461;
wire x_19462;
wire x_19463;
wire x_19464;
wire x_19465;
wire x_19466;
wire x_19467;
wire x_19468;
wire x_19469;
wire x_19470;
wire x_19471;
wire x_19472;
wire x_19473;
wire x_19474;
wire x_19475;
wire x_19476;
wire x_19477;
wire x_19478;
wire x_19479;
wire x_19480;
wire x_19481;
wire x_19482;
wire x_19483;
wire x_19484;
wire x_19485;
wire x_19486;
wire x_19487;
wire x_19488;
wire x_19489;
wire x_19490;
wire x_19491;
wire x_19492;
wire x_19493;
wire x_19494;
wire x_19495;
wire x_19496;
wire x_19497;
wire x_19498;
wire x_19499;
wire x_19500;
wire x_19501;
wire x_19502;
wire x_19503;
wire x_19504;
wire x_19505;
wire x_19506;
wire x_19507;
wire x_19508;
wire x_19509;
wire x_19510;
wire x_19511;
wire x_19512;
wire x_19513;
wire x_19514;
wire x_19515;
wire x_19516;
wire x_19517;
wire x_19518;
wire x_19519;
wire x_19520;
wire x_19521;
wire x_19522;
wire x_19523;
wire x_19524;
wire x_19525;
wire x_19526;
wire x_19527;
wire x_19528;
wire x_19529;
wire x_19530;
wire x_19531;
wire x_19532;
wire x_19533;
wire x_19534;
wire x_19535;
wire x_19536;
wire x_19537;
wire x_19538;
wire x_19539;
wire x_19540;
wire x_19541;
wire x_19542;
wire x_19543;
wire x_19544;
wire x_19545;
wire x_19546;
wire x_19547;
wire x_19548;
wire x_19549;
wire x_19550;
wire x_19551;
wire x_19552;
wire x_19553;
wire x_19554;
wire x_19555;
wire x_19556;
wire x_19557;
wire x_19558;
wire x_19559;
wire x_19560;
wire x_19561;
wire x_19562;
wire x_19563;
wire x_19564;
wire x_19565;
wire x_19566;
wire x_19567;
wire x_19568;
wire x_19569;
wire x_19570;
wire x_19571;
wire x_19572;
wire x_19573;
wire x_19574;
wire x_19575;
wire x_19576;
wire x_19577;
wire x_19578;
wire x_19579;
wire x_19580;
wire x_19581;
wire x_19582;
wire x_19583;
wire x_19584;
wire x_19585;
wire x_19586;
wire x_19587;
wire x_19588;
wire x_19589;
wire x_19590;
wire x_19591;
wire x_19592;
wire x_19593;
wire x_19594;
wire x_19595;
wire x_19596;
wire x_19597;
wire x_19598;
wire x_19599;
wire x_19600;
wire x_19601;
wire x_19602;
wire x_19603;
wire x_19604;
wire x_19605;
wire x_19606;
wire x_19607;
wire x_19608;
wire x_19609;
wire x_19610;
wire x_19611;
wire x_19612;
wire x_19613;
wire x_19614;
wire x_19615;
wire x_19616;
wire x_19617;
wire x_19618;
wire x_19619;
wire x_19620;
wire x_19621;
wire x_19622;
wire x_19623;
wire x_19624;
wire x_19625;
wire x_19626;
wire x_19627;
wire x_19628;
wire x_19629;
wire x_19630;
wire x_19631;
wire x_19632;
wire x_19633;
wire x_19634;
wire x_19635;
wire x_19636;
wire x_19637;
wire x_19638;
wire x_19639;
wire x_19640;
wire x_19641;
wire x_19642;
wire x_19643;
wire x_19644;
wire x_19645;
wire x_19646;
wire x_19647;
wire x_19648;
wire x_19649;
wire x_19650;
wire x_19651;
wire x_19652;
wire x_19653;
wire x_19654;
wire x_19655;
wire x_19656;
wire x_19657;
wire x_19658;
wire x_19659;
wire x_19660;
wire x_19661;
wire x_19662;
wire x_19663;
wire x_19664;
wire x_19665;
wire x_19666;
wire x_19667;
wire x_19668;
wire x_19669;
wire x_19670;
wire x_19671;
wire x_19672;
wire x_19673;
wire x_19674;
wire x_19675;
wire x_19676;
wire x_19677;
wire x_19678;
wire x_19679;
wire x_19680;
wire x_19681;
wire x_19682;
wire x_19683;
wire x_19684;
wire x_19685;
wire x_19686;
wire x_19687;
wire x_19688;
wire x_19689;
wire x_19690;
wire x_19691;
wire x_19692;
wire x_19693;
wire x_19694;
wire x_19695;
wire x_19696;
wire x_19697;
wire x_19698;
wire x_19699;
wire x_19700;
wire x_19701;
wire x_19702;
wire x_19703;
wire x_19704;
wire x_19705;
wire x_19706;
wire x_19707;
wire x_19708;
wire x_19709;
wire x_19710;
wire x_19711;
wire x_19712;
wire x_19713;
wire x_19714;
wire x_19715;
wire x_19716;
wire x_19717;
wire x_19718;
wire x_19719;
wire x_19720;
wire x_19721;
wire x_19722;
wire x_19723;
wire x_19724;
wire x_19725;
wire x_19726;
wire x_19727;
wire x_19728;
wire x_19729;
wire x_19730;
wire x_19731;
wire x_19732;
wire x_19733;
wire x_19734;
wire x_19735;
wire x_19736;
wire x_19737;
wire x_19738;
wire x_19739;
wire x_19740;
wire x_19741;
wire x_19742;
wire x_19743;
wire x_19744;
wire x_19745;
wire x_19746;
wire x_19747;
wire x_19748;
wire x_19749;
wire x_19750;
wire x_19751;
wire x_19752;
wire x_19753;
wire x_19754;
wire x_19755;
wire x_19756;
wire x_19757;
wire x_19758;
wire x_19759;
wire x_19760;
wire x_19761;
wire x_19762;
wire x_19763;
wire x_19764;
wire x_19765;
wire x_19766;
wire x_19767;
wire x_19768;
wire x_19769;
wire x_19770;
wire x_19771;
wire x_19772;
wire x_19773;
wire x_19774;
wire x_19775;
wire x_19776;
wire x_19777;
wire x_19778;
wire x_19779;
wire x_19780;
wire x_19781;
wire x_19782;
wire x_19783;
wire x_19784;
wire x_19785;
wire x_19786;
wire x_19787;
wire x_19788;
wire x_19789;
wire x_19790;
wire x_19791;
wire x_19792;
wire x_19793;
wire x_19794;
wire x_19795;
wire x_19796;
wire x_19797;
wire x_19798;
wire x_19799;
wire x_19800;
wire x_19801;
wire x_19802;
wire x_19803;
wire x_19804;
wire x_19805;
wire x_19806;
wire x_19807;
wire x_19808;
wire x_19809;
wire x_19810;
wire x_19811;
wire x_19812;
wire x_19813;
wire x_19814;
wire x_19815;
wire x_19816;
wire x_19817;
wire x_19818;
wire x_19819;
wire x_19820;
wire x_19821;
wire x_19822;
wire x_19823;
wire x_19824;
wire x_19825;
wire x_19826;
wire x_19827;
wire x_19828;
wire x_19829;
wire x_19830;
wire x_19831;
wire x_19832;
wire x_19833;
wire x_19834;
wire x_19835;
wire x_19836;
wire x_19837;
wire x_19838;
wire x_19839;
wire x_19840;
wire x_19841;
wire x_19842;
wire x_19843;
wire x_19844;
wire x_19845;
wire x_19846;
wire x_19847;
wire x_19848;
wire x_19849;
wire x_19850;
wire x_19851;
wire x_19852;
wire x_19853;
wire x_19854;
wire x_19855;
wire x_19856;
wire x_19857;
wire x_19858;
wire x_19859;
wire x_19860;
wire x_19861;
wire x_19862;
wire x_19863;
wire x_19864;
wire x_19865;
wire x_19866;
wire x_19867;
wire x_19868;
wire x_19869;
wire x_19870;
wire x_19871;
wire x_19872;
wire x_19873;
wire x_19874;
wire x_19875;
wire x_19876;
wire x_19877;
wire x_19878;
wire x_19879;
wire x_19880;
wire x_19881;
wire x_19882;
wire x_19883;
wire x_19884;
wire x_19885;
wire x_19886;
wire x_19887;
wire x_19888;
wire x_19889;
wire x_19890;
wire x_19891;
wire x_19892;
wire x_19893;
wire x_19894;
wire x_19895;
wire x_19896;
wire x_19897;
wire x_19898;
wire x_19899;
wire x_19900;
wire x_19901;
wire x_19902;
wire x_19903;
wire x_19904;
wire x_19905;
wire x_19906;
wire x_19907;
wire x_19908;
wire x_19909;
wire x_19910;
wire x_19911;
wire x_19912;
wire x_19913;
wire x_19914;
wire x_19915;
wire x_19916;
wire x_19917;
wire x_19918;
wire x_19919;
wire x_19920;
wire x_19921;
wire x_19922;
wire x_19923;
wire x_19924;
wire x_19925;
wire x_19926;
wire x_19927;
wire x_19928;
wire x_19929;
wire x_19930;
wire x_19931;
wire x_19932;
wire x_19933;
wire x_19934;
wire x_19935;
wire x_19936;
wire x_19937;
wire x_19938;
wire x_19939;
wire x_19940;
wire x_19941;
wire x_19942;
wire x_19943;
wire x_19944;
wire x_19945;
wire x_19946;
wire x_19947;
wire x_19948;
wire x_19949;
wire x_19950;
wire x_19951;
wire x_19952;
wire x_19953;
wire x_19954;
wire x_19955;
wire x_19956;
wire x_19957;
wire x_19958;
wire x_19959;
wire x_19960;
wire x_19961;
wire x_19962;
wire x_19963;
wire x_19964;
wire x_19965;
wire x_19966;
wire x_19967;
wire x_19968;
wire x_19969;
wire x_19970;
wire x_19971;
wire x_19972;
wire x_19973;
wire x_19974;
wire x_19975;
wire x_19976;
wire x_19977;
wire x_19978;
wire x_19979;
wire x_19980;
wire x_19981;
wire x_19982;
wire x_19983;
wire x_19984;
wire x_19985;
wire x_19986;
wire x_19987;
wire x_19988;
wire x_19989;
wire x_19990;
wire x_19991;
wire x_19992;
wire x_19993;
wire x_19994;
wire x_19995;
wire x_19996;
wire x_19997;
wire x_19998;
wire x_19999;
wire x_20000;
wire x_20001;
wire x_20002;
wire x_20003;
wire x_20004;
wire x_20005;
wire x_20006;
wire x_20007;
wire x_20008;
wire x_20009;
wire x_20010;
wire x_20011;
wire x_20012;
wire x_20013;
wire x_20014;
wire x_20015;
wire x_20016;
wire x_20017;
wire x_20018;
wire x_20019;
wire x_20020;
wire x_20021;
wire x_20022;
wire x_20023;
wire x_20024;
wire x_20025;
wire x_20026;
wire x_20027;
wire x_20028;
wire x_20029;
wire x_20030;
wire x_20031;
wire x_20032;
wire x_20033;
wire x_20034;
wire x_20035;
wire x_20036;
wire x_20037;
wire x_20038;
wire x_20039;
wire x_20040;
wire x_20041;
wire x_20042;
wire x_20043;
wire x_20044;
wire x_20045;
wire x_20046;
wire x_20047;
wire x_20048;
wire x_20049;
wire x_20050;
wire x_20051;
wire x_20052;
wire x_20053;
wire x_20054;
wire x_20055;
wire x_20056;
wire x_20057;
wire x_20058;
wire x_20059;
wire x_20060;
wire x_20061;
wire x_20062;
wire x_20063;
wire x_20064;
wire x_20065;
wire x_20066;
wire x_20067;
wire x_20068;
wire x_20069;
wire x_20070;
wire x_20071;
wire x_20072;
wire x_20073;
wire x_20074;
wire x_20075;
wire x_20076;
wire x_20077;
wire x_20078;
wire x_20079;
wire x_20080;
wire x_20081;
wire x_20082;
wire x_20083;
wire x_20084;
wire x_20085;
wire x_20086;
wire x_20087;
wire x_20088;
wire x_20089;
wire x_20090;
wire x_20091;
wire x_20092;
wire x_20093;
wire x_20094;
wire x_20095;
wire x_20096;
wire x_20097;
wire x_20098;
wire x_20099;
wire x_20100;
wire x_20101;
wire x_20102;
wire x_20103;
wire x_20104;
wire x_20105;
wire x_20106;
wire x_20107;
wire x_20108;
wire x_20109;
wire x_20110;
wire x_20111;
wire x_20112;
wire x_20113;
wire x_20114;
wire x_20115;
wire x_20116;
wire x_20117;
wire x_20118;
wire x_20119;
wire x_20120;
wire x_20121;
wire x_20122;
wire x_20123;
wire x_20124;
wire x_20125;
wire x_20126;
wire x_20127;
wire x_20128;
wire x_20129;
wire x_20130;
wire x_20131;
wire x_20132;
wire x_20133;
wire x_20134;
wire x_20135;
wire x_20136;
wire x_20137;
wire x_20138;
wire x_20139;
wire x_20140;
wire x_20141;
wire x_20142;
wire x_20143;
wire x_20144;
wire x_20145;
wire x_20146;
wire x_20147;
wire x_20148;
wire x_20149;
wire x_20150;
wire x_20151;
wire x_20152;
wire x_20153;
wire x_20154;
wire x_20155;
wire x_20156;
wire x_20157;
wire x_20158;
wire x_20159;
wire x_20160;
wire x_20161;
wire x_20162;
wire x_20163;
wire x_20164;
wire x_20165;
wire x_20166;
wire x_20167;
wire x_20168;
wire x_20169;
wire x_20170;
wire x_20171;
wire x_20172;
wire x_20173;
wire x_20174;
wire x_20175;
wire x_20176;
wire x_20177;
wire x_20178;
wire x_20179;
wire x_20180;
wire x_20181;
wire x_20182;
wire x_20183;
wire x_20184;
wire x_20185;
wire x_20186;
wire x_20187;
wire x_20188;
wire x_20189;
wire x_20190;
wire x_20191;
wire x_20192;
wire x_20193;
wire x_20194;
wire x_20195;
wire x_20196;
wire x_20197;
wire x_20198;
wire x_20199;
wire x_20200;
wire x_20201;
wire x_20202;
wire x_20203;
wire x_20204;
wire x_20205;
wire x_20206;
wire x_20207;
wire x_20208;
wire x_20209;
wire x_20210;
wire x_20211;
wire x_20212;
wire x_20213;
wire x_20214;
wire x_20215;
wire x_20216;
wire x_20217;
wire x_20218;
wire x_20219;
wire x_20220;
wire x_20221;
wire x_20222;
wire x_20223;
wire x_20224;
wire x_20225;
wire x_20226;
wire x_20227;
wire x_20228;
wire x_20229;
wire x_20230;
wire x_20231;
wire x_20232;
wire x_20233;
wire x_20234;
wire x_20235;
wire x_20236;
wire x_20237;
wire x_20238;
wire x_20239;
wire x_20240;
wire x_20241;
wire x_20242;
wire x_20243;
wire x_20244;
wire x_20245;
wire x_20246;
wire x_20247;
wire x_20248;
wire x_20249;
wire x_20250;
wire x_20251;
wire x_20252;
wire x_20253;
wire x_20254;
wire x_20255;
wire x_20256;
wire x_20257;
wire x_20258;
wire x_20259;
wire x_20260;
wire x_20261;
wire x_20262;
wire x_20263;
wire x_20264;
wire x_20265;
wire x_20266;
wire x_20267;
wire x_20268;
wire x_20269;
wire x_20270;
wire x_20271;
wire x_20272;
wire x_20273;
wire x_20274;
wire x_20275;
wire x_20276;
wire x_20277;
wire x_20278;
wire x_20279;
wire x_20280;
wire x_20281;
wire x_20282;
wire x_20283;
wire x_20284;
wire x_20285;
wire x_20286;
wire x_20287;
wire x_20288;
wire x_20289;
wire x_20290;
wire x_20291;
wire x_20292;
wire x_20293;
wire x_20294;
wire x_20295;
wire x_20296;
wire x_20297;
wire x_20298;
wire x_20299;
wire x_20300;
wire x_20301;
wire x_20302;
wire x_20303;
wire x_20304;
wire x_20305;
wire x_20306;
wire x_20307;
wire x_20308;
wire x_20309;
wire x_20310;
wire x_20311;
wire x_20312;
wire x_20313;
wire x_20314;
wire x_20315;
wire x_20316;
wire x_20317;
wire x_20318;
wire x_20319;
wire x_20320;
wire x_20321;
wire x_20322;
wire x_20323;
wire x_20324;
wire x_20325;
wire x_20326;
wire x_20327;
wire x_20328;
wire x_20329;
wire x_20330;
wire x_20331;
wire x_20332;
wire x_20333;
wire x_20334;
wire x_20335;
wire x_20336;
wire x_20337;
wire x_20338;
wire x_20339;
wire x_20340;
wire x_20341;
wire x_20342;
wire x_20343;
wire x_20344;
wire x_20345;
wire x_20346;
wire x_20347;
wire x_20348;
wire x_20349;
wire x_20350;
wire x_20351;
wire x_20352;
wire x_20353;
wire x_20354;
wire x_20355;
wire x_20356;
wire x_20357;
wire x_20358;
wire x_20359;
wire x_20360;
wire x_20361;
wire x_20362;
wire x_20363;
wire x_20364;
wire x_20365;
wire x_20366;
wire x_20367;
wire x_20368;
wire x_20369;
wire x_20370;
wire x_20371;
wire x_20372;
wire x_20373;
wire x_20374;
wire x_20375;
wire x_20376;
wire x_20377;
wire x_20378;
wire x_20379;
wire x_20380;
wire x_20381;
wire x_20382;
wire x_20383;
wire x_20384;
wire x_20385;
wire x_20386;
wire x_20387;
wire x_20388;
wire x_20389;
wire x_20390;
wire x_20391;
wire x_20392;
wire x_20393;
wire x_20394;
wire x_20395;
wire x_20396;
wire x_20397;
wire x_20398;
wire x_20399;
wire x_20400;
wire x_20401;
wire x_20402;
wire x_20403;
wire x_20404;
wire x_20405;
wire x_20406;
wire x_20407;
wire x_20408;
wire x_20409;
wire x_20410;
wire x_20411;
wire x_20412;
wire x_20413;
wire x_20414;
wire x_20415;
wire x_20416;
wire x_20417;
wire x_20418;
wire x_20419;
wire x_20420;
wire x_20421;
wire x_20422;
wire x_20423;
wire x_20424;
wire x_20425;
wire x_20426;
wire x_20427;
wire x_20428;
wire x_20429;
wire x_20430;
wire x_20431;
wire x_20432;
wire x_20433;
wire x_20434;
wire x_20435;
wire x_20436;
wire x_20437;
wire x_20438;
wire x_20439;
wire x_20440;
wire x_20441;
wire x_20442;
wire x_20443;
wire x_20444;
wire x_20445;
wire x_20446;
wire x_20447;
wire x_20448;
wire x_20449;
wire x_20450;
wire x_20451;
wire x_20452;
wire x_20453;
wire x_20454;
wire x_20455;
wire x_20456;
wire x_20457;
wire x_20458;
wire x_20459;
wire x_20460;
wire x_20461;
wire x_20462;
wire x_20463;
wire x_20464;
wire x_20465;
wire x_20466;
wire x_20467;
wire x_20468;
wire x_20469;
wire x_20470;
wire x_20471;
wire x_20472;
wire x_20473;
wire x_20474;
wire x_20475;
wire x_20476;
wire x_20477;
wire x_20478;
wire x_20479;
wire x_20480;
wire x_20481;
wire x_20482;
wire x_20483;
wire x_20484;
wire x_20485;
wire x_20486;
wire x_20487;
wire x_20488;
wire x_20489;
wire x_20490;
wire x_20491;
wire x_20492;
wire x_20493;
wire x_20494;
wire x_20495;
wire x_20496;
wire x_20497;
wire x_20498;
wire x_20499;
wire x_20500;
wire x_20501;
wire x_20502;
wire x_20503;
wire x_20504;
wire x_20505;
wire x_20506;
wire x_20507;
wire x_20508;
wire x_20509;
wire x_20510;
wire x_20511;
wire x_20512;
wire x_20513;
wire x_20514;
wire x_20515;
wire x_20516;
wire x_20517;
wire x_20518;
wire x_20519;
wire x_20520;
wire x_20521;
wire x_20522;
wire x_20523;
wire x_20524;
wire x_20525;
wire x_20526;
wire x_20527;
wire x_20528;
wire x_20529;
wire x_20530;
wire x_20531;
wire x_20532;
wire x_20533;
wire x_20534;
wire x_20535;
wire x_20536;
wire x_20537;
wire x_20538;
wire x_20539;
wire x_20540;
wire x_20541;
wire x_20542;
wire x_20543;
wire x_20544;
wire x_20545;
wire x_20546;
wire x_20547;
wire x_20548;
wire x_20549;
wire x_20550;
wire x_20551;
wire x_20552;
wire x_20553;
wire x_20554;
wire x_20555;
wire x_20556;
wire x_20557;
wire x_20558;
wire x_20559;
wire x_20560;
wire x_20561;
wire x_20562;
wire x_20563;
wire x_20564;
wire x_20565;
wire x_20566;
wire x_20567;
wire x_20568;
wire x_20569;
wire x_20570;
wire x_20571;
wire x_20572;
wire x_20573;
wire x_20574;
wire x_20575;
wire x_20576;
wire x_20577;
wire x_20578;
wire x_20579;
wire x_20580;
wire x_20581;
wire x_20582;
wire x_20583;
wire x_20584;
wire x_20585;
wire x_20586;
wire x_20587;
wire x_20588;
wire x_20589;
wire x_20590;
wire x_20591;
wire x_20592;
wire x_20593;
wire x_20594;
wire x_20595;
wire x_20596;
wire x_20597;
wire x_20598;
wire x_20599;
wire x_20600;
wire x_20601;
wire x_20602;
wire x_20603;
wire x_20604;
wire x_20605;
wire x_20606;
wire x_20607;
wire x_20608;
wire x_20609;
wire x_20610;
wire x_20611;
wire x_20612;
wire x_20613;
wire x_20614;
wire x_20615;
wire x_20616;
wire x_20617;
wire x_20618;
wire x_20619;
wire x_20620;
wire x_20621;
wire x_20622;
wire x_20623;
wire x_20624;
wire x_20625;
wire x_20626;
wire x_20627;
wire x_20628;
wire x_20629;
wire x_20630;
wire x_20631;
wire x_20632;
wire x_20633;
wire x_20634;
wire x_20635;
wire x_20636;
wire x_20637;
wire x_20638;
wire x_20639;
wire x_20640;
wire x_20641;
wire x_20642;
wire x_20643;
wire x_20644;
wire x_20645;
wire x_20646;
wire x_20647;
wire x_20648;
wire x_20649;
wire x_20650;
wire x_20651;
wire x_20652;
wire x_20653;
wire x_20654;
wire x_20655;
wire x_20656;
wire x_20657;
wire x_20658;
wire x_20659;
wire x_20660;
wire x_20661;
wire x_20662;
wire x_20663;
wire x_20664;
wire x_20665;
wire x_20666;
wire x_20667;
wire x_20668;
wire x_20669;
wire x_20670;
wire x_20671;
wire x_20672;
wire x_20673;
wire x_20674;
wire x_20675;
wire x_20676;
wire x_20677;
wire x_20678;
wire x_20679;
wire x_20680;
wire x_20681;
wire x_20682;
wire x_20683;
wire x_20684;
wire x_20685;
wire x_20686;
wire x_20687;
wire x_20688;
wire x_20689;
wire x_20690;
wire x_20691;
wire x_20692;
wire x_20693;
wire x_20694;
wire x_20695;
wire x_20696;
wire x_20697;
wire x_20698;
wire x_20699;
wire x_20700;
wire x_20701;
wire x_20702;
wire x_20703;
wire x_20704;
wire x_20705;
wire x_20706;
wire x_20707;
wire x_20708;
wire x_20709;
wire x_20710;
wire x_20711;
wire x_20712;
wire x_20713;
wire x_20714;
wire x_20715;
wire x_20716;
wire x_20717;
wire x_20718;
wire x_20719;
wire x_20720;
wire x_20721;
wire x_20722;
wire x_20723;
wire x_20724;
wire x_20725;
wire x_20726;
wire x_20727;
wire x_20728;
wire x_20729;
wire x_20730;
wire x_20731;
wire x_20732;
wire x_20733;
wire x_20734;
wire x_20735;
wire x_20736;
wire x_20737;
wire x_20738;
wire x_20739;
wire x_20740;
wire x_20741;
wire x_20742;
wire x_20743;
wire x_20744;
wire x_20745;
wire x_20746;
wire x_20747;
wire x_20748;
wire x_20749;
wire x_20750;
wire x_20751;
wire x_20752;
wire x_20753;
wire x_20754;
wire x_20755;
wire x_20756;
wire x_20757;
wire x_20758;
wire x_20759;
wire x_20760;
wire x_20761;
wire x_20762;
wire x_20763;
wire x_20764;
wire x_20765;
wire x_20766;
wire x_20767;
wire x_20768;
wire x_20769;
wire x_20770;
wire x_20771;
wire x_20772;
wire x_20773;
wire x_20774;
wire x_20775;
wire x_20776;
wire x_20777;
wire x_20778;
wire x_20779;
wire x_20780;
wire x_20781;
wire x_20782;
wire x_20783;
wire x_20784;
wire x_20785;
wire x_20786;
wire x_20787;
wire x_20788;
wire x_20789;
wire x_20790;
wire x_20791;
wire x_20792;
wire x_20793;
wire x_20794;
wire x_20795;
wire x_20796;
wire x_20797;
wire x_20798;
wire x_20799;
wire x_20800;
wire x_20801;
wire x_20802;
wire x_20803;
wire x_20804;
wire x_20805;
wire x_20806;
wire x_20807;
wire x_20808;
wire x_20809;
wire x_20810;
wire x_20811;
wire x_20812;
wire x_20813;
wire x_20814;
wire x_20815;
wire x_20816;
wire x_20817;
wire x_20818;
wire x_20819;
wire x_20820;
wire x_20821;
wire x_20822;
wire x_20823;
wire x_20824;
wire x_20825;
wire x_20826;
wire x_20827;
wire x_20828;
wire x_20829;
wire x_20830;
wire x_20831;
wire x_20832;
wire x_20833;
wire x_20834;
wire x_20835;
wire x_20836;
wire x_20837;
wire x_20838;
wire x_20839;
wire x_20840;
wire x_20841;
wire x_20842;
wire x_20843;
wire x_20844;
wire x_20845;
wire x_20846;
wire x_20847;
wire x_20848;
wire x_20849;
wire x_20850;
wire x_20851;
wire x_20852;
wire x_20853;
wire x_20854;
wire x_20855;
wire x_20856;
wire x_20857;
wire x_20858;
wire x_20859;
wire x_20860;
wire x_20861;
wire x_20862;
wire x_20863;
wire x_20864;
wire x_20865;
wire x_20866;
wire x_20867;
wire x_20868;
wire x_20869;
wire x_20870;
wire x_20871;
wire x_20872;
wire x_20873;
wire x_20874;
wire x_20875;
wire x_20876;
wire x_20877;
wire x_20878;
wire x_20879;
wire x_20880;
wire x_20881;
wire x_20882;
wire x_20883;
wire x_20884;
wire x_20885;
wire x_20886;
wire x_20887;
wire x_20888;
wire x_20889;
wire x_20890;
wire x_20891;
wire x_20892;
wire x_20893;
wire x_20894;
wire x_20895;
wire x_20896;
wire x_20897;
wire x_20898;
wire x_20899;
wire x_20900;
wire x_20901;
wire x_20902;
wire x_20903;
wire x_20904;
wire x_20905;
wire x_20906;
wire x_20907;
wire x_20908;
wire x_20909;
wire x_20910;
wire x_20911;
wire x_20912;
wire x_20913;
wire x_20914;
wire x_20915;
wire x_20916;
wire x_20917;
wire x_20918;
wire x_20919;
wire x_20920;
wire x_20921;
wire x_20922;
wire x_20923;
wire x_20924;
wire x_20925;
wire x_20926;
wire x_20927;
wire x_20928;
wire x_20929;
wire x_20930;
wire x_20931;
wire x_20932;
wire x_20933;
wire x_20934;
wire x_20935;
wire x_20936;
wire x_20937;
wire x_20938;
wire x_20939;
wire x_20940;
wire x_20941;
wire x_20942;
wire x_20943;
wire x_20944;
wire x_20945;
wire x_20946;
wire x_20947;
wire x_20948;
wire x_20949;
wire x_20950;
wire x_20951;
wire x_20952;
wire x_20953;
wire x_20954;
wire x_20955;
wire x_20956;
wire x_20957;
wire x_20958;
wire x_20959;
wire x_20960;
wire x_20961;
wire x_20962;
wire x_20963;
wire x_20964;
wire x_20965;
wire x_20966;
wire x_20967;
wire x_20968;
wire x_20969;
wire x_20970;
wire x_20971;
wire x_20972;
wire x_20973;
wire x_20974;
wire x_20975;
wire x_20976;
wire x_20977;
wire x_20978;
wire x_20979;
wire x_20980;
wire x_20981;
wire x_20982;
wire x_20983;
wire x_20984;
wire x_20985;
wire x_20986;
wire x_20987;
wire x_20988;
wire x_20989;
wire x_20990;
wire x_20991;
wire x_20992;
wire x_20993;
wire x_20994;
wire x_20995;
wire x_20996;
wire x_20997;
wire x_20998;
wire x_20999;
wire x_21000;
wire x_21001;
wire x_21002;
wire x_21003;
wire x_21004;
wire x_21005;
wire x_21006;
wire x_21007;
wire x_21008;
wire x_21009;
wire x_21010;
wire x_21011;
wire x_21012;
wire x_21013;
wire x_21014;
wire x_21015;
wire x_21016;
wire x_21017;
wire x_21018;
wire x_21019;
wire x_21020;
wire x_21021;
wire x_21022;
wire x_21023;
wire x_21024;
wire x_21025;
wire x_21026;
wire x_21027;
wire x_21028;
wire x_21029;
wire x_21030;
wire x_21031;
wire x_21032;
wire x_21033;
wire x_21034;
wire x_21035;
wire x_21036;
wire x_21037;
wire x_21038;
wire x_21039;
wire x_21040;
wire x_21041;
wire x_21042;
wire x_21043;
wire x_21044;
wire x_21045;
wire x_21046;
wire x_21047;
wire x_21048;
wire x_21049;
wire x_21050;
wire x_21051;
wire x_21052;
wire x_21053;
wire x_21054;
wire x_21055;
wire x_21056;
wire x_21057;
wire x_21058;
wire x_21059;
wire x_21060;
wire x_21061;
wire x_21062;
wire x_21063;
wire x_21064;
wire x_21065;
wire x_21066;
wire x_21067;
wire x_21068;
wire x_21069;
wire x_21070;
wire x_21071;
wire x_21072;
wire x_21073;
wire x_21074;
wire x_21075;
wire x_21076;
wire x_21077;
wire x_21078;
wire x_21079;
wire x_21080;
wire x_21081;
wire x_21082;
wire x_21083;
wire x_21084;
wire x_21085;
wire x_21086;
wire x_21087;
wire x_21088;
wire x_21089;
wire x_21090;
wire x_21091;
wire x_21092;
wire x_21093;
wire x_21094;
wire x_21095;
wire x_21096;
wire x_21097;
wire x_21098;
wire x_21099;
wire x_21100;
wire x_21101;
wire x_21102;
wire x_21103;
wire x_21104;
wire x_21105;
wire x_21106;
wire x_21107;
wire x_21108;
wire x_21109;
wire x_21110;
wire x_21111;
wire x_21112;
wire x_21113;
wire x_21114;
wire x_21115;
wire x_21116;
wire x_21117;
wire x_21118;
wire x_21119;
wire x_21120;
wire x_21121;
wire x_21122;
wire x_21123;
wire x_21124;
wire x_21125;
wire x_21126;
wire x_21127;
wire x_21128;
wire x_21129;
wire x_21130;
wire x_21131;
wire x_21132;
wire x_21133;
wire x_21134;
wire x_21135;
wire x_21136;
wire x_21137;
wire x_21138;
wire x_21139;
wire x_21140;
wire x_21141;
wire x_21142;
wire x_21143;
wire x_21144;
wire x_21145;
wire x_21146;
wire x_21147;
wire x_21148;
wire x_21149;
wire x_21150;
wire x_21151;
wire x_21152;
wire x_21153;
wire x_21154;
wire x_21155;
wire x_21156;
wire x_21157;
wire x_21158;
wire x_21159;
wire x_21160;
wire x_21161;
wire x_21162;
wire x_21163;
wire x_21164;
wire x_21165;
wire x_21166;
wire x_21167;
wire x_21168;
wire x_21169;
wire x_21170;
wire x_21171;
wire x_21172;
wire x_21173;
wire x_21174;
wire x_21175;
wire x_21176;
wire x_21177;
wire x_21178;
wire x_21179;
wire x_21180;
wire x_21181;
wire x_21182;
wire x_21183;
wire x_21184;
wire x_21185;
wire x_21186;
wire x_21187;
wire x_21188;
wire x_21189;
wire x_21190;
wire x_21191;
wire x_21192;
wire x_21193;
wire x_21194;
wire x_21195;
wire x_21196;
wire x_21197;
wire x_21198;
wire x_21199;
wire x_21200;
wire x_21201;
wire x_21202;
wire x_21203;
wire x_21204;
wire x_21205;
wire x_21206;
wire x_21207;
wire x_21208;
wire x_21209;
wire x_21210;
wire x_21211;
wire x_21212;
wire x_21213;
wire x_21214;
wire x_21215;
wire x_21216;
wire x_21217;
wire x_21218;
wire x_21219;
wire x_21220;
wire x_21221;
wire x_21222;
wire x_21223;
wire x_21224;
wire x_21225;
wire x_21226;
wire x_21227;
wire x_21228;
wire x_21229;
wire x_21230;
wire x_21231;
wire x_21232;
wire x_21233;
wire x_21234;
wire x_21235;
wire x_21236;
wire x_21237;
wire x_21238;
wire x_21239;
wire x_21240;
wire x_21241;
wire x_21242;
wire x_21243;
wire x_21244;
wire x_21245;
wire x_21246;
wire x_21247;
wire x_21248;
wire x_21249;
wire x_21250;
wire x_21251;
wire x_21252;
wire x_21253;
wire x_21254;
wire x_21255;
wire x_21256;
wire x_21257;
wire x_21258;
wire x_21259;
wire x_21260;
wire x_21261;
wire x_21262;
wire x_21263;
wire x_21264;
wire x_21265;
wire x_21266;
wire x_21267;
wire x_21268;
wire x_21269;
wire x_21270;
wire x_21271;
wire x_21272;
wire x_21273;
wire x_21274;
wire x_21275;
wire x_21276;
wire x_21277;
wire x_21278;
wire x_21279;
wire x_21280;
wire x_21281;
wire x_21282;
wire x_21283;
wire x_21284;
wire x_21285;
wire x_21286;
wire x_21287;
wire x_21288;
wire x_21289;
wire x_21290;
wire x_21291;
wire x_21292;
wire x_21293;
wire x_21294;
wire x_21295;
wire x_21296;
wire x_21297;
wire x_21298;
wire x_21299;
wire x_21300;
wire x_21301;
wire x_21302;
wire x_21303;
wire x_21304;
wire x_21305;
wire x_21306;
wire x_21307;
wire x_21308;
wire x_21309;
wire x_21310;
wire x_21311;
wire x_21312;
wire x_21313;
wire x_21314;
wire x_21315;
wire x_21316;
wire x_21317;
wire x_21318;
wire x_21319;
wire x_21320;
wire x_21321;
wire x_21322;
wire x_21323;
wire x_21324;
wire x_21325;
wire x_21326;
wire x_21327;
wire x_21328;
wire x_21329;
wire x_21330;
wire x_21331;
wire x_21332;
wire x_21333;
wire x_21334;
wire x_21335;
wire x_21336;
wire x_21337;
wire x_21338;
wire x_21339;
wire x_21340;
wire x_21341;
wire x_21342;
wire x_21343;
wire x_21344;
wire x_21345;
wire x_21346;
wire x_21347;
wire x_21348;
wire x_21349;
wire x_21350;
wire x_21351;
wire x_21352;
wire x_21353;
wire x_21354;
wire x_21355;
wire x_21356;
wire x_21357;
wire x_21358;
wire x_21359;
wire x_21360;
wire x_21361;
wire x_21362;
wire x_21363;
wire x_21364;
wire x_21365;
wire x_21366;
wire x_21367;
wire x_21368;
wire x_21369;
wire x_21370;
wire x_21371;
wire x_21372;
wire x_21373;
wire x_21374;
wire x_21375;
wire x_21376;
wire x_21377;
wire x_21378;
wire x_21379;
wire x_21380;
wire x_21381;
wire x_21382;
wire x_21383;
wire x_21384;
wire x_21385;
wire x_21386;
wire x_21387;
wire x_21388;
wire x_21389;
wire x_21390;
wire x_21391;
wire x_21392;
wire x_21393;
wire x_21394;
wire x_21395;
wire x_21396;
wire x_21397;
wire x_21398;
wire x_21399;
wire x_21400;
wire x_21401;
wire x_21402;
wire x_21403;
wire x_21404;
wire x_21405;
wire x_21406;
wire x_21407;
wire x_21408;
wire x_21409;
wire x_21410;
wire x_21411;
wire x_21412;
wire x_21413;
wire x_21414;
wire x_21415;
wire x_21416;
wire x_21417;
wire x_21418;
wire x_21419;
wire x_21420;
wire x_21421;
wire x_21422;
wire x_21423;
wire x_21424;
wire x_21425;
wire x_21426;
wire x_21427;
wire x_21428;
wire x_21429;
wire x_21430;
wire x_21431;
wire x_21432;
wire x_21433;
wire x_21434;
wire x_21435;
wire x_21436;
wire x_21437;
wire x_21438;
wire x_21439;
wire x_21440;
wire x_21441;
wire x_21442;
wire x_21443;
wire x_21444;
wire x_21445;
wire x_21446;
wire x_21447;
wire x_21448;
wire x_21449;
wire x_21450;
wire x_21451;
wire x_21452;
wire x_21453;
wire x_21454;
wire x_21455;
wire x_21456;
wire x_21457;
wire x_21458;
wire x_21459;
wire x_21460;
wire x_21461;
wire x_21462;
wire x_21463;
wire x_21464;
wire x_21465;
wire x_21466;
wire x_21467;
wire x_21468;
wire x_21469;
wire x_21470;
wire x_21471;
wire x_21472;
wire x_21473;
wire x_21474;
wire x_21475;
wire x_21476;
wire x_21477;
wire x_21478;
wire x_21479;
wire x_21480;
wire x_21481;
wire x_21482;
wire x_21483;
wire x_21484;
wire x_21485;
wire x_21486;
wire x_21487;
wire x_21488;
wire x_21489;
wire x_21490;
wire x_21491;
wire x_21492;
wire x_21493;
wire x_21494;
wire x_21495;
wire x_21496;
wire x_21497;
wire x_21498;
wire x_21499;
wire x_21500;
wire x_21501;
wire x_21502;
wire x_21503;
wire x_21504;
wire x_21505;
wire x_21506;
wire x_21507;
wire x_21508;
wire x_21509;
wire x_21510;
wire x_21511;
wire x_21512;
wire x_21513;
wire x_21514;
wire x_21515;
wire x_21516;
wire x_21517;
wire x_21518;
wire x_21519;
wire x_21520;
wire x_21521;
wire x_21522;
wire x_21523;
wire x_21524;
wire x_21525;
wire x_21526;
wire x_21527;
wire x_21528;
wire x_21529;
wire x_21530;
wire x_21531;
wire x_21532;
wire x_21533;
wire x_21534;
wire x_21535;
wire x_21536;
wire x_21537;
wire x_21538;
wire x_21539;
wire x_21540;
wire x_21541;
wire x_21542;
wire x_21543;
wire x_21544;
wire x_21545;
wire x_21546;
wire x_21547;
wire x_21548;
wire x_21549;
wire x_21550;
wire x_21551;
wire x_21552;
wire x_21553;
wire x_21554;
wire x_21555;
wire x_21556;
wire x_21557;
wire x_21558;
wire x_21559;
wire x_21560;
wire x_21561;
wire x_21562;
wire x_21563;
wire x_21564;
wire x_21565;
wire x_21566;
wire x_21567;
wire x_21568;
wire x_21569;
wire x_21570;
wire x_21571;
wire x_21572;
wire x_21573;
wire x_21574;
wire x_21575;
wire x_21576;
wire x_21577;
wire x_21578;
wire x_21579;
wire x_21580;
wire x_21581;
wire x_21582;
wire x_21583;
wire x_21584;
wire x_21585;
wire x_21586;
wire x_21587;
wire x_21588;
wire x_21589;
wire x_21590;
wire x_21591;
wire x_21592;
wire x_21593;
wire x_21594;
wire x_21595;
wire x_21596;
wire x_21597;
wire x_21598;
wire x_21599;
wire x_21600;
wire x_21601;
wire x_21602;
wire x_21603;
wire x_21604;
wire x_21605;
wire x_21606;
wire x_21607;
wire x_21608;
wire x_21609;
wire x_21610;
wire x_21611;
wire x_21612;
wire x_21613;
wire x_21614;
wire x_21615;
wire x_21616;
wire x_21617;
wire x_21618;
wire x_21619;
wire x_21620;
wire x_21621;
wire x_21622;
wire x_21623;
wire x_21624;
wire x_21625;
wire x_21626;
wire x_21627;
wire x_21628;
wire x_21629;
wire x_21630;
wire x_21631;
wire x_21632;
wire x_21633;
wire x_21634;
wire x_21635;
wire x_21636;
wire x_21637;
wire x_21638;
wire x_21639;
wire x_21640;
wire x_21641;
wire x_21642;
wire x_21643;
wire x_21644;
wire x_21645;
wire x_21646;
wire x_21647;
wire x_21648;
wire x_21649;
wire x_21650;
wire x_21651;
wire x_21652;
wire x_21653;
wire x_21654;
wire x_21655;
wire x_21656;
wire x_21657;
wire x_21658;
wire x_21659;
wire x_21660;
wire x_21661;
wire x_21662;
wire x_21663;
wire x_21664;
wire x_21665;
wire x_21666;
wire x_21667;
wire x_21668;
wire x_21669;
wire x_21670;
wire x_21671;
wire x_21672;
wire x_21673;
wire x_21674;
wire x_21675;
wire x_21676;
wire x_21677;
wire x_21678;
wire x_21679;
wire x_21680;
wire x_21681;
wire x_21682;
wire x_21683;
wire x_21684;
wire x_21685;
wire x_21686;
wire x_21687;
wire x_21688;
wire x_21689;
wire x_21690;
wire x_21691;
wire x_21692;
wire x_21693;
wire x_21694;
wire x_21695;
wire x_21696;
wire x_21697;
wire x_21698;
wire x_21699;
wire x_21700;
wire x_21701;
wire x_21702;
wire x_21703;
wire x_21704;
wire x_21705;
wire x_21706;
wire x_21707;
wire x_21708;
wire x_21709;
wire x_21710;
wire x_21711;
wire x_21712;
wire x_21713;
wire x_21714;
wire x_21715;
wire x_21716;
wire x_21717;
wire x_21718;
wire x_21719;
wire x_21720;
wire x_21721;
wire x_21722;
wire x_21723;
wire x_21724;
wire x_21725;
wire x_21726;
wire x_21727;
wire x_21728;
wire x_21729;
wire x_21730;
wire x_21731;
wire x_21732;
wire x_21733;
wire x_21734;
wire x_21735;
wire x_21736;
wire x_21737;
wire x_21738;
wire x_21739;
wire x_21740;
wire x_21741;
wire x_21742;
wire x_21743;
wire x_21744;
wire x_21745;
wire x_21746;
wire x_21747;
wire x_21748;
wire x_21749;
wire x_21750;
wire x_21751;
wire x_21752;
wire x_21753;
wire x_21754;
wire x_21755;
wire x_21756;
wire x_21757;
wire x_21758;
wire x_21759;
wire x_21760;
wire x_21761;
wire x_21762;
wire x_21763;
wire x_21764;
wire x_21765;
wire x_21766;
wire x_21767;
wire x_21768;
wire x_21769;
wire x_21770;
wire x_21771;
wire x_21772;
wire x_21773;
wire x_21774;
wire x_21775;
wire x_21776;
wire x_21777;
wire x_21778;
wire x_21779;
wire x_21780;
wire x_21781;
wire x_21782;
wire x_21783;
wire x_21784;
wire x_21785;
wire x_21786;
wire x_21787;
wire x_21788;
wire x_21789;
wire x_21790;
wire x_21791;
wire x_21792;
wire x_21793;
wire x_21794;
wire x_21795;
wire x_21796;
wire x_21797;
wire x_21798;
wire x_21799;
wire x_21800;
wire x_21801;
wire x_21802;
wire x_21803;
wire x_21804;
wire x_21805;
wire x_21806;
wire x_21807;
wire x_21808;
wire x_21809;
wire x_21810;
wire x_21811;
wire x_21812;
wire x_21813;
wire x_21814;
wire x_21815;
wire x_21816;
wire x_21817;
wire x_21818;
wire x_21819;
wire x_21820;
wire x_21821;
wire x_21822;
wire x_21823;
wire x_21824;
wire x_21825;
wire x_21826;
wire x_21827;
wire x_21828;
wire x_21829;
wire x_21830;
wire x_21831;
wire x_21832;
wire x_21833;
wire x_21834;
wire x_21835;
wire x_21836;
wire x_21837;
wire x_21838;
wire x_21839;
wire x_21840;
wire x_21841;
wire x_21842;
wire x_21843;
wire x_21844;
wire x_21845;
wire x_21846;
wire x_21847;
wire x_21848;
wire x_21849;
wire x_21850;
wire x_21851;
wire x_21852;
wire x_21853;
wire x_21854;
wire x_21855;
wire x_21856;
wire x_21857;
wire x_21858;
wire x_21859;
wire x_21860;
wire x_21861;
wire x_21862;
wire x_21863;
wire x_21864;
wire x_21865;
wire x_21866;
wire x_21867;
wire x_21868;
wire x_21869;
wire x_21870;
wire x_21871;
wire x_21872;
wire x_21873;
wire x_21874;
wire x_21875;
wire x_21876;
wire x_21877;
wire x_21878;
wire x_21879;
wire x_21880;
wire x_21881;
wire x_21882;
wire x_21883;
wire x_21884;
wire x_21885;
wire x_21886;
wire x_21887;
wire x_21888;
wire x_21889;
wire x_21890;
wire x_21891;
wire x_21892;
wire x_21893;
wire x_21894;
wire x_21895;
wire x_21896;
wire x_21897;
wire x_21898;
wire x_21899;
wire x_21900;
wire x_21901;
wire x_21902;
wire x_21903;
wire x_21904;
wire x_21905;
wire x_21906;
wire x_21907;
wire x_21908;
wire x_21909;
wire x_21910;
wire x_21911;
wire x_21912;
wire x_21913;
wire x_21914;
wire x_21915;
wire x_21916;
wire x_21917;
wire x_21918;
wire x_21919;
wire x_21920;
wire x_21921;
wire x_21922;
wire x_21923;
wire x_21924;
wire x_21925;
wire x_21926;
wire x_21927;
wire x_21928;
wire x_21929;
wire x_21930;
wire x_21931;
wire x_21932;
wire x_21933;
wire x_21934;
wire x_21935;
wire x_21936;
wire x_21937;
wire x_21938;
wire x_21939;
wire x_21940;
wire x_21941;
wire x_21942;
wire x_21943;
wire x_21944;
wire x_21945;
wire x_21946;
wire x_21947;
wire x_21948;
wire x_21949;
wire x_21950;
wire x_21951;
wire x_21952;
wire x_21953;
wire x_21954;
wire x_21955;
wire x_21956;
wire x_21957;
wire x_21958;
wire x_21959;
wire x_21960;
wire x_21961;
wire x_21962;
wire x_21963;
wire x_21964;
wire x_21965;
wire x_21966;
wire x_21967;
wire x_21968;
wire x_21969;
wire x_21970;
wire x_21971;
wire x_21972;
wire x_21973;
wire x_21974;
wire x_21975;
wire x_21976;
wire x_21977;
wire x_21978;
wire x_21979;
wire x_21980;
wire x_21981;
wire x_21982;
wire x_21983;
wire x_21984;
wire x_21985;
wire x_21986;
wire x_21987;
wire x_21988;
wire x_21989;
wire x_21990;
wire x_21991;
wire x_21992;
wire x_21993;
wire x_21994;
wire x_21995;
wire x_21996;
wire x_21997;
wire x_21998;
wire x_21999;
wire x_22000;
wire x_22001;
wire x_22002;
wire x_22003;
wire x_22004;
wire x_22005;
wire x_22006;
wire x_22007;
wire x_22008;
wire x_22009;
wire x_22010;
wire x_22011;
wire x_22012;
wire x_22013;
wire x_22014;
wire x_22015;
wire x_22016;
wire x_22017;
wire x_22018;
wire x_22019;
wire x_22020;
wire x_22021;
wire x_22022;
wire x_22023;
wire x_22024;
wire x_22025;
wire x_22026;
wire x_22027;
wire x_22028;
wire x_22029;
wire x_22030;
wire x_22031;
wire x_22032;
wire x_22033;
wire x_22034;
wire x_22035;
wire x_22036;
wire x_22037;
wire x_22038;
wire x_22039;
wire x_22040;
wire x_22041;
wire x_22042;
wire x_22043;
wire x_22044;
wire x_22045;
wire x_22046;
wire x_22047;
wire x_22048;
wire x_22049;
wire x_22050;
wire x_22051;
wire x_22052;
wire x_22053;
wire x_22054;
wire x_22055;
wire x_22056;
wire x_22057;
wire x_22058;
wire x_22059;
wire x_22060;
wire x_22061;
wire x_22062;
wire x_22063;
wire x_22064;
wire x_22065;
wire x_22066;
wire x_22067;
wire x_22068;
wire x_22069;
wire x_22070;
wire x_22071;
wire x_22072;
wire x_22073;
wire x_22074;
wire x_22075;
wire x_22076;
wire x_22077;
wire x_22078;
wire x_22079;
wire x_22080;
wire x_22081;
wire x_22082;
wire x_22083;
wire x_22084;
wire x_22085;
wire x_22086;
wire x_22087;
wire x_22088;
wire x_22089;
wire x_22090;
wire x_22091;
wire x_22092;
wire x_22093;
wire x_22094;
wire x_22095;
wire x_22096;
wire x_22097;
wire x_22098;
wire x_22099;
wire x_22100;
wire x_22101;
wire x_22102;
wire x_22103;
wire x_22104;
wire x_22105;
wire x_22106;
wire x_22107;
wire x_22108;
wire x_22109;
wire x_22110;
wire x_22111;
wire x_22112;
wire x_22113;
wire x_22114;
wire x_22115;
wire x_22116;
wire x_22117;
wire x_22118;
wire x_22119;
wire x_22120;
wire x_22121;
wire x_22122;
wire x_22123;
wire x_22124;
wire x_22125;
wire x_22126;
wire x_22127;
wire x_22128;
wire x_22129;
wire x_22130;
wire x_22131;
wire x_22132;
wire x_22133;
wire x_22134;
wire x_22135;
wire x_22136;
wire x_22137;
wire x_22138;
wire x_22139;
wire x_22140;
wire x_22141;
wire x_22142;
wire x_22143;
wire x_22144;
wire x_22145;
wire x_22146;
wire x_22147;
wire x_22148;
wire x_22149;
wire x_22150;
wire x_22151;
wire x_22152;
wire x_22153;
wire x_22154;
wire x_22155;
wire x_22156;
wire x_22157;
wire x_22158;
wire x_22159;
wire x_22160;
wire x_22161;
wire x_22162;
wire x_22163;
wire x_22164;
wire x_22165;
wire x_22166;
wire x_22167;
wire x_22168;
wire x_22169;
wire x_22170;
wire x_22171;
wire x_22172;
wire x_22173;
wire x_22174;
wire x_22175;
wire x_22176;
wire x_22177;
wire x_22178;
wire x_22179;
wire x_22180;
wire x_22181;
wire x_22182;
wire x_22183;
wire x_22184;
wire x_22185;
wire x_22186;
wire x_22187;
wire x_22188;
wire x_22189;
wire x_22190;
wire x_22191;
wire x_22192;
wire x_22193;
wire x_22194;
wire x_22195;
wire x_22196;
wire x_22197;
wire x_22198;
wire x_22199;
wire x_22200;
wire x_22201;
wire x_22202;
wire x_22203;
wire x_22204;
wire x_22205;
wire x_22206;
wire x_22207;
wire x_22208;
wire x_22209;
wire x_22210;
wire x_22211;
wire x_22212;
wire x_22213;
wire x_22214;
wire x_22215;
wire x_22216;
wire x_22217;
wire x_22218;
wire x_22219;
wire x_22220;
wire x_22221;
wire x_22222;
wire x_22223;
wire x_22224;
wire x_22225;
wire x_22226;
wire x_22227;
wire x_22228;
wire x_22229;
wire x_22230;
wire x_22231;
wire x_22232;
wire x_22233;
wire x_22234;
wire x_22235;
wire x_22236;
wire x_22237;
wire x_22238;
wire x_22239;
wire x_22240;
wire x_22241;
wire x_22242;
wire x_22243;
wire x_22244;
wire x_22245;
wire x_22246;
wire x_22247;
wire x_22248;
wire x_22249;
wire x_22250;
wire x_22251;
wire x_22252;
wire x_22253;
wire x_22254;
wire x_22255;
wire x_22256;
wire x_22257;
wire x_22258;
wire x_22259;
wire x_22260;
wire x_22261;
wire x_22262;
wire x_22263;
wire x_22264;
wire x_22265;
wire x_22266;
wire x_22267;
wire x_22268;
wire x_22269;
wire x_22270;
wire x_22271;
wire x_22272;
wire x_22273;
wire x_22274;
wire x_22275;
wire x_22276;
wire x_22277;
wire x_22278;
wire x_22279;
wire x_22280;
wire x_22281;
wire x_22282;
wire x_22283;
wire x_22284;
wire x_22285;
wire x_22286;
wire x_22287;
wire x_22288;
wire x_22289;
wire x_22290;
wire x_22291;
wire x_22292;
wire x_22293;
wire x_22294;
wire x_22295;
wire x_22296;
wire x_22297;
wire x_22298;
wire x_22299;
wire x_22300;
wire x_22301;
wire x_22302;
wire x_22303;
wire x_22304;
wire x_22305;
wire x_22306;
wire x_22307;
wire x_22308;
wire x_22309;
wire x_22310;
wire x_22311;
wire x_22312;
wire x_22313;
wire x_22314;
wire x_22315;
wire x_22316;
wire x_22317;
wire x_22318;
wire x_22319;
wire x_22320;
wire x_22321;
wire x_22322;
wire x_22323;
wire x_22324;
wire x_22325;
wire x_22326;
wire x_22327;
wire x_22328;
wire x_22329;
wire x_22330;
wire x_22331;
wire x_22332;
wire x_22333;
wire x_22334;
wire x_22335;
wire x_22336;
wire x_22337;
wire x_22338;
wire x_22339;
wire x_22340;
wire x_22341;
wire x_22342;
wire x_22343;
wire x_22344;
wire x_22345;
wire x_22346;
wire x_22347;
wire x_22348;
wire x_22349;
wire x_22350;
wire x_22351;
wire x_22352;
wire x_22353;
wire x_22354;
wire x_22355;
wire x_22356;
wire x_22357;
wire x_22358;
wire x_22359;
wire x_22360;
wire x_22361;
wire x_22362;
wire x_22363;
wire x_22364;
wire x_22365;
wire x_22366;
wire x_22367;
wire x_22368;
wire x_22369;
wire x_22370;
wire x_22371;
wire x_22372;
wire x_22373;
wire x_22374;
wire x_22375;
wire x_22376;
wire x_22377;
wire x_22378;
wire x_22379;
wire x_22380;
wire x_22381;
wire x_22382;
wire x_22383;
wire x_22384;
wire x_22385;
wire x_22386;
wire x_22387;
wire x_22388;
wire x_22389;
wire x_22390;
wire x_22391;
wire x_22392;
wire x_22393;
wire x_22394;
wire x_22395;
wire x_22396;
wire x_22397;
wire x_22398;
wire x_22399;
wire x_22400;
wire x_22401;
wire x_22402;
wire x_22403;
wire x_22404;
wire x_22405;
wire x_22406;
wire x_22407;
wire x_22408;
wire x_22409;
wire x_22410;
wire x_22411;
wire x_22412;
wire x_22413;
wire x_22414;
wire x_22415;
wire x_22416;
wire x_22417;
wire x_22418;
wire x_22419;
wire x_22420;
wire x_22421;
wire x_22422;
wire x_22423;
wire x_22424;
wire x_22425;
wire x_22426;
wire x_22427;
wire x_22428;
wire x_22429;
wire x_22430;
wire x_22431;
wire x_22432;
wire x_22433;
wire x_22434;
wire x_22435;
wire x_22436;
wire x_22437;
wire x_22438;
wire x_22439;
wire x_22440;
wire x_22441;
wire x_22442;
wire x_22443;
wire x_22444;
wire x_22445;
wire x_22446;
wire x_22447;
wire x_22448;
wire x_22449;
wire x_22450;
wire x_22451;
wire x_22452;
wire x_22453;
wire x_22454;
wire x_22455;
wire x_22456;
wire x_22457;
wire x_22458;
wire x_22459;
wire x_22460;
wire x_22461;
wire x_22462;
wire x_22463;
wire x_22464;
wire x_22465;
wire x_22466;
wire x_22467;
wire x_22468;
wire x_22469;
wire x_22470;
wire x_22471;
wire x_22472;
wire x_22473;
wire x_22474;
wire x_22475;
wire x_22476;
wire x_22477;
wire x_22478;
wire x_22479;
wire x_22480;
wire x_22481;
wire x_22482;
wire x_22483;
wire x_22484;
wire x_22485;
wire x_22486;
wire x_22487;
wire x_22488;
wire x_22489;
wire x_22490;
wire x_22491;
wire x_22492;
wire x_22493;
wire x_22494;
wire x_22495;
wire x_22496;
wire x_22497;
wire x_22498;
wire x_22499;
wire x_22500;
wire x_22501;
wire x_22502;
wire x_22503;
wire x_22504;
wire x_22505;
wire x_22506;
wire x_22507;
wire x_22508;
wire x_22509;
wire x_22510;
wire x_22511;
wire x_22512;
wire x_22513;
wire x_22514;
wire x_22515;
wire x_22516;
wire x_22517;
wire x_22518;
wire x_22519;
wire x_22520;
wire x_22521;
wire x_22522;
wire x_22523;
wire x_22524;
wire x_22525;
wire x_22526;
wire x_22527;
wire x_22528;
wire x_22529;
wire x_22530;
wire x_22531;
wire x_22532;
wire x_22533;
wire x_22534;
wire x_22535;
wire x_22536;
wire x_22537;
wire x_22538;
wire x_22539;
wire x_22540;
wire x_22541;
wire x_22542;
wire x_22543;
wire x_22544;
wire x_22545;
wire x_22546;
wire x_22547;
wire x_22548;
wire x_22549;
wire x_22550;
wire x_22551;
wire x_22552;
wire x_22553;
wire x_22554;
wire x_22555;
wire x_22556;
wire x_22557;
wire x_22558;
wire x_22559;
wire x_22560;
wire x_22561;
wire x_22562;
wire x_22563;
wire x_22564;
wire x_22565;
wire x_22566;
wire x_22567;
wire x_22568;
wire x_22569;
wire x_22570;
wire x_22571;
wire x_22572;
wire x_22573;
wire x_22574;
wire x_22575;
wire x_22576;
wire x_22577;
wire x_22578;
wire x_22579;
wire x_22580;
wire x_22581;
wire x_22582;
wire x_22583;
wire x_22584;
wire x_22585;
wire x_22586;
wire x_22587;
wire x_22588;
wire x_22589;
wire x_22590;
wire x_22591;
wire x_22592;
wire x_22593;
wire x_22594;
wire x_22595;
wire x_22596;
wire x_22597;
wire x_22598;
wire x_22599;
wire x_22600;
wire x_22601;
wire x_22602;
wire x_22603;
wire x_22604;
wire x_22605;
wire x_22606;
wire x_22607;
wire x_22608;
wire x_22609;
wire x_22610;
wire x_22611;
wire x_22612;
wire x_22613;
wire x_22614;
wire x_22615;
wire x_22616;
wire x_22617;
wire x_22618;
wire x_22619;
wire x_22620;
wire x_22621;
wire x_22622;
wire x_22623;
wire x_22624;
wire x_22625;
wire x_22626;
wire x_22627;
wire x_22628;
wire x_22629;
wire x_22630;
wire x_22631;
wire x_22632;
wire x_22633;
wire x_22634;
wire x_22635;
wire x_22636;
wire x_22637;
wire x_22638;
wire x_22639;
wire x_22640;
wire x_22641;
wire x_22642;
wire x_22643;
wire x_22644;
wire x_22645;
wire x_22646;
wire x_22647;
wire x_22648;
wire x_22649;
wire x_22650;
wire x_22651;
wire x_22652;
wire x_22653;
wire x_22654;
wire x_22655;
wire x_22656;
wire x_22657;
wire x_22658;
wire x_22659;
wire x_22660;
wire x_22661;
wire x_22662;
wire x_22663;
wire x_22664;
wire x_22665;
wire x_22666;
wire x_22667;
wire x_22668;
wire x_22669;
wire x_22670;
wire x_22671;
wire x_22672;
wire x_22673;
wire x_22674;
wire x_22675;
wire x_22676;
wire x_22677;
wire x_22678;
wire x_22679;
wire x_22680;
wire x_22681;
wire x_22682;
wire x_22683;
wire x_22684;
wire x_22685;
wire x_22686;
wire x_22687;
wire x_22688;
wire x_22689;
wire x_22690;
wire x_22691;
wire x_22692;
wire x_22693;
wire x_22694;
wire x_22695;
wire x_22696;
wire x_22697;
wire x_22698;
wire x_22699;
wire x_22700;
wire x_22701;
wire x_22702;
wire x_22703;
wire x_22704;
wire x_22705;
wire x_22706;
wire x_22707;
wire x_22708;
wire x_22709;
wire x_22710;
wire x_22711;
wire x_22712;
wire x_22713;
wire x_22714;
wire x_22715;
wire x_22716;
wire x_22717;
wire x_22718;
wire x_22719;
wire x_22720;
wire x_22721;
wire x_22722;
wire x_22723;
wire x_22724;
wire x_22725;
wire x_22726;
wire x_22727;
wire x_22728;
wire x_22729;
wire x_22730;
wire x_22731;
wire x_22732;
wire x_22733;
wire x_22734;
wire x_22735;
wire x_22736;
wire x_22737;
wire x_22738;
wire x_22739;
wire x_22740;
wire x_22741;
wire x_22742;
wire x_22743;
wire x_22744;
wire x_22745;
wire x_22746;
wire x_22747;
wire x_22748;
wire x_22749;
wire x_22750;
wire x_22751;
wire x_22752;
wire x_22753;
wire x_22754;
wire x_22755;
wire x_22756;
wire x_22757;
wire x_22758;
wire x_22759;
wire x_22760;
wire x_22761;
wire x_22762;
wire x_22763;
wire x_22764;
wire x_22765;
wire x_22766;
wire x_22767;
wire x_22768;
wire x_22769;
wire x_22770;
wire x_22771;
wire x_22772;
wire x_22773;
wire x_22774;
wire x_22775;
wire x_22776;
wire x_22777;
wire x_22778;
wire x_22779;
wire x_22780;
wire x_22781;
wire x_22782;
wire x_22783;
wire x_22784;
wire x_22785;
wire x_22786;
wire x_22787;
wire x_22788;
wire x_22789;
wire x_22790;
wire x_22791;
wire x_22792;
wire x_22793;
wire x_22794;
wire x_22795;
wire x_22796;
wire x_22797;
wire x_22798;
wire x_22799;
wire x_22800;
wire x_22801;
wire x_22802;
wire x_22803;
wire x_22804;
wire x_22805;
wire x_22806;
wire x_22807;
wire x_22808;
wire x_22809;
wire x_22810;
wire x_22811;
wire x_22812;
wire x_22813;
wire x_22814;
wire x_22815;
wire x_22816;
wire x_22817;
wire x_22818;
wire x_22819;
wire x_22820;
wire x_22821;
wire x_22822;
wire x_22823;
wire x_22824;
wire x_22825;
wire x_22826;
wire x_22827;
wire x_22828;
wire x_22829;
wire x_22830;
wire x_22831;
wire x_22832;
wire x_22833;
wire x_22834;
wire x_22835;
wire x_22836;
wire x_22837;
wire x_22838;
wire x_22839;
wire x_22840;
wire x_22841;
wire x_22842;
wire x_22843;
wire x_22844;
wire x_22845;
wire x_22846;
wire x_22847;
wire x_22848;
wire x_22849;
wire x_22850;
wire x_22851;
wire x_22852;
wire x_22853;
wire x_22854;
wire x_22855;
wire x_22856;
wire x_22857;
wire x_22858;
wire x_22859;
wire x_22860;
wire x_22861;
wire x_22862;
wire x_22863;
wire x_22864;
wire x_22865;
wire x_22866;
wire x_22867;
wire x_22868;
wire x_22869;
wire x_22870;
wire x_22871;
wire x_22872;
wire x_22873;
wire x_22874;
wire x_22875;
wire x_22876;
wire x_22877;
wire x_22878;
wire x_22879;
wire x_22880;
wire x_22881;
wire x_22882;
wire x_22883;
wire x_22884;
wire x_22885;
wire x_22886;
wire x_22887;
wire x_22888;
wire x_22889;
wire x_22890;
wire x_22891;
wire x_22892;
wire x_22893;
wire x_22894;
wire x_22895;
wire x_22896;
wire x_22897;
wire x_22898;
wire x_22899;
wire x_22900;
wire x_22901;
wire x_22902;
wire x_22903;
wire x_22904;
wire x_22905;
wire x_22906;
wire x_22907;
wire x_22908;
wire x_22909;
wire x_22910;
wire x_22911;
wire x_22912;
wire x_22913;
wire x_22914;
wire x_22915;
wire x_22916;
wire x_22917;
wire x_22918;
wire x_22919;
wire x_22920;
wire x_22921;
wire x_22922;
wire x_22923;
wire x_22924;
wire x_22925;
wire x_22926;
wire x_22927;
wire x_22928;
wire x_22929;
wire x_22930;
wire x_22931;
wire x_22932;
wire x_22933;
wire x_22934;
wire x_22935;
wire x_22936;
wire x_22937;
wire x_22938;
wire x_22939;
wire x_22940;
wire x_22941;
wire x_22942;
wire x_22943;
wire x_22944;
wire x_22945;
wire x_22946;
wire x_22947;
wire x_22948;
wire x_22949;
wire x_22950;
wire x_22951;
wire x_22952;
wire x_22953;
wire x_22954;
wire x_22955;
wire x_22956;
wire x_22957;
wire x_22958;
wire x_22959;
wire x_22960;
wire x_22961;
wire x_22962;
wire x_22963;
wire x_22964;
wire x_22965;
wire x_22966;
wire x_22967;
wire x_22968;
wire x_22969;
wire x_22970;
wire x_22971;
wire x_22972;
wire x_22973;
wire x_22974;
wire x_22975;
wire x_22976;
wire x_22977;
wire x_22978;
wire x_22979;
wire x_22980;
wire x_22981;
wire x_22982;
wire x_22983;
wire x_22984;
wire x_22985;
wire x_22986;
wire x_22987;
wire x_22988;
wire x_22989;
wire x_22990;
wire x_22991;
wire x_22992;
wire x_22993;
wire x_22994;
wire x_22995;
wire x_22996;
wire x_22997;
wire x_22998;
wire x_22999;
wire x_23000;
wire x_23001;
wire x_23002;
wire x_23003;
wire x_23004;
wire x_23005;
wire x_23006;
wire x_23007;
wire x_23008;
wire x_23009;
wire x_23010;
wire x_23011;
wire x_23012;
wire x_23013;
wire x_23014;
wire x_23015;
wire x_23016;
wire x_23017;
wire x_23018;
wire x_23019;
wire x_23020;
wire x_23021;
wire x_23022;
wire x_23023;
wire x_23024;
wire x_23025;
wire x_23026;
wire x_23027;
wire x_23028;
wire x_23029;
wire x_23030;
wire x_23031;
wire x_23032;
wire x_23033;
wire x_23034;
wire x_23035;
wire x_23036;
wire x_23037;
wire x_23038;
wire x_23039;
wire x_23040;
wire x_23041;
wire x_23042;
wire x_23043;
wire x_23044;
wire x_23045;
wire x_23046;
wire x_23047;
wire x_23048;
wire x_23049;
wire x_23050;
wire x_23051;
wire x_23052;
wire x_23053;
wire x_23054;
wire x_23055;
wire x_23056;
wire x_23057;
wire x_23058;
wire x_23059;
wire x_23060;
wire x_23061;
wire x_23062;
wire x_23063;
wire x_23064;
wire x_23065;
wire x_23066;
wire x_23067;
wire x_23068;
wire x_23069;
wire x_23070;
wire x_23071;
wire x_23072;
wire x_23073;
wire x_23074;
wire x_23075;
wire x_23076;
wire x_23077;
wire x_23078;
wire x_23079;
wire x_23080;
wire x_23081;
wire x_23082;
wire x_23083;
wire x_23084;
wire x_23085;
wire x_23086;
wire x_23087;
wire x_23088;
wire x_23089;
wire x_23090;
wire x_23091;
wire x_23092;
wire x_23093;
wire x_23094;
wire x_23095;
wire x_23096;
wire x_23097;
wire x_23098;
wire x_23099;
wire x_23100;
wire x_23101;
wire x_23102;
wire x_23103;
wire x_23104;
wire x_23105;
wire x_23106;
wire x_23107;
wire x_23108;
wire x_23109;
wire x_23110;
wire x_23111;
wire x_23112;
wire x_23113;
wire x_23114;
wire x_23115;
wire x_23116;
wire x_23117;
wire x_23118;
wire x_23119;
wire x_23120;
wire x_23121;
wire x_23122;
wire x_23123;
wire x_23124;
wire x_23125;
wire x_23126;
wire x_23127;
wire x_23128;
wire x_23129;
wire x_23130;
wire x_23131;
wire x_23132;
wire x_23133;
wire x_23134;
wire x_23135;
wire x_23136;
wire x_23137;
wire x_23138;
wire x_23139;
wire x_23140;
wire x_23141;
wire x_23142;
wire x_23143;
wire x_23144;
wire x_23145;
wire x_23146;
wire x_23147;
wire x_23148;
wire x_23149;
wire x_23150;
wire x_23151;
wire x_23152;
wire x_23153;
wire x_23154;
wire x_23155;
wire x_23156;
wire x_23157;
wire x_23158;
wire x_23159;
wire x_23160;
wire x_23161;
wire x_23162;
wire x_23163;
wire x_23164;
wire x_23165;
wire x_23166;
wire x_23167;
wire x_23168;
wire x_23169;
wire x_23170;
wire x_23171;
wire x_23172;
wire x_23173;
wire x_23174;
wire x_23175;
wire x_23176;
wire x_23177;
wire x_23178;
wire x_23179;
wire x_23180;
wire x_23181;
wire x_23182;
wire x_23183;
wire x_23184;
wire x_23185;
wire x_23186;
wire x_23187;
wire x_23188;
wire x_23189;
wire x_23190;
wire x_23191;
wire x_23192;
wire x_23193;
wire x_23194;
wire x_23195;
wire x_23196;
wire x_23197;
wire x_23198;
wire x_23199;
wire x_23200;
wire x_23201;
wire x_23202;
wire x_23203;
wire x_23204;
wire x_23205;
wire x_23206;
wire x_23207;
wire x_23208;
wire x_23209;
wire x_23210;
wire x_23211;
wire x_23212;
wire x_23213;
wire x_23214;
wire x_23215;
wire x_23216;
wire x_23217;
wire x_23218;
wire x_23219;
wire x_23220;
wire x_23221;
wire x_23222;
wire x_23223;
wire x_23224;
wire x_23225;
wire x_23226;
wire x_23227;
wire x_23228;
wire x_23229;
wire x_23230;
wire x_23231;
wire x_23232;
wire x_23233;
wire x_23234;
wire x_23235;
wire x_23236;
wire x_23237;
wire x_23238;
wire x_23239;
wire x_23240;
wire x_23241;
wire x_23242;
wire x_23243;
wire x_23244;
wire x_23245;
wire x_23246;
wire x_23247;
wire x_23248;
wire x_23249;
wire x_23250;
wire x_23251;
wire x_23252;
wire x_23253;
wire x_23254;
wire x_23255;
wire x_23256;
wire x_23257;
wire x_23258;
wire x_23259;
wire x_23260;
wire x_23261;
wire x_23262;
wire x_23263;
wire x_23264;
wire x_23265;
wire x_23266;
wire x_23267;
wire x_23268;
wire x_23269;
wire x_23270;
wire x_23271;
wire x_23272;
wire x_23273;
wire x_23274;
wire x_23275;
wire x_23276;
wire x_23277;
wire x_23278;
wire x_23279;
wire x_23280;
wire x_23281;
wire x_23282;
wire x_23283;
wire x_23284;
wire x_23285;
wire x_23286;
wire x_23287;
wire x_23288;
wire x_23289;
wire x_23290;
wire x_23291;
wire x_23292;
wire x_23293;
wire x_23294;
wire x_23295;
wire x_23296;
wire x_23297;
wire x_23298;
wire x_23299;
wire x_23300;
wire x_23301;
wire x_23302;
wire x_23303;
wire x_23304;
wire x_23305;
wire x_23306;
wire x_23307;
wire x_23308;
wire x_23309;
wire x_23310;
wire x_23311;
wire x_23312;
wire x_23313;
wire x_23314;
wire x_23315;
wire x_23316;
wire x_23317;
wire x_23318;
wire x_23319;
wire x_23320;
wire x_23321;
wire x_23322;
wire x_23323;
wire x_23324;
wire x_23325;
wire x_23326;
wire x_23327;
wire x_23328;
wire x_23329;
wire x_23330;
wire x_23331;
wire x_23332;
wire x_23333;
wire x_23334;
wire x_23335;
wire x_23336;
wire x_23337;
wire x_23338;
wire x_23339;
wire x_23340;
wire x_23341;
wire x_23342;
wire x_23343;
wire x_23344;
wire x_23345;
wire x_23346;
wire x_23347;
wire x_23348;
wire x_23349;
wire x_23350;
wire x_23351;
wire x_23352;
wire x_23353;
wire x_23354;
wire x_23355;
wire x_23356;
wire x_23357;
wire x_23358;
wire x_23359;
wire x_23360;
wire x_23361;
wire x_23362;
wire x_23363;
wire x_23364;
wire x_23365;
wire x_23366;
wire x_23367;
wire x_23368;
wire x_23369;
wire x_23370;
wire x_23371;
wire x_23372;
wire x_23373;
wire x_23374;
wire x_23375;
wire x_23376;
wire x_23377;
wire x_23378;
wire x_23379;
wire x_23380;
wire x_23381;
wire x_23382;
wire x_23383;
wire x_23384;
wire x_23385;
wire x_23386;
wire x_23387;
wire x_23388;
wire x_23389;
wire x_23390;
wire x_23391;
wire x_23392;
wire x_23393;
wire x_23394;
wire x_23395;
wire x_23396;
wire x_23397;
wire x_23398;
wire x_23399;
wire x_23400;
wire x_23401;
wire x_23402;
wire x_23403;
wire x_23404;
wire x_23405;
wire x_23406;
wire x_23407;
wire x_23408;
wire x_23409;
wire x_23410;
wire x_23411;
wire x_23412;
wire x_23413;
wire x_23414;
wire x_23415;
wire x_23416;
wire x_23417;
wire x_23418;
wire x_23419;
wire x_23420;
wire x_23421;
wire x_23422;
wire x_23423;
wire x_23424;
wire x_23425;
wire x_23426;
wire x_23427;
wire x_23428;
wire x_23429;
wire x_23430;
wire x_23431;
wire x_23432;
wire x_23433;
wire x_23434;
wire x_23435;
wire x_23436;
wire x_23437;
wire x_23438;
wire x_23439;
wire x_23440;
wire x_23441;
wire x_23442;
wire x_23443;
wire x_23444;
wire x_23445;
wire x_23446;
wire x_23447;
wire x_23448;
wire x_23449;
wire x_23450;
wire x_23451;
wire x_23452;
wire x_23453;
wire x_23454;
wire x_23455;
wire x_23456;
wire x_23457;
wire x_23458;
wire x_23459;
wire x_23460;
wire x_23461;
wire x_23462;
wire x_23463;
wire x_23464;
wire x_23465;
wire x_23466;
wire x_23467;
wire x_23468;
wire x_23469;
wire x_23470;
wire x_23471;
wire x_23472;
wire x_23473;
wire x_23474;
wire x_23475;
wire x_23476;
wire x_23477;
wire x_23478;
wire x_23479;
wire x_23480;
wire x_23481;
wire x_23482;
wire x_23483;
wire x_23484;
wire x_23485;
wire x_23486;
wire x_23487;
wire x_23488;
wire x_23489;
wire x_23490;
wire x_23491;
wire x_23492;
wire x_23493;
wire x_23494;
wire x_23495;
wire x_23496;
wire x_23497;
wire x_23498;
wire x_23499;
wire x_23500;
wire x_23501;
wire x_23502;
wire x_23503;
wire x_23504;
wire x_23505;
wire x_23506;
wire x_23507;
wire x_23508;
wire x_23509;
wire x_23510;
wire x_23511;
wire x_23512;
wire x_23513;
wire x_23514;
wire x_23515;
wire x_23516;
wire x_23517;
wire x_23518;
wire x_23519;
wire x_23520;
wire x_23521;
wire x_23522;
wire x_23523;
wire x_23524;
wire x_23525;
wire x_23526;
wire x_23527;
wire x_23528;
wire x_23529;
wire x_23530;
wire x_23531;
wire x_23532;
wire x_23533;
wire x_23534;
wire x_23535;
wire x_23536;
wire x_23537;
wire x_23538;
wire x_23539;
wire x_23540;
wire x_23541;
wire x_23542;
wire x_23543;
wire x_23544;
wire x_23545;
wire x_23546;
wire x_23547;
wire x_23548;
wire x_23549;
wire x_23550;
wire x_23551;
wire x_23552;
wire x_23553;
wire x_23554;
wire x_23555;
wire x_23556;
wire x_23557;
wire x_23558;
wire x_23559;
wire x_23560;
wire x_23561;
wire x_23562;
wire x_23563;
wire x_23564;
wire x_23565;
wire x_23566;
wire x_23567;
wire x_23568;
wire x_23569;
wire x_23570;
wire x_23571;
wire x_23572;
wire x_23573;
wire x_23574;
wire x_23575;
wire x_23576;
wire x_23577;
wire x_23578;
wire x_23579;
wire x_23580;
wire x_23581;
wire x_23582;
wire x_23583;
wire x_23584;
wire x_23585;
wire x_23586;
wire x_23587;
wire x_23588;
wire x_23589;
wire x_23590;
wire x_23591;
wire x_23592;
wire x_23593;
wire x_23594;
wire x_23595;
wire x_23596;
wire x_23597;
wire x_23598;
wire x_23599;
wire x_23600;
wire x_23601;
wire x_23602;
wire x_23603;
wire x_23604;
wire x_23605;
wire x_23606;
wire x_23607;
wire x_23608;
wire x_23609;
wire x_23610;
wire x_23611;
wire x_23612;
wire x_23613;
wire x_23614;
wire x_23615;
wire x_23616;
wire x_23617;
wire x_23618;
wire x_23619;
wire x_23620;
wire x_23621;
wire x_23622;
wire x_23623;
wire x_23624;
wire x_23625;
wire x_23626;
wire x_23627;
wire x_23628;
wire x_23629;
wire x_23630;
wire x_23631;
wire x_23632;
wire x_23633;
wire x_23634;
wire x_23635;
wire x_23636;
wire x_23637;
wire x_23638;
wire x_23639;
wire x_23640;
wire x_23641;
wire x_23642;
wire x_23643;
wire x_23644;
wire x_23645;
wire x_23646;
wire x_23647;
wire x_23648;
wire x_23649;
wire x_23650;
wire x_23651;
wire x_23652;
wire x_23653;
wire x_23654;
wire x_23655;
wire x_23656;
wire x_23657;
wire x_23658;
wire x_23659;
wire x_23660;
wire x_23661;
wire x_23662;
wire x_23663;
wire x_23664;
wire x_23665;
wire x_23666;
wire x_23667;
wire x_23668;
wire x_23669;
wire x_23670;
wire x_23671;
wire x_23672;
wire x_23673;
wire x_23674;
wire x_23675;
wire x_23676;
wire x_23677;
wire x_23678;
wire x_23679;
wire x_23680;
wire x_23681;
wire x_23682;
wire x_23683;
wire x_23684;
wire x_23685;
wire x_23686;
wire x_23687;
wire x_23688;
wire x_23689;
wire x_23690;
wire x_23691;
wire x_23692;
wire x_23693;
wire x_23694;
wire x_23695;
wire x_23696;
wire x_23697;
wire x_23698;
wire x_23699;
wire x_23700;
wire x_23701;
wire x_23702;
wire x_23703;
wire x_23704;
wire x_23705;
wire x_23706;
wire x_23707;
wire x_23708;
wire x_23709;
wire x_23710;
wire x_23711;
wire x_23712;
wire x_23713;
wire x_23714;
wire x_23715;
wire x_23716;
wire x_23717;
wire x_23718;
wire x_23719;
wire x_23720;
wire x_23721;
wire x_23722;
wire x_23723;
wire x_23724;
wire x_23725;
wire x_23726;
wire x_23727;
wire x_23728;
wire x_23729;
wire x_23730;
wire x_23731;
wire x_23732;
wire x_23733;
wire x_23734;
wire x_23735;
wire x_23736;
wire x_23737;
wire x_23738;
wire x_23739;
wire x_23740;
wire x_23741;
wire x_23742;
wire x_23743;
wire x_23744;
wire x_23745;
wire x_23746;
wire x_23747;
wire x_23748;
wire x_23749;
wire x_23750;
wire x_23751;
wire x_23752;
wire x_23753;
wire x_23754;
wire x_23755;
wire x_23756;
wire x_23757;
wire x_23758;
wire x_23759;
wire x_23760;
wire x_23761;
wire x_23762;
wire x_23763;
wire x_23764;
wire x_23765;
wire x_23766;
wire x_23767;
wire x_23768;
wire x_23769;
wire x_23770;
wire x_23771;
wire x_23772;
wire x_23773;
wire x_23774;
wire x_23775;
wire x_23776;
wire x_23777;
wire x_23778;
wire x_23779;
wire x_23780;
wire x_23781;
wire x_23782;
wire x_23783;
wire x_23784;
wire x_23785;
wire x_23786;
wire x_23787;
wire x_23788;
wire x_23789;
wire x_23790;
wire x_23791;
wire x_23792;
wire x_23793;
wire x_23794;
wire x_23795;
wire x_23796;
wire x_23797;
wire x_23798;
wire x_23799;
wire x_23800;
wire x_23801;
wire x_23802;
wire x_23803;
wire x_23804;
wire x_23805;
wire x_23806;
wire x_23807;
wire x_23808;
wire x_23809;
wire x_23810;
wire x_23811;
wire x_23812;
wire x_23813;
wire x_23814;
wire x_23815;
wire x_23816;
wire x_23817;
wire x_23818;
wire x_23819;
wire x_23820;
wire x_23821;
wire x_23822;
wire x_23823;
wire x_23824;
wire x_23825;
wire x_23826;
wire x_23827;
wire x_23828;
wire x_23829;
wire x_23830;
wire x_23831;
wire x_23832;
wire x_23833;
wire x_23834;
wire x_23835;
wire x_23836;
wire x_23837;
wire x_23838;
wire x_23839;
wire x_23840;
wire x_23841;
wire x_23842;
wire x_23843;
wire x_23844;
wire x_23845;
wire x_23846;
wire x_23847;
wire x_23848;
wire x_23849;
wire x_23850;
wire x_23851;
wire x_23852;
wire x_23853;
wire x_23854;
wire x_23855;
wire x_23856;
wire x_23857;
wire x_23858;
wire x_23859;
wire x_23860;
wire x_23861;
wire x_23862;
wire x_23863;
wire x_23864;
wire x_23865;
wire x_23866;
wire x_23867;
wire x_23868;
wire x_23869;
wire x_23870;
wire x_23871;
wire x_23872;
wire x_23873;
wire x_23874;
wire x_23875;
wire x_23876;
wire x_23877;
wire x_23878;
wire x_23879;
wire x_23880;
wire x_23881;
wire x_23882;
wire x_23883;
wire x_23884;
wire x_23885;
wire x_23886;
wire x_23887;
wire x_23888;
wire x_23889;
wire x_23890;
wire x_23891;
wire x_23892;
wire x_23893;
wire x_23894;
wire x_23895;
wire x_23896;
wire x_23897;
wire x_23898;
wire x_23899;
wire x_23900;
wire x_23901;
wire x_23902;
wire x_23903;
wire x_23904;
wire x_23905;
wire x_23906;
wire x_23907;
wire x_23908;
wire x_23909;
wire x_23910;
wire x_23911;
wire x_23912;
wire x_23913;
wire x_23914;
wire x_23915;
wire x_23916;
wire x_23917;
wire x_23918;
wire x_23919;
wire x_23920;
wire x_23921;
wire x_23922;
wire x_23923;
wire x_23924;
wire x_23925;
wire x_23926;
wire x_23927;
wire x_23928;
wire x_23929;
wire x_23930;
wire x_23931;
wire x_23932;
wire x_23933;
wire x_23934;
wire x_23935;
wire x_23936;
wire x_23937;
wire x_23938;
wire x_23939;
wire x_23940;
wire x_23941;
wire x_23942;
wire x_23943;
wire x_23944;
wire x_23945;
wire x_23946;
wire x_23947;
wire x_23948;
wire x_23949;
wire x_23950;
wire x_23951;
wire x_23952;
wire x_23953;
wire x_23954;
wire x_23955;
wire x_23956;
wire x_23957;
wire x_23958;
wire x_23959;
wire x_23960;
wire x_23961;
wire x_23962;
wire x_23963;
wire x_23964;
wire x_23965;
wire x_23966;
wire x_23967;
wire x_23968;
wire x_23969;
wire x_23970;
wire x_23971;
wire x_23972;
wire x_23973;
wire x_23974;
wire x_23975;
wire x_23976;
wire x_23977;
wire x_23978;
wire x_23979;
wire x_23980;
wire x_23981;
wire x_23982;
wire x_23983;
wire x_23984;
wire x_23985;
wire x_23986;
wire x_23987;
wire x_23988;
wire x_23989;
wire x_23990;
wire x_23991;
wire x_23992;
wire x_23993;
wire x_23994;
wire x_23995;
wire x_23996;
wire x_23997;
wire x_23998;
wire x_23999;
wire x_24000;
wire x_24001;
wire x_24002;
wire x_24003;
wire x_24004;
wire x_24005;
wire x_24006;
wire x_24007;
wire x_24008;
wire x_24009;
wire x_24010;
wire x_24011;
wire x_24012;
wire x_24013;
wire x_24014;
wire x_24015;
wire x_24016;
wire x_24017;
wire x_24018;
wire x_24019;
wire x_24020;
wire x_24021;
wire x_24022;
wire x_24023;
wire x_24024;
wire x_24025;
wire x_24026;
wire x_24027;
wire x_24028;
wire x_24029;
wire x_24030;
wire x_24031;
wire x_24032;
wire x_24033;
wire x_24034;
wire x_24035;
wire x_24036;
wire x_24037;
wire x_24038;
wire x_24039;
wire x_24040;
wire x_24041;
wire x_24042;
wire x_24043;
wire x_24044;
wire x_24045;
wire x_24046;
wire x_24047;
wire x_24048;
wire x_24049;
wire x_24050;
wire x_24051;
wire x_24052;
wire x_24053;
wire x_24054;
wire x_24055;
wire x_24056;
wire x_24057;
wire x_24058;
wire x_24059;
wire x_24060;
wire x_24061;
wire x_24062;
wire x_24063;
wire x_24064;
wire x_24065;
wire x_24066;
wire x_24067;
wire x_24068;
wire x_24069;
wire x_24070;
wire x_24071;
wire x_24072;
wire x_24073;
wire x_24074;
wire x_24075;
wire x_24076;
wire x_24077;
wire x_24078;
wire x_24079;
wire x_24080;
wire x_24081;
wire x_24082;
wire x_24083;
wire x_24084;
wire x_24085;
wire x_24086;
wire x_24087;
wire x_24088;
wire x_24089;
wire x_24090;
wire x_24091;
wire x_24092;
wire x_24093;
wire x_24094;
wire x_24095;
wire x_24096;
wire x_24097;
wire x_24098;
wire x_24099;
wire x_24100;
wire x_24101;
wire x_24102;
wire x_24103;
wire x_24104;
wire x_24105;
wire x_24106;
wire x_24107;
wire x_24108;
wire x_24109;
wire x_24110;
wire x_24111;
wire x_24112;
wire x_24113;
wire x_24114;
wire x_24115;
wire x_24116;
wire x_24117;
wire x_24118;
wire x_24119;
wire x_24120;
wire x_24121;
wire x_24122;
wire x_24123;
wire x_24124;
wire x_24125;
wire x_24126;
wire x_24127;
wire x_24128;
wire x_24129;
wire x_24130;
wire x_24131;
wire x_24132;
wire x_24133;
wire x_24134;
wire x_24135;
wire x_24136;
wire x_24137;
wire x_24138;
wire x_24139;
wire x_24140;
wire x_24141;
wire x_24142;
wire x_24143;
wire x_24144;
wire x_24145;
wire x_24146;
wire x_24147;
wire x_24148;
wire x_24149;
wire x_24150;
wire x_24151;
wire x_24152;
wire x_24153;
wire x_24154;
wire x_24155;
wire x_24156;
wire x_24157;
wire x_24158;
wire x_24159;
wire x_24160;
wire x_24161;
wire x_24162;
wire x_24163;
wire x_24164;
wire x_24165;
wire x_24166;
wire x_24167;
wire x_24168;
wire x_24169;
wire x_24170;
wire x_24171;
wire x_24172;
wire x_24173;
wire x_24174;
wire x_24175;
wire x_24176;
wire x_24177;
wire x_24178;
wire x_24179;
wire x_24180;
wire x_24181;
wire x_24182;
wire x_24183;
wire x_24184;
wire x_24185;
wire x_24186;
wire x_24187;
wire x_24188;
wire x_24189;
wire x_24190;
wire x_24191;
wire x_24192;
wire x_24193;
wire x_24194;
wire x_24195;
wire x_24196;
wire x_24197;
wire x_24198;
wire x_24199;
wire x_24200;
wire x_24201;
wire x_24202;
wire x_24203;
wire x_24204;
wire x_24205;
wire x_24206;
wire x_24207;
wire x_24208;
wire x_24209;
wire x_24210;
wire x_24211;
wire x_24212;
wire x_24213;
wire x_24214;
wire x_24215;
wire x_24216;
wire x_24217;
wire x_24218;
wire x_24219;
wire x_24220;
wire x_24221;
wire x_24222;
wire x_24223;
wire x_24224;
wire x_24225;
wire x_24226;
wire x_24227;
wire x_24228;
wire x_24229;
wire x_24230;
wire x_24231;
wire x_24232;
wire x_24233;
wire x_24234;
wire x_24235;
wire x_24236;
wire x_24237;
wire x_24238;
wire x_24239;
wire x_24240;
wire x_24241;
wire x_24242;
wire x_24243;
wire x_24244;
wire x_24245;
wire x_24246;
wire x_24247;
wire x_24248;
wire x_24249;
wire x_24250;
wire x_24251;
wire x_24252;
wire x_24253;
wire x_24254;
wire x_24255;
wire x_24256;
wire x_24257;
wire x_24258;
wire x_24259;
wire x_24260;
wire x_24261;
wire x_24262;
wire x_24263;
wire x_24264;
wire x_24265;
wire x_24266;
wire x_24267;
wire x_24268;
wire x_24269;
wire x_24270;
wire x_24271;
wire x_24272;
wire x_24273;
wire x_24274;
wire x_24275;
wire x_24276;
wire x_24277;
wire x_24278;
wire x_24279;
wire x_24280;
wire x_24281;
wire x_24282;
wire x_24283;
wire x_24284;
wire x_24285;
wire x_24286;
wire x_24287;
wire x_24288;
wire x_24289;
wire x_24290;
wire x_24291;
wire x_24292;
wire x_24293;
wire x_24294;
wire x_24295;
wire x_24296;
wire x_24297;
wire x_24298;
wire x_24299;
wire x_24300;
wire x_24301;
wire x_24302;
wire x_24303;
wire x_24304;
wire x_24305;
wire x_24306;
wire x_24307;
wire x_24308;
wire x_24309;
wire x_24310;
wire x_24311;
wire x_24312;
wire x_24313;
wire x_24314;
wire x_24315;
wire x_24316;
wire x_24317;
wire x_24318;
wire x_24319;
wire x_24320;
wire x_24321;
wire x_24322;
wire x_24323;
wire x_24324;
wire x_24325;
wire x_24326;
wire x_24327;
wire x_24328;
wire x_24329;
wire x_24330;
wire x_24331;
wire x_24332;
wire x_24333;
wire x_24334;
wire x_24335;
wire x_24336;
wire x_24337;
wire x_24338;
wire x_24339;
wire x_24340;
wire x_24341;
wire x_24342;
wire x_24343;
wire x_24344;
wire x_24345;
wire x_24346;
wire x_24347;
wire x_24348;
wire x_24349;
wire x_24350;
wire x_24351;
wire x_24352;
wire x_24353;
wire x_24354;
wire x_24355;
wire x_24356;
wire x_24357;
wire x_24358;
wire x_24359;
wire x_24360;
wire x_24361;
wire x_24362;
wire x_24363;
wire x_24364;
wire x_24365;
wire x_24366;
wire x_24367;
wire x_24368;
wire x_24369;
wire x_24370;
wire x_24371;
wire x_24372;
wire x_24373;
wire x_24374;
wire x_24375;
wire x_24376;
wire x_24377;
wire x_24378;
wire x_24379;
wire x_24380;
wire x_24381;
wire x_24382;
wire x_24383;
wire x_24384;
wire x_24385;
wire x_24386;
wire x_24387;
wire x_24388;
wire x_24389;
wire x_24390;
wire x_24391;
wire x_24392;
wire x_24393;
wire x_24394;
wire x_24395;
wire x_24396;
wire x_24397;
wire x_24398;
wire x_24399;
wire x_24400;
wire x_24401;
wire x_24402;
wire x_24403;
wire x_24404;
wire x_24405;
wire x_24406;
wire x_24407;
wire x_24408;
wire x_24409;
wire x_24410;
wire x_24411;
wire x_24412;
wire x_24413;
wire x_24414;
wire x_24415;
wire x_24416;
wire x_24417;
wire x_24418;
wire x_24419;
wire x_24420;
wire x_24421;
wire x_24422;
wire x_24423;
wire x_24424;
wire x_24425;
wire x_24426;
wire x_24427;
wire x_24428;
wire x_24429;
wire x_24430;
wire x_24431;
wire x_24432;
wire x_24433;
wire x_24434;
wire x_24435;
wire x_24436;
wire x_24437;
wire x_24438;
wire x_24439;
wire x_24440;
wire x_24441;
wire x_24442;
wire x_24443;
wire x_24444;
wire x_24445;
wire x_24446;
wire x_24447;
wire x_24448;
wire x_24449;
wire x_24450;
wire x_24451;
wire x_24452;
wire x_24453;
wire x_24454;
wire x_24455;
wire x_24456;
wire x_24457;
wire x_24458;
wire x_24459;
wire x_24460;
wire x_24461;
wire x_24462;
wire x_24463;
wire x_24464;
wire x_24465;
wire x_24466;
wire x_24467;
wire x_24468;
wire x_24469;
wire x_24470;
wire x_24471;
wire x_24472;
wire x_24473;
wire x_24474;
wire x_24475;
wire x_24476;
wire x_24477;
wire x_24478;
wire x_24479;
wire x_24480;
wire x_24481;
wire x_24482;
wire x_24483;
wire x_24484;
wire x_24485;
wire x_24486;
wire x_24487;
wire x_24488;
wire x_24489;
wire x_24490;
wire x_24491;
wire x_24492;
wire x_24493;
wire x_24494;
wire x_24495;
wire x_24496;
wire x_24497;
wire x_24498;
wire x_24499;
wire x_24500;
wire x_24501;
wire x_24502;
wire x_24503;
wire x_24504;
wire x_24505;
wire x_24506;
wire x_24507;
wire x_24508;
wire x_24509;
wire x_24510;
wire x_24511;
wire x_24512;
wire x_24513;
wire x_24514;
wire x_24515;
wire x_24516;
wire x_24517;
wire x_24518;
wire x_24519;
wire x_24520;
wire x_24521;
wire x_24522;
wire x_24523;
wire x_24524;
wire x_24525;
wire x_24526;
wire x_24527;
wire x_24528;
wire x_24529;
wire x_24530;
wire x_24531;
wire x_24532;
wire x_24533;
wire x_24534;
wire x_24535;
wire x_24536;
wire x_24537;
wire x_24538;
wire x_24539;
wire x_24540;
wire x_24541;
wire x_24542;
wire x_24543;
wire x_24544;
wire x_24545;
wire x_24546;
wire x_24547;
wire x_24548;
wire x_24549;
wire x_24550;
wire x_24551;
wire x_24552;
wire x_24553;
wire x_24554;
wire x_24555;
wire x_24556;
wire x_24557;
wire x_24558;
wire x_24559;
wire x_24560;
wire x_24561;
wire x_24562;
wire x_24563;
wire x_24564;
wire x_24565;
wire x_24566;
wire x_24567;
wire x_24568;
wire x_24569;
wire x_24570;
wire x_24571;
wire x_24572;
wire x_24573;
wire x_24574;
wire x_24575;
wire x_24576;
wire x_24577;
wire x_24578;
wire x_24579;
wire x_24580;
wire x_24581;
wire x_24582;
wire x_24583;
wire x_24584;
wire x_24585;
wire x_24586;
wire x_24587;
wire x_24588;
wire x_24589;
wire x_24590;
wire x_24591;
wire x_24592;
wire x_24593;
wire x_24594;
wire x_24595;
wire x_24596;
wire x_24597;
wire x_24598;
wire x_24599;
wire x_24600;
wire x_24601;
wire x_24602;
wire x_24603;
wire x_24604;
wire x_24605;
wire x_24606;
wire x_24607;
wire x_24608;
wire x_24609;
wire x_24610;
wire x_24611;
wire x_24612;
wire x_24613;
wire x_24614;
wire x_24615;
wire x_24616;
wire x_24617;
wire x_24618;
wire x_24619;
wire x_24620;
wire x_24621;
wire x_24622;
wire x_24623;
wire x_24624;
wire x_24625;
wire x_24626;
wire x_24627;
wire x_24628;
wire x_24629;
wire x_24630;
wire x_24631;
wire x_24632;
wire x_24633;
wire x_24634;
wire x_24635;
wire x_24636;
wire x_24637;
wire x_24638;
wire x_24639;
wire x_24640;
wire x_24641;
wire x_24642;
wire x_24643;
wire x_24644;
wire x_24645;
wire x_24646;
wire x_24647;
wire x_24648;
wire x_24649;
wire x_24650;
wire x_24651;
wire x_24652;
wire x_24653;
wire x_24654;
wire x_24655;
wire x_24656;
wire x_24657;
wire x_24658;
wire x_24659;
wire x_24660;
wire x_24661;
wire x_24662;
wire x_24663;
wire x_24664;
wire x_24665;
wire x_24666;
wire x_24667;
wire x_24668;
wire x_24669;
wire x_24670;
wire x_24671;
wire x_24672;
wire x_24673;
wire x_24674;
wire x_24675;
wire x_24676;
wire x_24677;
wire x_24678;
wire x_24679;
wire x_24680;
wire x_24681;
wire x_24682;
wire x_24683;
wire x_24684;
wire x_24685;
wire x_24686;
wire x_24687;
wire x_24688;
wire x_24689;
wire x_24690;
wire x_24691;
wire x_24692;
wire x_24693;
wire x_24694;
wire x_24695;
wire x_24696;
wire x_24697;
wire x_24698;
wire x_24699;
wire x_24700;
wire x_24701;
wire x_24702;
wire x_24703;
wire x_24704;
wire x_24705;
wire x_24706;
wire x_24707;
wire x_24708;
wire x_24709;
wire x_24710;
wire x_24711;
wire x_24712;
wire x_24713;
wire x_24714;
wire x_24715;
wire x_24716;
wire x_24717;
wire x_24718;
wire x_24719;
wire x_24720;
wire x_24721;
wire x_24722;
wire x_24723;
wire x_24724;
wire x_24725;
wire x_24726;
wire x_24727;
wire x_24728;
wire x_24729;
wire x_24730;
wire x_24731;
wire x_24732;
wire x_24733;
wire x_24734;
wire x_24735;
wire x_24736;
wire x_24737;
wire x_24738;
wire x_24739;
wire x_24740;
wire x_24741;
wire x_24742;
wire x_24743;
wire x_24744;
wire x_24745;
wire x_24746;
wire x_24747;
wire x_24748;
wire x_24749;
wire x_24750;
wire x_24751;
wire x_24752;
wire x_24753;
wire x_24754;
wire x_24755;
wire x_24756;
wire x_24757;
wire x_24758;
wire x_24759;
wire x_24760;
wire x_24761;
wire x_24762;
wire x_24763;
wire x_24764;
wire x_24765;
wire x_24766;
wire x_24767;
wire x_24768;
wire x_24769;
wire x_24770;
wire x_24771;
wire x_24772;
wire x_24773;
wire x_24774;
wire x_24775;
wire x_24776;
wire x_24777;
wire x_24778;
wire x_24779;
wire x_24780;
wire x_24781;
wire x_24782;
wire x_24783;
wire x_24784;
wire x_24785;
wire x_24786;
wire x_24787;
wire x_24788;
wire x_24789;
wire x_24790;
wire x_24791;
wire x_24792;
wire x_24793;
wire x_24794;
wire x_24795;
wire x_24796;
wire x_24797;
wire x_24798;
wire x_24799;
wire x_24800;
wire x_24801;
wire x_24802;
wire x_24803;
wire x_24804;
wire x_24805;
wire x_24806;
wire x_24807;
wire x_24808;
wire x_24809;
wire x_24810;
wire x_24811;
wire x_24812;
wire x_24813;
wire x_24814;
wire x_24815;
wire x_24816;
wire x_24817;
wire x_24818;
wire x_24819;
wire x_24820;
wire x_24821;
wire x_24822;
wire x_24823;
wire x_24824;
wire x_24825;
wire x_24826;
wire x_24827;
wire x_24828;
wire x_24829;
wire x_24830;
wire x_24831;
wire x_24832;
wire x_24833;
wire x_24834;
wire x_24835;
wire x_24836;
wire x_24837;
wire x_24838;
wire x_24839;
wire x_24840;
wire x_24841;
wire x_24842;
wire x_24843;
wire x_24844;
wire x_24845;
wire x_24846;
wire x_24847;
wire x_24848;
wire x_24849;
wire x_24850;
wire x_24851;
wire x_24852;
wire x_24853;
wire x_24854;
wire x_24855;
wire x_24856;
wire x_24857;
wire x_24858;
wire x_24859;
wire x_24860;
wire x_24861;
wire x_24862;
wire x_24863;
wire x_24864;
wire x_24865;
wire x_24866;
wire x_24867;
wire x_24868;
wire x_24869;
wire x_24870;
wire x_24871;
wire x_24872;
wire x_24873;
wire x_24874;
wire x_24875;
wire x_24876;
wire x_24877;
wire x_24878;
wire x_24879;
wire x_24880;
wire x_24881;
wire x_24882;
wire x_24883;
wire x_24884;
wire x_24885;
wire x_24886;
wire x_24887;
wire x_24888;
wire x_24889;
wire x_24890;
wire x_24891;
wire x_24892;
wire x_24893;
wire x_24894;
wire x_24895;
wire x_24896;
wire x_24897;
wire x_24898;
wire x_24899;
wire x_24900;
wire x_24901;
wire x_24902;
wire x_24903;
wire x_24904;
wire x_24905;
wire x_24906;
wire x_24907;
wire x_24908;
wire x_24909;
wire x_24910;
wire x_24911;
wire x_24912;
wire x_24913;
wire x_24914;
wire x_24915;
wire x_24916;
wire x_24917;
wire x_24918;
wire x_24919;
wire x_24920;
wire x_24921;
wire x_24922;
wire x_24923;
wire x_24924;
wire x_24925;
wire x_24926;
wire x_24927;
wire x_24928;
wire x_24929;
wire x_24930;
wire x_24931;
wire x_24932;
wire x_24933;
wire x_24934;
wire x_24935;
wire x_24936;
wire x_24937;
wire x_24938;
wire x_24939;
wire x_24940;
wire x_24941;
wire x_24942;
wire x_24943;
wire x_24944;
wire x_24945;
wire x_24946;
wire x_24947;
wire x_24948;
wire x_24949;
wire x_24950;
wire x_24951;
wire x_24952;
wire x_24953;
wire x_24954;
wire x_24955;
wire x_24956;
wire x_24957;
wire x_24958;
wire x_24959;
wire x_24960;
wire x_24961;
wire x_24962;
wire x_24963;
wire x_24964;
wire x_24965;
wire x_24966;
wire x_24967;
wire x_24968;
wire x_24969;
wire x_24970;
wire x_24971;
wire x_24972;
wire x_24973;
wire x_24974;
wire x_24975;
wire x_24976;
wire x_24977;
wire x_24978;
wire x_24979;
wire x_24980;
wire x_24981;
wire x_24982;
wire x_24983;
wire x_24984;
wire x_24985;
wire x_24986;
wire x_24987;
wire x_24988;
wire x_24989;
wire x_24990;
wire x_24991;
wire x_24992;
wire x_24993;
wire x_24994;
wire x_24995;
wire x_24996;
wire x_24997;
wire x_24998;
wire x_24999;
wire x_25000;
wire x_25001;
wire x_25002;
wire x_25003;
wire x_25004;
wire x_25005;
wire x_25006;
wire x_25007;
wire x_25008;
wire x_25009;
wire x_25010;
wire x_25011;
wire x_25012;
wire x_25013;
wire x_25014;
wire x_25015;
wire x_25016;
wire x_25017;
wire x_25018;
wire x_25019;
wire x_25020;
wire x_25021;
wire x_25022;
wire x_25023;
wire x_25024;
wire x_25025;
wire x_25026;
wire x_25027;
wire x_25028;
wire x_25029;
wire x_25030;
wire x_25031;
wire x_25032;
wire x_25033;
wire x_25034;
wire x_25035;
wire x_25036;
wire x_25037;
wire x_25038;
wire x_25039;
wire x_25040;
wire x_25041;
wire x_25042;
wire x_25043;
wire x_25044;
wire x_25045;
wire x_25046;
wire x_25047;
wire x_25048;
wire x_25049;
wire x_25050;
wire x_25051;
wire x_25052;
wire x_25053;
wire x_25054;
wire x_25055;
wire x_25056;
wire x_25057;
wire x_25058;
wire x_25059;
wire x_25060;
wire x_25061;
wire x_25062;
wire x_25063;
wire x_25064;
wire x_25065;
wire x_25066;
wire x_25067;
wire x_25068;
wire x_25069;
wire x_25070;
wire x_25071;
wire x_25072;
wire x_25073;
wire x_25074;
wire x_25075;
wire x_25076;
wire x_25077;
wire x_25078;
wire x_25079;
wire x_25080;
wire x_25081;
wire x_25082;
wire x_25083;
wire x_25084;
wire x_25085;
wire x_25086;
wire x_25087;
wire x_25088;
wire x_25089;
wire x_25090;
wire x_25091;
wire x_25092;
wire x_25093;
wire x_25094;
wire x_25095;
wire x_25096;
wire x_25097;
wire x_25098;
wire x_25099;
wire x_25100;
wire x_25101;
wire x_25102;
wire x_25103;
wire x_25104;
wire x_25105;
wire x_25106;
wire x_25107;
wire x_25108;
wire x_25109;
wire x_25110;
wire x_25111;
wire x_25112;
wire x_25113;
wire x_25114;
wire x_25115;
wire x_25116;
wire x_25117;
wire x_25118;
wire x_25119;
wire x_25120;
wire x_25121;
wire x_25122;
wire x_25123;
wire x_25124;
wire x_25125;
wire x_25126;
wire x_25127;
wire x_25128;
wire x_25129;
wire x_25130;
wire x_25131;
wire x_25132;
wire x_25133;
wire x_25134;
wire x_25135;
wire x_25136;
wire x_25137;
wire x_25138;
wire x_25139;
wire x_25140;
wire x_25141;
wire x_25142;
wire x_25143;
wire x_25144;
wire x_25145;
wire x_25146;
wire x_25147;
wire x_25148;
wire x_25149;
wire x_25150;
wire x_25151;
wire x_25152;
wire x_25153;
wire x_25154;
wire x_25155;
wire x_25156;
wire x_25157;
wire x_25158;
wire x_25159;
wire x_25160;
wire x_25161;
wire x_25162;
wire x_25163;
wire x_25164;
wire x_25165;
wire x_25166;
wire x_25167;
wire x_25168;
wire x_25169;
wire x_25170;
wire x_25171;
wire x_25172;
wire x_25173;
wire x_25174;
wire x_25175;
wire x_25176;
wire x_25177;
wire x_25178;
wire x_25179;
wire x_25180;
wire x_25181;
wire x_25182;
wire x_25183;
wire x_25184;
wire x_25185;
wire x_25186;
wire x_25187;
wire x_25188;
wire x_25189;
wire x_25190;
wire x_25191;
wire x_25192;
wire x_25193;
wire x_25194;
wire x_25195;
wire x_25196;
wire x_25197;
wire x_25198;
wire x_25199;
wire x_25200;
wire x_25201;
wire x_25202;
wire x_25203;
wire x_25204;
wire x_25205;
wire x_25206;
wire x_25207;
wire x_25208;
wire x_25209;
wire x_25210;
wire x_25211;
wire x_25212;
wire x_25213;
wire x_25214;
wire x_25215;
wire x_25216;
wire x_25217;
wire x_25218;
wire x_25219;
wire x_25220;
wire x_25221;
wire x_25222;
wire x_25223;
wire x_25224;
wire x_25225;
wire x_25226;
wire x_25227;
wire x_25228;
wire x_25229;
wire x_25230;
wire x_25231;
wire x_25232;
wire x_25233;
wire x_25234;
wire x_25235;
wire x_25236;
wire x_25237;
wire x_25238;
wire x_25239;
wire x_25240;
wire x_25241;
wire x_25242;
wire x_25243;
wire x_25244;
wire x_25245;
wire x_25246;
wire x_25247;
wire x_25248;
wire x_25249;
wire x_25250;
wire x_25251;
wire x_25252;
wire x_25253;
wire x_25254;
wire x_25255;
wire x_25256;
wire x_25257;
wire x_25258;
wire x_25259;
wire x_25260;
wire x_25261;
wire x_25262;
wire x_25263;
wire x_25264;
wire x_25265;
wire x_25266;
wire x_25267;
wire x_25268;
wire x_25269;
wire x_25270;
wire x_25271;
wire x_25272;
wire x_25273;
wire x_25274;
wire x_25275;
wire x_25276;
wire x_25277;
wire x_25278;
wire x_25279;
wire x_25280;
wire x_25281;
wire x_25282;
wire x_25283;
wire x_25284;
wire x_25285;
wire x_25286;
wire x_25287;
wire x_25288;
wire x_25289;
wire x_25290;
wire x_25291;
wire x_25292;
wire x_25293;
wire x_25294;
wire x_25295;
wire x_25296;
wire x_25297;
wire x_25298;
wire x_25299;
wire x_25300;
wire x_25301;
wire x_25302;
wire x_25303;
wire x_25304;
wire x_25305;
wire x_25306;
wire x_25307;
wire x_25308;
wire x_25309;
wire x_25310;
wire x_25311;
wire x_25312;
wire x_25313;
wire x_25314;
wire x_25315;
wire x_25316;
wire x_25317;
wire x_25318;
wire x_25319;
wire x_25320;
wire x_25321;
wire x_25322;
wire x_25323;
wire x_25324;
wire x_25325;
wire x_25326;
wire x_25327;
wire x_25328;
wire x_25329;
wire x_25330;
wire x_25331;
wire x_25332;
wire x_25333;
wire x_25334;
wire x_25335;
wire x_25336;
wire x_25337;
wire x_25338;
wire x_25339;
wire x_25340;
wire x_25341;
wire x_25342;
wire x_25343;
wire x_25344;
wire x_25345;
wire x_25346;
wire x_25347;
wire x_25348;
wire x_25349;
wire x_25350;
wire x_25351;
wire x_25352;
wire x_25353;
wire x_25354;
wire x_25355;
wire x_25356;
wire x_25357;
wire x_25358;
wire x_25359;
wire x_25360;
wire x_25361;
wire x_25362;
wire x_25363;
wire x_25364;
wire x_25365;
wire x_25366;
wire x_25367;
wire x_25368;
wire x_25369;
wire x_25370;
wire x_25371;
wire x_25372;
wire x_25373;
wire x_25374;
wire x_25375;
wire x_25376;
wire x_25377;
wire x_25378;
wire x_25379;
wire x_25380;
wire x_25381;
wire x_25382;
wire x_25383;
wire x_25384;
wire x_25385;
wire x_25386;
wire x_25387;
wire x_25388;
wire x_25389;
wire x_25390;
wire x_25391;
wire x_25392;
wire x_25393;
wire x_25394;
wire x_25395;
wire x_25396;
wire x_25397;
wire x_25398;
wire x_25399;
wire x_25400;
wire x_25401;
wire x_25402;
wire x_25403;
wire x_25404;
wire x_25405;
wire x_25406;
wire x_25407;
wire x_25408;
wire x_25409;
wire x_25410;
wire x_25411;
wire x_25412;
wire x_25413;
wire x_25414;
wire x_25415;
wire x_25416;
wire x_25417;
wire x_25418;
wire x_25419;
wire x_25420;
wire x_25421;
wire x_25422;
wire x_25423;
wire x_25424;
wire x_25425;
wire x_25426;
wire x_25427;
wire x_25428;
wire x_25429;
wire x_25430;
wire x_25431;
wire x_25432;
wire x_25433;
wire x_25434;
wire x_25435;
wire x_25436;
wire x_25437;
wire x_25438;
wire x_25439;
wire x_25440;
wire x_25441;
wire x_25442;
wire x_25443;
wire x_25444;
wire x_25445;
wire x_25446;
wire x_25447;
wire x_25448;
wire x_25449;
wire x_25450;
wire x_25451;
wire x_25452;
wire x_25453;
wire x_25454;
wire x_25455;
wire x_25456;
wire x_25457;
wire x_25458;
wire x_25459;
wire x_25460;
wire x_25461;
wire x_25462;
wire x_25463;
wire x_25464;
wire x_25465;
wire x_25466;
wire x_25467;
wire x_25468;
wire x_25469;
wire x_25470;
wire x_25471;
wire x_25472;
wire x_25473;
wire x_25474;
wire x_25475;
wire x_25476;
wire x_25477;
wire x_25478;
wire x_25479;
wire x_25480;
wire x_25481;
wire x_25482;
wire x_25483;
wire x_25484;
wire x_25485;
wire x_25486;
wire x_25487;
wire x_25488;
wire x_25489;
wire x_25490;
wire x_25491;
wire x_25492;
wire x_25493;
wire x_25494;
wire x_25495;
wire x_25496;
wire x_25497;
wire x_25498;
wire x_25499;
wire x_25500;
wire x_25501;
wire x_25502;
wire x_25503;
wire x_25504;
wire x_25505;
wire x_25506;
wire x_25507;
wire x_25508;
wire x_25509;
wire x_25510;
wire x_25511;
wire x_25512;
wire x_25513;
wire x_25514;
wire x_25515;
wire x_25516;
wire x_25517;
wire x_25518;
wire x_25519;
wire x_25520;
wire x_25521;
wire x_25522;
wire x_25523;
wire x_25524;
wire x_25525;
wire x_25526;
wire x_25527;
wire x_25528;
wire x_25529;
wire x_25530;
wire x_25531;
wire x_25532;
wire x_25533;
wire x_25534;
wire x_25535;
wire x_25536;
wire x_25537;
wire x_25538;
wire x_25539;
wire x_25540;
wire x_25541;
wire x_25542;
wire x_25543;
wire x_25544;
wire x_25545;
wire x_25546;
wire x_25547;
wire x_25548;
wire x_25549;
wire x_25550;
wire x_25551;
wire x_25552;
wire x_25553;
wire x_25554;
wire x_25555;
wire x_25556;
wire x_25557;
wire x_25558;
wire x_25559;
wire x_25560;
wire x_25561;
wire x_25562;
wire x_25563;
wire x_25564;
wire x_25565;
wire x_25566;
wire x_25567;
wire x_25568;
wire x_25569;
wire x_25570;
wire x_25571;
wire x_25572;
wire x_25573;
wire x_25574;
wire x_25575;
wire x_25576;
wire x_25577;
wire x_25578;
wire x_25579;
wire x_25580;
wire x_25581;
wire x_25582;
wire x_25583;
wire x_25584;
wire x_25585;
wire x_25586;
wire x_25587;
wire x_25588;
wire x_25589;
wire x_25590;
wire x_25591;
wire x_25592;
wire x_25593;
wire x_25594;
wire x_25595;
wire x_25596;
wire x_25597;
wire x_25598;
wire x_25599;
wire x_25600;
wire x_25601;
wire x_25602;
wire x_25603;
wire x_25604;
wire x_25605;
wire x_25606;
wire x_25607;
wire x_25608;
wire x_25609;
wire x_25610;
wire x_25611;
wire x_25612;
wire x_25613;
wire x_25614;
wire x_25615;
wire x_25616;
wire x_25617;
wire x_25618;
wire x_25619;
wire x_25620;
wire x_25621;
wire x_25622;
wire x_25623;
wire x_25624;
wire x_25625;
wire x_25626;
wire x_25627;
wire x_25628;
wire x_25629;
wire x_25630;
wire x_25631;
wire x_25632;
wire x_25633;
wire x_25634;
wire x_25635;
wire x_25636;
wire x_25637;
wire x_25638;
wire x_25639;
wire x_25640;
wire x_25641;
wire x_25642;
wire x_25643;
wire x_25644;
wire x_25645;
wire x_25646;
wire x_25647;
wire x_25648;
wire x_25649;
wire x_25650;
wire x_25651;
wire x_25652;
wire x_25653;
wire x_25654;
wire x_25655;
wire x_25656;
wire x_25657;
wire x_25658;
wire x_25659;
wire x_25660;
wire x_25661;
wire x_25662;
wire x_25663;
wire x_25664;
wire x_25665;
wire x_25666;
wire x_25667;
wire x_25668;
wire x_25669;
wire x_25670;
wire x_25671;
wire x_25672;
wire x_25673;
wire x_25674;
wire x_25675;
wire x_25676;
wire x_25677;
wire x_25678;
wire x_25679;
wire x_25680;
wire x_25681;
wire x_25682;
wire x_25683;
wire x_25684;
wire x_25685;
wire x_25686;
wire x_25687;
wire x_25688;
wire x_25689;
wire x_25690;
wire x_25691;
wire x_25692;
wire x_25693;
wire x_25694;
wire x_25695;
wire x_25696;
wire x_25697;
wire x_25698;
wire x_25699;
wire x_25700;
wire x_25701;
wire x_25702;
wire x_25703;
wire x_25704;
wire x_25705;
wire x_25706;
wire x_25707;
wire x_25708;
wire x_25709;
wire x_25710;
wire x_25711;
wire x_25712;
wire x_25713;
wire x_25714;
wire x_25715;
wire x_25716;
wire x_25717;
wire x_25718;
wire x_25719;
wire x_25720;
wire x_25721;
wire x_25722;
wire x_25723;
wire x_25724;
wire x_25725;
wire x_25726;
wire x_25727;
wire x_25728;
wire x_25729;
wire x_25730;
wire x_25731;
wire x_25732;
wire x_25733;
wire x_25734;
wire x_25735;
wire x_25736;
wire x_25737;
wire x_25738;
wire x_25739;
wire x_25740;
wire x_25741;
wire x_25742;
wire x_25743;
wire x_25744;
wire x_25745;
wire x_25746;
wire x_25747;
wire x_25748;
wire x_25749;
wire x_25750;
wire x_25751;
wire x_25752;
wire x_25753;
wire x_25754;
wire x_25755;
wire x_25756;
wire x_25757;
wire x_25758;
wire x_25759;
wire x_25760;
wire x_25761;
wire x_25762;
wire x_25763;
wire x_25764;
wire x_25765;
wire x_25766;
wire x_25767;
wire x_25768;
wire x_25769;
wire x_25770;
wire x_25771;
wire x_25772;
wire x_25773;
wire x_25774;
wire x_25775;
wire x_25776;
wire x_25777;
wire x_25778;
wire x_25779;
wire x_25780;
wire x_25781;
wire x_25782;
wire x_25783;
wire x_25784;
wire x_25785;
wire x_25786;
wire x_25787;
wire x_25788;
wire x_25789;
wire x_25790;
wire x_25791;
wire x_25792;
wire x_25793;
wire x_25794;
wire x_25795;
wire x_25796;
wire x_25797;
wire x_25798;
wire x_25799;
wire x_25800;
wire x_25801;
wire x_25802;
wire x_25803;
wire x_25804;
wire x_25805;
wire x_25806;
wire x_25807;
wire x_25808;
wire x_25809;
wire x_25810;
wire x_25811;
wire x_25812;
wire x_25813;
wire x_25814;
wire x_25815;
wire x_25816;
wire x_25817;
wire x_25818;
wire x_25819;
wire x_25820;
wire x_25821;
wire x_25822;
wire x_25823;
wire x_25824;
wire x_25825;
wire x_25826;
wire x_25827;
wire x_25828;
wire x_25829;
wire x_25830;
wire x_25831;
wire x_25832;
wire x_25833;
wire x_25834;
wire x_25835;
wire x_25836;
wire x_25837;
wire x_25838;
wire x_25839;
wire x_25840;
wire x_25841;
wire x_25842;
wire x_25843;
wire x_25844;
wire x_25845;
wire x_25846;
wire x_25847;
wire x_25848;
wire x_25849;
wire x_25850;
wire x_25851;
wire x_25852;
wire x_25853;
wire x_25854;
wire x_25855;
wire x_25856;
wire x_25857;
wire x_25858;
wire x_25859;
wire x_25860;
wire x_25861;
wire x_25862;
wire x_25863;
wire x_25864;
wire x_25865;
wire x_25866;
wire x_25867;
wire x_25868;
wire x_25869;
wire x_25870;
wire x_25871;
wire x_25872;
wire x_25873;
wire x_25874;
wire x_25875;
wire x_25876;
wire x_25877;
wire x_25878;
wire x_25879;
wire x_25880;
wire x_25881;
wire x_25882;
wire x_25883;
wire x_25884;
wire x_25885;
wire x_25886;
wire x_25887;
wire x_25888;
wire x_25889;
wire x_25890;
wire x_25891;
wire x_25892;
wire x_25893;
wire x_25894;
wire x_25895;
wire x_25896;
wire x_25897;
wire x_25898;
wire x_25899;
wire x_25900;
wire x_25901;
wire x_25902;
wire x_25903;
wire x_25904;
wire x_25905;
wire x_25906;
wire x_25907;
wire x_25908;
wire x_25909;
wire x_25910;
wire x_25911;
wire x_25912;
wire x_25913;
wire x_25914;
wire x_25915;
wire x_25916;
wire x_25917;
wire x_25918;
wire x_25919;
wire x_25920;
wire x_25921;
wire x_25922;
wire x_25923;
wire x_25924;
wire x_25925;
wire x_25926;
wire x_25927;
wire x_25928;
wire x_25929;
wire x_25930;
wire x_25931;
wire x_25932;
wire x_25933;
wire x_25934;
wire x_25935;
wire x_25936;
wire x_25937;
wire x_25938;
wire x_25939;
wire x_25940;
wire x_25941;
wire x_25942;
wire x_25943;
wire x_25944;
wire x_25945;
wire x_25946;
wire x_25947;
wire x_25948;
wire x_25949;
wire x_25950;
wire x_25951;
wire x_25952;
wire x_25953;
wire x_25954;
wire x_25955;
wire x_25956;
wire x_25957;
wire x_25958;
wire x_25959;
wire x_25960;
wire x_25961;
wire x_25962;
wire x_25963;
wire x_25964;
wire x_25965;
wire x_25966;
wire x_25967;
wire x_25968;
wire x_25969;
wire x_25970;
wire x_25971;
wire x_25972;
wire x_25973;
wire x_25974;
wire x_25975;
wire x_25976;
wire x_25977;
wire x_25978;
wire x_25979;
wire x_25980;
wire x_25981;
wire x_25982;
wire x_25983;
wire x_25984;
wire x_25985;
wire x_25986;
wire x_25987;
wire x_25988;
wire x_25989;
wire x_25990;
wire x_25991;
wire x_25992;
wire x_25993;
wire x_25994;
wire x_25995;
wire x_25996;
wire x_25997;
wire x_25998;
wire x_25999;
wire x_26000;
wire x_26001;
wire x_26002;
wire x_26003;
wire x_26004;
wire x_26005;
wire x_26006;
wire x_26007;
wire x_26008;
wire x_26009;
wire x_26010;
wire x_26011;
wire x_26012;
wire x_26013;
wire x_26014;
wire x_26015;
wire x_26016;
wire x_26017;
wire x_26018;
wire x_26019;
wire x_26020;
wire x_26021;
wire x_26022;
wire x_26023;
wire x_26024;
wire x_26025;
wire x_26026;
wire x_26027;
wire x_26028;
wire x_26029;
wire x_26030;
wire x_26031;
wire x_26032;
wire x_26033;
wire x_26034;
wire x_26035;
wire x_26036;
wire x_26037;
wire x_26038;
wire x_26039;
wire x_26040;
wire x_26041;
wire x_26042;
wire x_26043;
wire x_26044;
wire x_26045;
wire x_26046;
wire x_26047;
wire x_26048;
wire x_26049;
wire x_26050;
wire x_26051;
wire x_26052;
wire x_26053;
wire x_26054;
wire x_26055;
wire x_26056;
wire x_26057;
wire x_26058;
wire x_26059;
wire x_26060;
wire x_26061;
wire x_26062;
wire x_26063;
wire x_26064;
wire x_26065;
wire x_26066;
wire x_26067;
wire x_26068;
wire x_26069;
wire x_26070;
wire x_26071;
wire x_26072;
wire x_26073;
wire x_26074;
wire x_26075;
wire x_26076;
wire x_26077;
wire x_26078;
wire x_26079;
wire x_26080;
wire x_26081;
wire x_26082;
wire x_26083;
wire x_26084;
wire x_26085;
wire x_26086;
wire x_26087;
wire x_26088;
wire x_26089;
wire x_26090;
wire x_26091;
wire x_26092;
wire x_26093;
wire x_26094;
wire x_26095;
wire x_26096;
wire x_26097;
wire x_26098;
wire x_26099;
wire x_26100;
wire x_26101;
wire x_26102;
wire x_26103;
wire x_26104;
wire x_26105;
wire x_26106;
wire x_26107;
wire x_26108;
wire x_26109;
wire x_26110;
wire x_26111;
wire x_26112;
wire x_26113;
wire x_26114;
wire x_26115;
wire x_26116;
wire x_26117;
wire x_26118;
wire x_26119;
wire x_26120;
wire x_26121;
wire x_26122;
wire x_26123;
wire x_26124;
wire x_26125;
wire x_26126;
wire x_26127;
wire x_26128;
wire x_26129;
wire x_26130;
wire x_26131;
wire x_26132;
wire x_26133;
wire x_26134;
wire x_26135;
wire x_26136;
wire x_26137;
wire x_26138;
wire x_26139;
wire x_26140;
wire x_26141;
wire x_26142;
wire x_26143;
wire x_26144;
wire x_26145;
wire x_26146;
wire x_26147;
wire x_26148;
wire x_26149;
wire x_26150;
wire x_26151;
wire x_26152;
wire x_26153;
wire x_26154;
wire x_26155;
wire x_26156;
wire x_26157;
wire x_26158;
wire x_26159;
wire x_26160;
wire x_26161;
wire x_26162;
wire x_26163;
wire x_26164;
wire x_26165;
wire x_26166;
wire x_26167;
wire x_26168;
wire x_26169;
wire x_26170;
wire x_26171;
wire x_26172;
wire x_26173;
wire x_26174;
wire x_26175;
wire x_26176;
wire x_26177;
wire x_26178;
wire x_26179;
wire x_26180;
wire x_26181;
wire x_26182;
wire x_26183;
wire x_26184;
wire x_26185;
wire x_26186;
wire x_26187;
wire x_26188;
wire x_26189;
wire x_26190;
wire x_26191;
wire x_26192;
wire x_26193;
wire x_26194;
wire x_26195;
wire x_26196;
wire x_26197;
wire x_26198;
wire x_26199;
wire x_26200;
wire x_26201;
wire x_26202;
wire x_26203;
wire x_26204;
wire x_26205;
wire x_26206;
wire x_26207;
wire x_26208;
wire x_26209;
wire x_26210;
wire x_26211;
wire x_26212;
wire x_26213;
wire x_26214;
wire x_26215;
wire x_26216;
wire x_26217;
wire x_26218;
wire x_26219;
wire x_26220;
wire x_26221;
wire x_26222;
wire x_26223;
wire x_26224;
wire x_26225;
wire x_26226;
wire x_26227;
wire x_26228;
wire x_26229;
wire x_26230;
wire x_26231;
wire x_26232;
wire x_26233;
wire x_26234;
wire x_26235;
wire x_26236;
wire x_26237;
wire x_26238;
wire x_26239;
wire x_26240;
wire x_26241;
wire x_26242;
wire x_26243;
wire x_26244;
wire x_26245;
wire x_26246;
wire x_26247;
wire x_26248;
wire x_26249;
wire x_26250;
wire x_26251;
wire x_26252;
wire x_26253;
wire x_26254;
wire x_26255;
wire x_26256;
wire x_26257;
wire x_26258;
wire x_26259;
wire x_26260;
wire x_26261;
wire x_26262;
wire x_26263;
wire x_26264;
wire x_26265;
wire x_26266;
wire x_26267;
wire x_26268;
wire x_26269;
wire x_26270;
wire x_26271;
wire x_26272;
wire x_26273;
wire x_26274;
wire x_26275;
wire x_26276;
wire x_26277;
wire x_26278;
wire x_26279;
wire x_26280;
wire x_26281;
wire x_26282;
wire x_26283;
wire x_26284;
wire x_26285;
wire x_26286;
wire x_26287;
wire x_26288;
wire x_26289;
wire x_26290;
wire x_26291;
wire x_26292;
wire x_26293;
wire x_26294;
wire x_26295;
wire x_26296;
wire x_26297;
wire x_26298;
wire x_26299;
wire x_26300;
wire x_26301;
wire x_26302;
wire x_26303;
wire x_26304;
wire x_26305;
wire x_26306;
wire x_26307;
wire x_26308;
wire x_26309;
wire x_26310;
wire x_26311;
wire x_26312;
wire x_26313;
wire x_26314;
wire x_26315;
wire x_26316;
wire x_26317;
wire x_26318;
wire x_26319;
wire x_26320;
wire x_26321;
wire x_26322;
wire x_26323;
wire x_26324;
wire x_26325;
wire x_26326;
wire x_26327;
wire x_26328;
wire x_26329;
wire x_26330;
wire x_26331;
wire x_26332;
wire x_26333;
wire x_26334;
wire x_26335;
wire x_26336;
wire x_26337;
wire x_26338;
wire x_26339;
wire x_26340;
wire x_26341;
wire x_26342;
wire x_26343;
wire x_26344;
wire x_26345;
wire x_26346;
wire x_26347;
wire x_26348;
wire x_26349;
wire x_26350;
wire x_26351;
wire x_26352;
wire x_26353;
wire x_26354;
wire x_26355;
wire x_26356;
wire x_26357;
wire x_26358;
wire x_26359;
wire x_26360;
wire x_26361;
wire x_26362;
wire x_26363;
wire x_26364;
wire x_26365;
wire x_26366;
wire x_26367;
wire x_26368;
wire x_26369;
wire x_26370;
wire x_26371;
wire x_26372;
wire x_26373;
wire x_26374;
wire x_26375;
wire x_26376;
wire x_26377;
wire x_26378;
wire x_26379;
wire x_26380;
wire x_26381;
wire x_26382;
wire x_26383;
wire x_26384;
wire x_26385;
wire x_26386;
wire x_26387;
wire x_26388;
wire x_26389;
wire x_26390;
wire x_26391;
wire x_26392;
wire x_26393;
wire x_26394;
wire x_26395;
wire x_26396;
wire x_26397;
wire x_26398;
wire x_26399;
wire x_26400;
wire x_26401;
wire x_26402;
wire x_26403;
wire x_26404;
wire x_26405;
wire x_26406;
wire x_26407;
wire x_26408;
wire x_26409;
wire x_26410;
wire x_26411;
wire x_26412;
wire x_26413;
wire x_26414;
wire x_26415;
wire x_26416;
wire x_26417;
wire x_26418;
wire x_26419;
wire x_26420;
wire x_26421;
wire x_26422;
wire x_26423;
wire x_26424;
wire x_26425;
wire x_26426;
wire x_26427;
wire x_26428;
wire x_26429;
wire x_26430;
wire x_26431;
wire x_26432;
wire x_26433;
wire x_26434;
wire x_26435;
wire x_26436;
wire x_26437;
wire x_26438;
wire x_26439;
wire x_26440;
wire x_26441;
wire x_26442;
wire x_26443;
wire x_26444;
wire x_26445;
wire x_26446;
wire x_26447;
wire x_26448;
wire x_26449;
wire x_26450;
wire x_26451;
wire x_26452;
wire x_26453;
wire x_26454;
wire x_26455;
wire x_26456;
wire x_26457;
wire x_26458;
wire x_26459;
wire x_26460;
wire x_26461;
wire x_26462;
wire x_26463;
wire x_26464;
wire x_26465;
wire x_26466;
wire x_26467;
wire x_26468;
wire x_26469;
wire x_26470;
wire x_26471;
wire x_26472;
wire x_26473;
wire x_26474;
wire x_26475;
wire x_26476;
wire x_26477;
wire x_26478;
wire x_26479;
wire x_26480;
wire x_26481;
wire x_26482;
wire x_26483;
wire x_26484;
wire x_26485;
wire x_26486;
wire x_26487;
wire x_26488;
wire x_26489;
wire x_26490;
wire x_26491;
wire x_26492;
wire x_26493;
wire x_26494;
wire x_26495;
wire x_26496;
wire x_26497;
wire x_26498;
wire x_26499;
wire x_26500;
wire x_26501;
wire x_26502;
wire x_26503;
wire x_26504;
wire x_26505;
wire x_26506;
wire x_26507;
wire x_26508;
wire x_26509;
wire x_26510;
wire x_26511;
wire x_26512;
wire x_26513;
wire x_26514;
wire x_26515;
wire x_26516;
wire x_26517;
wire x_26518;
wire x_26519;
wire x_26520;
wire x_26521;
wire x_26522;
wire x_26523;
wire x_26524;
wire x_26525;
wire x_26526;
wire x_26527;
wire x_26528;
wire x_26529;
wire x_26530;
wire x_26531;
wire x_26532;
wire x_26533;
wire x_26534;
wire x_26535;
wire x_26536;
wire x_26537;
wire x_26538;
wire x_26539;
wire x_26540;
wire x_26541;
wire x_26542;
wire x_26543;
wire x_26544;
wire x_26545;
wire x_26546;
wire x_26547;
wire x_26548;
wire x_26549;
wire x_26550;
wire x_26551;
wire x_26552;
wire x_26553;
wire x_26554;
wire x_26555;
wire x_26556;
wire x_26557;
wire x_26558;
wire x_26559;
wire x_26560;
wire x_26561;
wire x_26562;
wire x_26563;
wire x_26564;
wire x_26565;
wire x_26566;
wire x_26567;
wire x_26568;
wire x_26569;
wire x_26570;
wire x_26571;
wire x_26572;
wire x_26573;
wire x_26574;
wire x_26575;
wire x_26576;
wire x_26577;
wire x_26578;
wire x_26579;
wire x_26580;
wire x_26581;
wire x_26582;
wire x_26583;
wire x_26584;
wire x_26585;
wire x_26586;
wire x_26587;
wire x_26588;
wire x_26589;
wire x_26590;
wire x_26591;
wire x_26592;
wire x_26593;
wire x_26594;
wire x_26595;
wire x_26596;
wire x_26597;
wire x_26598;
wire x_26599;
wire x_26600;
wire x_26601;
wire x_26602;
wire x_26603;
wire x_26604;
wire x_26605;
wire x_26606;
wire x_26607;
wire x_26608;
wire x_26609;
wire x_26610;
wire x_26611;
wire x_26612;
wire x_26613;
wire x_26614;
wire x_26615;
wire x_26616;
wire x_26617;
wire x_26618;
wire x_26619;
wire x_26620;
wire x_26621;
wire x_26622;
wire x_26623;
wire x_26624;
wire x_26625;
wire x_26626;
wire x_26627;
wire x_26628;
wire x_26629;
wire x_26630;
wire x_26631;
wire x_26632;
wire x_26633;
wire x_26634;
wire x_26635;
wire x_26636;
wire x_26637;
wire x_26638;
wire x_26639;
wire x_26640;
wire x_26641;
wire x_26642;
wire x_26643;
wire x_26644;
wire x_26645;
wire x_26646;
wire x_26647;
wire x_26648;
wire x_26649;
wire x_26650;
wire x_26651;
wire x_26652;
wire x_26653;
wire x_26654;
wire x_26655;
wire x_26656;
wire x_26657;
wire x_26658;
wire x_26659;
wire x_26660;
wire x_26661;
wire x_26662;
wire x_26663;
wire x_26664;
wire x_26665;
wire x_26666;
wire x_26667;
wire x_26668;
wire x_26669;
wire x_26670;
wire x_26671;
wire x_26672;
wire x_26673;
wire x_26674;
wire x_26675;
wire x_26676;
wire x_26677;
wire x_26678;
wire x_26679;
wire x_26680;
wire x_26681;
wire x_26682;
wire x_26683;
wire x_26684;
wire x_26685;
wire x_26686;
wire x_26687;
wire x_26688;
wire x_26689;
wire x_26690;
wire x_26691;
wire x_26692;
wire x_26693;
wire x_26694;
wire x_26695;
wire x_26696;
wire x_26697;
wire x_26698;
wire x_26699;
wire x_26700;
wire x_26701;
wire x_26702;
wire x_26703;
wire x_26704;
wire x_26705;
wire x_26706;
wire x_26707;
wire x_26708;
wire x_26709;
wire x_26710;
wire x_26711;
wire x_26712;
wire x_26713;
wire x_26714;
wire x_26715;
wire x_26716;
wire x_26717;
wire x_26718;
wire x_26719;
wire x_26720;
wire x_26721;
wire x_26722;
wire x_26723;
wire x_26724;
wire x_26725;
wire x_26726;
wire x_26727;
wire x_26728;
wire x_26729;
wire x_26730;
wire x_26731;
wire x_26732;
wire x_26733;
wire x_26734;
wire x_26735;
wire x_26736;
wire x_26737;
wire x_26738;
wire x_26739;
wire x_26740;
wire x_26741;
wire x_26742;
wire x_26743;
wire x_26744;
wire x_26745;
wire x_26746;
wire x_26747;
wire x_26748;
wire x_26749;
wire x_26750;
wire x_26751;
wire x_26752;
wire x_26753;
wire x_26754;
wire x_26755;
wire x_26756;
wire x_26757;
wire x_26758;
wire x_26759;
wire x_26760;
wire x_26761;
wire x_26762;
wire x_26763;
wire x_26764;
wire x_26765;
wire x_26766;
wire x_26767;
wire x_26768;
wire x_26769;
wire x_26770;
wire x_26771;
wire x_26772;
wire x_26773;
wire x_26774;
wire x_26775;
wire x_26776;
wire x_26777;
wire x_26778;
wire x_26779;
wire x_26780;
wire x_26781;
wire x_26782;
wire x_26783;
wire x_26784;
wire x_26785;
wire x_26786;
wire x_26787;
wire x_26788;
wire x_26789;
wire x_26790;
wire x_26791;
wire x_26792;
wire x_26793;
wire x_26794;
wire x_26795;
wire x_26796;
wire x_26797;
wire x_26798;
wire x_26799;
wire x_26800;
wire x_26801;
wire x_26802;
wire x_26803;
wire x_26804;
wire x_26805;
wire x_26806;
wire x_26807;
wire x_26808;
wire x_26809;
wire x_26810;
wire x_26811;
wire x_26812;
wire x_26813;
wire x_26814;
wire x_26815;
wire x_26816;
wire x_26817;
wire x_26818;
wire x_26819;
wire x_26820;
wire x_26821;
wire x_26822;
wire x_26823;
wire x_26824;
wire x_26825;
wire x_26826;
wire x_26827;
wire x_26828;
wire x_26829;
wire x_26830;
wire x_26831;
wire x_26832;
wire x_26833;
wire x_26834;
wire x_26835;
wire x_26836;
wire x_26837;
wire x_26838;
wire x_26839;
wire x_26840;
wire x_26841;
wire x_26842;
wire x_26843;
wire x_26844;
wire x_26845;
wire x_26846;
wire x_26847;
wire x_26848;
wire x_26849;
wire x_26850;
wire x_26851;
wire x_26852;
wire x_26853;
wire x_26854;
wire x_26855;
wire x_26856;
wire x_26857;
wire x_26858;
wire x_26859;
wire x_26860;
wire x_26861;
wire x_26862;
wire x_26863;
wire x_26864;
wire x_26865;
wire x_26866;
wire x_26867;
wire x_26868;
wire x_26869;
wire x_26870;
wire x_26871;
wire x_26872;
wire x_26873;
wire x_26874;
wire x_26875;
wire x_26876;
wire x_26877;
wire x_26878;
wire x_26879;
wire x_26880;
wire x_26881;
wire x_26882;
wire x_26883;
wire x_26884;
wire x_26885;
wire x_26886;
wire x_26887;
wire x_26888;
wire x_26889;
wire x_26890;
wire x_26891;
wire x_26892;
wire x_26893;
wire x_26894;
wire x_26895;
wire x_26896;
wire x_26897;
wire x_26898;
wire x_26899;
wire x_26900;
wire x_26901;
wire x_26902;
wire x_26903;
wire x_26904;
wire x_26905;
wire x_26906;
wire x_26907;
wire x_26908;
wire x_26909;
wire x_26910;
wire x_26911;
wire x_26912;
wire x_26913;
wire x_26914;
wire x_26915;
wire x_26916;
wire x_26917;
wire x_26918;
wire x_26919;
wire x_26920;
wire x_26921;
wire x_26922;
wire x_26923;
wire x_26924;
wire x_26925;
wire x_26926;
wire x_26927;
wire x_26928;
wire x_26929;
wire x_26930;
wire x_26931;
wire x_26932;
wire x_26933;
wire x_26934;
wire x_26935;
wire x_26936;
wire x_26937;
wire x_26938;
wire x_26939;
wire x_26940;
wire x_26941;
wire x_26942;
wire x_26943;
wire x_26944;
wire x_26945;
wire x_26946;
wire x_26947;
wire x_26948;
wire x_26949;
wire x_26950;
wire x_26951;
wire x_26952;
wire x_26953;
wire x_26954;
wire x_26955;
wire x_26956;
wire x_26957;
wire x_26958;
wire x_26959;
wire x_26960;
wire x_26961;
wire x_26962;
wire x_26963;
wire x_26964;
wire x_26965;
wire x_26966;
wire x_26967;
wire x_26968;
wire x_26969;
wire x_26970;
wire x_26971;
wire x_26972;
wire x_26973;
wire x_26974;
wire x_26975;
wire x_26976;
wire x_26977;
wire x_26978;
wire x_26979;
wire x_26980;
wire x_26981;
wire x_26982;
wire x_26983;
wire x_26984;
wire x_26985;
wire x_26986;
wire x_26987;
wire x_26988;
wire x_26989;
wire x_26990;
wire x_26991;
wire x_26992;
wire x_26993;
wire x_26994;
wire x_26995;
wire x_26996;
wire x_26997;
wire x_26998;
wire x_26999;
wire x_27000;
wire x_27001;
wire x_27002;
wire x_27003;
wire x_27004;
wire x_27005;
wire x_27006;
wire x_27007;
wire x_27008;
wire x_27009;
wire x_27010;
wire x_27011;
wire x_27012;
wire x_27013;
wire x_27014;
wire x_27015;
wire x_27016;
wire x_27017;
wire x_27018;
wire x_27019;
wire x_27020;
wire x_27021;
wire x_27022;
wire x_27023;
wire x_27024;
wire x_27025;
wire x_27026;
wire x_27027;
wire x_27028;
wire x_27029;
wire x_27030;
wire x_27031;
wire x_27032;
wire x_27033;
wire x_27034;
wire x_27035;
wire x_27036;
wire x_27037;
wire x_27038;
wire x_27039;
wire x_27040;
wire x_27041;
wire x_27042;
wire x_27043;
wire x_27044;
wire x_27045;
wire x_27046;
wire x_27047;
wire x_27048;
wire x_27049;
wire x_27050;
wire x_27051;
wire x_27052;
wire x_27053;
wire x_27054;
wire x_27055;
wire x_27056;
wire x_27057;
wire x_27058;
wire x_27059;
wire x_27060;
wire x_27061;
wire x_27062;
wire x_27063;
wire x_27064;
wire x_27065;
wire x_27066;
wire x_27067;
wire x_27068;
wire x_27069;
wire x_27070;
wire x_27071;
wire x_27072;
wire x_27073;
wire x_27074;
wire x_27075;
wire x_27076;
wire x_27077;
wire x_27078;
wire x_27079;
wire x_27080;
wire x_27081;
wire x_27082;
wire x_27083;
wire x_27084;
wire x_27085;
wire x_27086;
wire x_27087;
wire x_27088;
wire x_27089;
wire x_27090;
wire x_27091;
wire x_27092;
wire x_27093;
wire x_27094;
wire x_27095;
wire x_27096;
wire x_27097;
wire x_27098;
wire x_27099;
wire x_27100;
wire x_27101;
wire x_27102;
wire x_27103;
wire x_27104;
wire x_27105;
wire x_27106;
wire x_27107;
wire x_27108;
wire x_27109;
wire x_27110;
wire x_27111;
wire x_27112;
wire x_27113;
wire x_27114;
wire x_27115;
wire x_27116;
wire x_27117;
wire x_27118;
wire x_27119;
wire x_27120;
wire x_27121;
wire x_27122;
wire x_27123;
wire x_27124;
wire x_27125;
wire x_27126;
wire x_27127;
wire x_27128;
wire x_27129;
wire x_27130;
wire x_27131;
wire x_27132;
wire x_27133;
wire x_27134;
wire x_27135;
wire x_27136;
wire x_27137;
wire x_27138;
wire x_27139;
wire x_27140;
wire x_27141;
wire x_27142;
wire x_27143;
wire x_27144;
wire x_27145;
wire x_27146;
wire x_27147;
wire x_27148;
wire x_27149;
wire x_27150;
wire x_27151;
wire x_27152;
wire x_27153;
wire x_27154;
wire x_27155;
wire x_27156;
wire x_27157;
wire x_27158;
wire x_27159;
wire x_27160;
wire x_27161;
wire x_27162;
wire x_27163;
wire x_27164;
wire x_27165;
wire x_27166;
wire x_27167;
wire x_27168;
wire x_27169;
wire x_27170;
wire x_27171;
wire x_27172;
wire x_27173;
wire x_27174;
wire x_27175;
wire x_27176;
wire x_27177;
wire x_27178;
wire x_27179;
wire x_27180;
wire x_27181;
wire x_27182;
wire x_27183;
wire x_27184;
wire x_27185;
wire x_27186;
wire x_27187;
wire x_27188;
wire x_27189;
wire x_27190;
wire x_27191;
wire x_27192;
wire x_27193;
wire x_27194;
wire x_27195;
wire x_27196;
wire x_27197;
wire x_27198;
wire x_27199;
wire x_27200;
wire x_27201;
wire x_27202;
wire x_27203;
wire x_27204;
wire x_27205;
wire x_27206;
wire x_27207;
wire x_27208;
wire x_27209;
wire x_27210;
wire x_27211;
wire x_27212;
wire x_27213;
wire x_27214;
wire x_27215;
wire x_27216;
wire x_27217;
wire x_27218;
wire x_27219;
wire x_27220;
wire x_27221;
wire x_27222;
wire x_27223;
wire x_27224;
wire x_27225;
wire x_27226;
wire x_27227;
wire x_27228;
wire x_27229;
wire x_27230;
wire x_27231;
wire x_27232;
wire x_27233;
wire x_27234;
wire x_27235;
wire x_27236;
wire x_27237;
wire x_27238;
wire x_27239;
wire x_27240;
wire x_27241;
wire x_27242;
wire x_27243;
wire x_27244;
wire x_27245;
wire x_27246;
wire x_27247;
wire x_27248;
wire x_27249;
wire x_27250;
wire x_27251;
wire x_27252;
wire x_27253;
wire x_27254;
wire x_27255;
wire x_27256;
wire x_27257;
wire x_27258;
wire x_27259;
wire x_27260;
wire x_27261;
wire x_27262;
wire x_27263;
wire x_27264;
wire x_27265;
wire x_27266;
wire x_27267;
wire x_27268;
wire x_27269;
wire x_27270;
wire x_27271;
wire x_27272;
wire x_27273;
wire x_27274;
wire x_27275;
wire x_27276;
wire x_27277;
wire x_27278;
wire x_27279;
wire x_27280;
wire x_27281;
wire x_27282;
wire x_27283;
wire x_27284;
wire x_27285;
wire x_27286;
wire x_27287;
wire x_27288;
wire x_27289;
wire x_27290;
wire x_27291;
wire x_27292;
wire x_27293;
wire x_27294;
wire x_27295;
wire x_27296;
wire x_27297;
wire x_27298;
wire x_27299;
wire x_27300;
wire x_27301;
wire x_27302;
wire x_27303;
wire x_27304;
wire x_27305;
wire x_27306;
wire x_27307;
wire x_27308;
wire x_27309;
wire x_27310;
wire x_27311;
wire x_27312;
wire x_27313;
wire x_27314;
wire x_27315;
wire x_27316;
wire x_27317;
wire x_27318;
wire x_27319;
wire x_27320;
wire x_27321;
wire x_27322;
wire x_27323;
wire x_27324;
wire x_27325;
wire x_27326;
wire x_27327;
wire x_27328;
wire x_27329;
wire x_27330;
wire x_27331;
wire x_27332;
wire x_27333;
wire x_27334;
wire x_27335;
wire x_27336;
wire x_27337;
wire x_27338;
wire x_27339;
wire x_27340;
wire x_27341;
wire x_27342;
wire x_27343;
wire x_27344;
wire x_27345;
wire x_27346;
wire x_27347;
wire x_27348;
wire x_27349;
wire x_27350;
wire x_27351;
wire x_27352;
wire x_27353;
wire x_27354;
wire x_27355;
wire x_27356;
wire x_27357;
wire x_27358;
wire x_27359;
wire x_27360;
wire x_27361;
wire x_27362;
wire x_27363;
wire x_27364;
wire x_27365;
wire x_27366;
wire x_27367;
wire x_27368;
wire x_27369;
wire x_27370;
wire x_27371;
wire x_27372;
wire x_27373;
wire x_27374;
wire x_27375;
wire x_27376;
wire x_27377;
wire x_27378;
wire x_27379;
wire x_27380;
wire x_27381;
wire x_27382;
wire x_27383;
wire x_27384;
wire x_27385;
wire x_27386;
wire x_27387;
wire x_27388;
wire x_27389;
wire x_27390;
wire x_27391;
wire x_27392;
wire x_27393;
wire x_27394;
wire x_27395;
wire x_27396;
wire x_27397;
wire x_27398;
wire x_27399;
wire x_27400;
wire x_27401;
wire x_27402;
wire x_27403;
wire x_27404;
wire x_27405;
wire x_27406;
wire x_27407;
wire x_27408;
wire x_27409;
wire x_27410;
wire x_27411;
wire x_27412;
wire x_27413;
wire x_27414;
wire x_27415;
wire x_27416;
wire x_27417;
wire x_27418;
wire x_27419;
wire x_27420;
wire x_27421;
wire x_27422;
wire x_27423;
wire x_27424;
wire x_27425;
wire x_27426;
wire x_27427;
wire x_27428;
wire x_27429;
wire x_27430;
wire x_27431;
wire x_27432;
wire x_27433;
wire x_27434;
wire x_27435;
wire x_27436;
wire x_27437;
wire x_27438;
wire x_27439;
wire x_27440;
wire x_27441;
wire x_27442;
wire x_27443;
wire x_27444;
wire x_27445;
wire x_27446;
wire x_27447;
wire x_27448;
wire x_27449;
wire x_27450;
wire x_27451;
wire x_27452;
wire x_27453;
wire x_27454;
wire x_27455;
wire x_27456;
wire x_27457;
wire x_27458;
wire x_27459;
wire x_27460;
wire x_27461;
wire x_27462;
wire x_27463;
wire x_27464;
wire x_27465;
wire x_27466;
wire x_27467;
wire x_27468;
wire x_27469;
wire x_27470;
wire x_27471;
wire x_27472;
wire x_27473;
wire x_27474;
wire x_27475;
wire x_27476;
wire x_27477;
wire x_27478;
wire x_27479;
wire x_27480;
wire x_27481;
wire x_27482;
wire x_27483;
wire x_27484;
wire x_27485;
wire x_27486;
wire x_27487;
wire x_27488;
wire x_27489;
wire x_27490;
wire x_27491;
wire x_27492;
wire x_27493;
wire x_27494;
wire x_27495;
wire x_27496;
wire x_27497;
wire x_27498;
wire x_27499;
wire x_27500;
wire x_27501;
wire x_27502;
wire x_27503;
wire x_27504;
wire x_27505;
wire x_27506;
wire x_27507;
wire x_27508;
wire x_27509;
wire x_27510;
wire x_27511;
wire x_27512;
wire x_27513;
wire x_27514;
wire x_27515;
wire x_27516;
wire x_27517;
wire x_27518;
wire x_27519;
wire x_27520;
wire x_27521;
wire x_27522;
wire x_27523;
wire x_27524;
wire x_27525;
wire x_27526;
wire x_27527;
wire x_27528;
wire x_27529;
wire x_27530;
wire x_27531;
wire x_27532;
wire x_27533;
wire x_27534;
wire x_27535;
wire x_27536;
wire x_27537;
wire x_27538;
wire x_27539;
wire x_27540;
wire x_27541;
wire x_27542;
wire x_27543;
wire x_27544;
wire x_27545;
wire x_27546;
wire x_27547;
wire x_27548;
wire x_27549;
wire x_27550;
wire x_27551;
wire x_27552;
wire x_27553;
wire x_27554;
wire x_27555;
wire x_27556;
wire x_27557;
wire x_27558;
wire x_27559;
wire x_27560;
wire x_27561;
wire x_27562;
wire x_27563;
wire x_27564;
wire x_27565;
wire x_27566;
wire x_27567;
wire x_27568;
wire x_27569;
wire x_27570;
wire x_27571;
wire x_27572;
wire x_27573;
wire x_27574;
wire x_27575;
wire x_27576;
wire x_27577;
wire x_27578;
wire x_27579;
wire x_27580;
wire x_27581;
wire x_27582;
wire x_27583;
wire x_27584;
wire x_27585;
wire x_27586;
wire x_27587;
wire x_27588;
wire x_27589;
wire x_27590;
wire x_27591;
wire x_27592;
wire x_27593;
wire x_27594;
wire x_27595;
wire x_27596;
wire x_27597;
wire x_27598;
wire x_27599;
wire x_27600;
wire x_27601;
wire x_27602;
wire x_27603;
wire x_27604;
wire x_27605;
wire x_27606;
wire x_27607;
wire x_27608;
wire x_27609;
wire x_27610;
wire x_27611;
wire x_27612;
wire x_27613;
wire x_27614;
wire x_27615;
wire x_27616;
wire x_27617;
wire x_27618;
wire x_27619;
wire x_27620;
wire x_27621;
wire x_27622;
wire x_27623;
wire x_27624;
wire x_27625;
wire x_27626;
wire x_27627;
wire x_27628;
wire x_27629;
wire x_27630;
wire x_27631;
wire x_27632;
wire x_27633;
wire x_27634;
wire x_27635;
wire x_27636;
wire x_27637;
wire x_27638;
wire x_27639;
wire x_27640;
wire x_27641;
wire x_27642;
wire x_27643;
wire x_27644;
wire x_27645;
wire x_27646;
wire x_27647;
wire x_27648;
wire x_27649;
wire x_27650;
wire x_27651;
wire x_27652;
wire x_27653;
wire x_27654;
wire x_27655;
wire x_27656;
wire x_27657;
wire x_27658;
wire x_27659;
wire x_27660;
wire x_27661;
wire x_27662;
wire x_27663;
wire x_27664;
wire x_27665;
wire x_27666;
wire x_27667;
wire x_27668;
wire x_27669;
wire x_27670;
wire x_27671;
wire x_27672;
wire x_27673;
wire x_27674;
wire x_27675;
wire x_27676;
wire x_27677;
wire x_27678;
wire x_27679;
wire x_27680;
wire x_27681;
wire x_27682;
wire x_27683;
wire x_27684;
wire x_27685;
wire x_27686;
wire x_27687;
wire x_27688;
wire x_27689;
wire x_27690;
wire x_27691;
wire x_27692;
wire x_27693;
wire x_27694;
wire x_27695;
wire x_27696;
wire x_27697;
wire x_27698;
wire x_27699;
wire x_27700;
wire x_27701;
wire x_27702;
wire x_27703;
wire x_27704;
wire x_27705;
wire x_27706;
wire x_27707;
wire x_27708;
wire x_27709;
wire x_27710;
wire x_27711;
wire x_27712;
wire x_27713;
wire x_27714;
wire x_27715;
wire x_27716;
wire x_27717;
wire x_27718;
wire x_27719;
wire x_27720;
wire x_27721;
wire x_27722;
wire x_27723;
wire x_27724;
wire x_27725;
wire x_27726;
wire x_27727;
wire x_27728;
wire x_27729;
wire x_27730;
wire x_27731;
wire x_27732;
wire x_27733;
wire x_27734;
wire x_27735;
wire x_27736;
wire x_27737;
wire x_27738;
wire x_27739;
wire x_27740;
wire x_27741;
wire x_27742;
wire x_27743;
wire x_27744;
wire x_27745;
wire x_27746;
wire x_27747;
wire x_27748;
wire x_27749;
wire x_27750;
wire x_27751;
wire x_27752;
wire x_27753;
wire x_27754;
wire x_27755;
wire x_27756;
wire x_27757;
wire x_27758;
wire x_27759;
wire x_27760;
wire x_27761;
wire x_27762;
wire x_27763;
wire x_27764;
wire x_27765;
wire x_27766;
wire x_27767;
wire x_27768;
wire x_27769;
wire x_27770;
wire x_27771;
wire x_27772;
wire x_27773;
wire x_27774;
wire x_27775;
wire x_27776;
wire x_27777;
wire x_27778;
wire x_27779;
wire x_27780;
wire x_27781;
wire x_27782;
wire x_27783;
wire x_27784;
wire x_27785;
wire x_27786;
wire x_27787;
wire x_27788;
wire x_27789;
wire x_27790;
wire x_27791;
wire x_27792;
wire x_27793;
wire x_27794;
wire x_27795;
wire x_27796;
wire x_27797;
wire x_27798;
wire x_27799;
wire x_27800;
wire x_27801;
wire x_27802;
wire x_27803;
wire x_27804;
wire x_27805;
wire x_27806;
wire x_27807;
wire x_27808;
wire x_27809;
wire x_27810;
wire x_27811;
wire x_27812;
wire x_27813;
wire x_27814;
wire x_27815;
wire x_27816;
wire x_27817;
wire x_27818;
wire x_27819;
wire x_27820;
wire x_27821;
wire x_27822;
wire x_27823;
wire x_27824;
wire x_27825;
wire x_27826;
wire x_27827;
wire x_27828;
wire x_27829;
wire x_27830;
wire x_27831;
wire x_27832;
wire x_27833;
wire x_27834;
wire x_27835;
wire x_27836;
wire x_27837;
wire x_27838;
wire x_27839;
wire x_27840;
wire x_27841;
wire x_27842;
wire x_27843;
wire x_27844;
wire x_27845;
wire x_27846;
wire x_27847;
wire x_27848;
wire x_27849;
wire x_27850;
wire x_27851;
wire x_27852;
wire x_27853;
wire x_27854;
wire x_27855;
wire x_27856;
wire x_27857;
wire x_27858;
wire x_27859;
wire x_27860;
wire x_27861;
wire x_27862;
wire x_27863;
wire x_27864;
wire x_27865;
wire x_27866;
wire x_27867;
wire x_27868;
wire x_27869;
wire x_27870;
wire x_27871;
wire x_27872;
wire x_27873;
wire x_27874;
wire x_27875;
wire x_27876;
wire x_27877;
wire x_27878;
wire x_27879;
wire x_27880;
wire x_27881;
wire x_27882;
wire x_27883;
wire x_27884;
wire x_27885;
wire x_27886;
wire x_27887;
wire x_27888;
wire x_27889;
wire x_27890;
wire x_27891;
wire x_27892;
wire x_27893;
wire x_27894;
wire x_27895;
wire x_27896;
wire x_27897;
wire x_27898;
wire x_27899;
wire x_27900;
wire x_27901;
wire x_27902;
wire x_27903;
wire x_27904;
wire x_27905;
wire x_27906;
wire x_27907;
wire x_27908;
wire x_27909;
wire x_27910;
wire x_27911;
wire x_27912;
wire x_27913;
wire x_27914;
wire x_27915;
wire x_27916;
wire x_27917;
wire x_27918;
wire x_27919;
wire x_27920;
wire x_27921;
wire x_27922;
wire x_27923;
wire x_27924;
wire x_27925;
wire x_27926;
wire x_27927;
wire x_27928;
wire x_27929;
wire x_27930;
wire x_27931;
wire x_27932;
wire x_27933;
wire x_27934;
wire x_27935;
wire x_27936;
wire x_27937;
wire x_27938;
wire x_27939;
wire x_27940;
wire x_27941;
wire x_27942;
wire x_27943;
wire x_27944;
wire x_27945;
wire x_27946;
wire x_27947;
wire x_27948;
wire x_27949;
wire x_27950;
wire x_27951;
wire x_27952;
wire x_27953;
wire x_27954;
wire x_27955;
wire x_27956;
wire x_27957;
wire x_27958;
wire x_27959;
wire x_27960;
wire x_27961;
wire x_27962;
wire x_27963;
wire x_27964;
wire x_27965;
wire x_27966;
wire x_27967;
wire x_27968;
wire x_27969;
wire x_27970;
wire x_27971;
wire x_27972;
wire x_27973;
wire x_27974;
wire x_27975;
wire x_27976;
wire x_27977;
wire x_27978;
wire x_27979;
wire x_27980;
wire x_27981;
wire x_27982;
wire x_27983;
wire x_27984;
wire x_27985;
wire x_27986;
wire x_27987;
wire x_27988;
wire x_27989;
wire x_27990;
wire x_27991;
wire x_27992;
wire x_27993;
wire x_27994;
wire x_27995;
wire x_27996;
wire x_27997;
wire x_27998;
wire x_27999;
wire x_28000;
wire x_28001;
wire x_28002;
wire x_28003;
wire x_28004;
wire x_28005;
wire x_28006;
wire x_28007;
wire x_28008;
wire x_28009;
wire x_28010;
wire x_28011;
wire x_28012;
wire x_28013;
wire x_28014;
wire x_28015;
wire x_28016;
wire x_28017;
wire x_28018;
wire x_28019;
wire x_28020;
wire x_28021;
wire x_28022;
wire x_28023;
wire x_28024;
wire x_28025;
wire x_28026;
wire x_28027;
wire x_28028;
wire x_28029;
wire x_28030;
wire x_28031;
wire x_28032;
wire x_28033;
wire x_28034;
wire x_28035;
wire x_28036;
wire x_28037;
wire x_28038;
wire x_28039;
wire x_28040;
wire x_28041;
wire x_28042;
wire x_28043;
wire x_28044;
wire x_28045;
wire x_28046;
wire x_28047;
wire x_28048;
wire x_28049;
wire x_28050;
wire x_28051;
wire x_28052;
wire x_28053;
wire x_28054;
wire x_28055;
wire x_28056;
wire x_28057;
wire x_28058;
wire x_28059;
wire x_28060;
wire x_28061;
wire x_28062;
wire x_28063;
wire x_28064;
wire x_28065;
wire x_28066;
wire x_28067;
wire x_28068;
wire x_28069;
wire x_28070;
wire x_28071;
wire x_28072;
wire x_28073;
wire x_28074;
wire x_28075;
wire x_28076;
wire x_28077;
wire x_28078;
wire x_28079;
wire x_28080;
wire x_28081;
wire x_28082;
wire x_28083;
wire x_28084;
wire x_28085;
wire x_28086;
wire x_28087;
wire x_28088;
wire x_28089;
wire x_28090;
wire x_28091;
wire x_28092;
wire x_28093;
wire x_28094;
wire x_28095;
wire x_28096;
wire x_28097;
wire x_28098;
wire x_28099;
wire x_28100;
wire x_28101;
wire x_28102;
wire x_28103;
wire x_28104;
wire x_28105;
wire x_28106;
wire x_28107;
wire x_28108;
wire x_28109;
wire x_28110;
wire x_28111;
wire x_28112;
wire x_28113;
wire x_28114;
wire x_28115;
wire x_28116;
wire x_28117;
wire x_28118;
wire x_28119;
wire x_28120;
wire x_28121;
wire x_28122;
wire x_28123;
wire x_28124;
wire x_28125;
wire x_28126;
wire x_28127;
wire x_28128;
wire x_28129;
wire x_28130;
wire x_28131;
wire x_28132;
wire x_28133;
wire x_28134;
wire x_28135;
wire x_28136;
wire x_28137;
wire x_28138;
wire x_28139;
wire x_28140;
wire x_28141;
wire x_28142;
wire x_28143;
wire x_28144;
wire x_28145;
wire x_28146;
wire x_28147;
wire x_28148;
wire x_28149;
wire x_28150;
wire x_28151;
wire x_28152;
wire x_28153;
wire x_28154;
wire x_28155;
wire x_28156;
wire x_28157;
wire x_28158;
wire x_28159;
wire x_28160;
wire x_28161;
wire x_28162;
wire x_28163;
wire x_28164;
wire x_28165;
wire x_28166;
wire x_28167;
wire x_28168;
wire x_28169;
wire x_28170;
wire x_28171;
wire x_28172;
wire x_28173;
wire x_28174;
wire x_28175;
wire x_28176;
wire x_28177;
wire x_28178;
wire x_28179;
wire x_28180;
wire x_28181;
wire x_28182;
wire x_28183;
wire x_28184;
wire x_28185;
wire x_28186;
wire x_28187;
wire x_28188;
wire x_28189;
wire x_28190;
wire x_28191;
wire x_28192;
wire x_28193;
wire x_28194;
wire x_28195;
wire x_28196;
wire x_28197;
wire x_28198;
wire x_28199;
wire x_28200;
wire x_28201;
wire x_28202;
wire x_28203;
wire x_28204;
wire x_28205;
wire x_28206;
wire x_28207;
wire x_28208;
wire x_28209;
wire x_28210;
wire x_28211;
wire x_28212;
wire x_28213;
wire x_28214;
wire x_28215;
wire x_28216;
wire x_28217;
wire x_28218;
wire x_28219;
wire x_28220;
wire x_28221;
wire x_28222;
wire x_28223;
wire x_28224;
wire x_28225;
wire x_28226;
wire x_28227;
wire x_28228;
wire x_28229;
wire x_28230;
wire x_28231;
wire x_28232;
wire x_28233;
wire x_28234;
wire x_28235;
wire x_28236;
wire x_28237;
wire x_28238;
wire x_28239;
wire x_28240;
wire x_28241;
wire x_28242;
wire x_28243;
wire x_28244;
wire x_28245;
wire x_28246;
wire x_28247;
wire x_28248;
wire x_28249;
wire x_28250;
wire x_28251;
wire x_28252;
wire x_28253;
wire x_28254;
wire x_28255;
wire x_28256;
wire x_28257;
wire x_28258;
wire x_28259;
wire x_28260;
wire x_28261;
wire x_28262;
wire x_28263;
wire x_28264;
wire x_28265;
wire x_28266;
wire x_28267;
wire x_28268;
wire x_28269;
wire x_28270;
wire x_28271;
wire x_28272;
wire x_28273;
wire x_28274;
wire x_28275;
wire x_28276;
wire x_28277;
wire x_28278;
wire x_28279;
wire x_28280;
wire x_28281;
wire x_28282;
wire x_28283;
wire x_28284;
wire x_28285;
wire x_28286;
wire x_28287;
wire x_28288;
wire x_28289;
wire x_28290;
wire x_28291;
wire x_28292;
wire x_28293;
wire x_28294;
wire x_28295;
wire x_28296;
wire x_28297;
wire x_28298;
wire x_28299;
wire x_28300;
wire x_28301;
wire x_28302;
wire x_28303;
wire x_28304;
wire x_28305;
wire x_28306;
wire x_28307;
wire x_28308;
wire x_28309;
wire x_28310;
wire x_28311;
wire x_28312;
wire x_28313;
wire x_28314;
wire x_28315;
wire x_28316;
wire x_28317;
wire x_28318;
wire x_28319;
wire x_28320;
wire x_28321;
wire x_28322;
wire x_28323;
wire x_28324;
wire x_28325;
wire x_28326;
wire x_28327;
wire x_28328;
wire x_28329;
wire x_28330;
wire x_28331;
wire x_28332;
wire x_28333;
wire x_28334;
wire x_28335;
wire x_28336;
wire x_28337;
wire x_28338;
wire x_28339;
wire x_28340;
wire x_28341;
wire x_28342;
wire x_28343;
wire x_28344;
wire x_28345;
wire x_28346;
wire x_28347;
wire x_28348;
wire x_28349;
wire x_28350;
wire x_28351;
wire x_28352;
wire x_28353;
wire x_28354;
wire x_28355;
wire x_28356;
wire x_28357;
wire x_28358;
wire x_28359;
wire x_28360;
wire x_28361;
wire x_28362;
wire x_28363;
wire x_28364;
wire x_28365;
wire x_28366;
wire x_28367;
wire x_28368;
wire x_28369;
wire x_28370;
wire x_28371;
wire x_28372;
wire x_28373;
wire x_28374;
wire x_28375;
wire x_28376;
wire x_28377;
wire x_28378;
wire x_28379;
wire x_28380;
wire x_28381;
wire x_28382;
wire x_28383;
wire x_28384;
wire x_28385;
wire x_28386;
wire x_28387;
wire x_28388;
wire x_28389;
wire x_28390;
wire x_28391;
wire x_28392;
wire x_28393;
wire x_28394;
wire x_28395;
wire x_28396;
wire x_28397;
wire x_28398;
wire x_28399;
wire x_28400;
wire x_28401;
wire x_28402;
wire x_28403;
wire x_28404;
wire x_28405;
wire x_28406;
wire x_28407;
wire x_28408;
wire x_28409;
wire x_28410;
wire x_28411;
wire x_28412;
wire x_28413;
wire x_28414;
wire x_28415;
wire x_28416;
wire x_28417;
wire x_28418;
wire x_28419;
wire x_28420;
wire x_28421;
wire x_28422;
wire x_28423;
wire x_28424;
wire x_28425;
wire x_28426;
wire x_28427;
wire x_28428;
wire x_28429;
wire x_28430;
wire x_28431;
wire x_28432;
wire x_28433;
wire x_28434;
wire x_28435;
wire x_28436;
wire x_28437;
wire x_28438;
wire x_28439;
wire x_28440;
wire x_28441;
wire x_28442;
wire x_28443;
wire x_28444;
wire x_28445;
wire x_28446;
wire x_28447;
wire x_28448;
wire x_28449;
wire x_28450;
wire x_28451;
wire x_28452;
wire x_28453;
wire x_28454;
wire x_28455;
wire x_28456;
wire x_28457;
wire x_28458;
wire x_28459;
wire x_28460;
wire x_28461;
wire x_28462;
wire x_28463;
wire x_28464;
wire x_28465;
wire x_28466;
wire x_28467;
wire x_28468;
wire x_28469;
wire x_28470;
wire x_28471;
wire x_28472;
wire x_28473;
wire x_28474;
wire x_28475;
wire x_28476;
wire x_28477;
wire x_28478;
wire x_28479;
wire x_28480;
wire x_28481;
wire x_28482;
wire x_28483;
wire x_28484;
wire x_28485;
wire x_28486;
wire x_28487;
wire x_28488;
wire x_28489;
wire x_28490;
wire x_28491;
wire x_28492;
wire x_28493;
wire x_28494;
wire x_28495;
wire x_28496;
wire x_28497;
wire x_28498;
wire x_28499;
wire x_28500;
wire x_28501;
wire x_28502;
wire x_28503;
wire x_28504;
wire x_28505;
wire x_28506;
wire x_28507;
wire x_28508;
wire x_28509;
wire x_28510;
wire x_28511;
wire x_28512;
wire x_28513;
wire x_28514;
wire x_28515;
wire x_28516;
wire x_28517;
wire x_28518;
wire x_28519;
wire x_28520;
wire x_28521;
wire x_28522;
wire x_28523;
wire x_28524;
wire x_28525;
wire x_28526;
wire x_28527;
wire x_28528;
wire x_28529;
wire x_28530;
wire x_28531;
wire x_28532;
wire x_28533;
wire x_28534;
wire x_28535;
wire x_28536;
wire x_28537;
wire x_28538;
wire x_28539;
wire x_28540;
wire x_28541;
wire x_28542;
wire x_28543;
wire x_28544;
wire x_28545;
wire x_28546;
wire x_28547;
wire x_28548;
wire x_28549;
wire x_28550;
wire x_28551;
wire x_28552;
wire x_28553;
wire x_28554;
wire x_28555;
wire x_28556;
wire x_28557;
wire x_28558;
wire x_28559;
wire x_28560;
wire x_28561;
wire x_28562;
wire x_28563;
wire x_28564;
wire x_28565;
wire x_28566;
wire x_28567;
wire x_28568;
wire x_28569;
wire x_28570;
wire x_28571;
wire x_28572;
wire x_28573;
wire x_28574;
wire x_28575;
wire x_28576;
wire x_28577;
wire x_28578;
wire x_28579;
wire x_28580;
wire x_28581;
wire x_28582;
wire x_28583;
wire x_28584;
wire x_28585;
wire x_28586;
wire x_28587;
wire x_28588;
wire x_28589;
wire x_28590;
wire x_28591;
wire x_28592;
wire x_28593;
wire x_28594;
wire x_28595;
wire x_28596;
wire x_28597;
wire x_28598;
wire x_28599;
wire x_28600;
wire x_28601;
wire x_28602;
wire x_28603;
wire x_28604;
wire x_28605;
wire x_28606;
wire x_28607;
wire x_28608;
wire x_28609;
wire x_28610;
wire x_28611;
wire x_28612;
wire x_28613;
wire x_28614;
wire x_28615;
wire x_28616;
wire x_28617;
wire x_28618;
wire x_28619;
wire x_28620;
wire x_28621;
wire x_28622;
wire x_28623;
wire x_28624;
wire x_28625;
wire x_28626;
wire x_28627;
wire x_28628;
wire x_28629;
wire x_28630;
wire x_28631;
wire x_28632;
wire x_28633;
wire x_28634;
wire x_28635;
wire x_28636;
wire x_28637;
wire x_28638;
wire x_28639;
wire x_28640;
wire x_28641;
wire x_28642;
wire x_28643;
wire x_28644;
wire x_28645;
wire x_28646;
wire x_28647;
wire x_28648;
wire x_28649;
wire x_28650;
wire x_28651;
wire x_28652;
wire x_28653;
wire x_28654;
wire x_28655;
wire x_28656;
wire x_28657;
wire x_28658;
wire x_28659;
wire x_28660;
wire x_28661;
wire x_28662;
wire x_28663;
wire x_28664;
wire x_28665;
wire x_28666;
wire x_28667;
wire x_28668;
wire x_28669;
wire x_28670;
wire x_28671;
wire x_28672;
wire x_28673;
wire x_28674;
wire x_28675;
wire x_28676;
wire x_28677;
wire x_28678;
wire x_28679;
wire x_28680;
wire x_28681;
wire x_28682;
wire x_28683;
wire x_28684;
wire x_28685;
wire x_28686;
wire x_28687;
wire x_28688;
wire x_28689;
wire x_28690;
wire x_28691;
wire x_28692;
wire x_28693;
wire x_28694;
wire x_28695;
wire x_28696;
wire x_28697;
wire x_28698;
wire x_28699;
wire x_28700;
wire x_28701;
wire x_28702;
wire x_28703;
wire x_28704;
wire x_28705;
wire x_28706;
wire x_28707;
wire x_28708;
wire x_28709;
wire x_28710;
wire x_28711;
wire x_28712;
wire x_28713;
wire x_28714;
wire x_28715;
wire x_28716;
wire x_28717;
wire x_28718;
wire x_28719;
wire x_28720;
wire x_28721;
wire x_28722;
wire x_28723;
wire x_28724;
wire x_28725;
wire x_28726;
wire x_28727;
wire x_28728;
wire x_28729;
wire x_28730;
wire x_28731;
wire x_28732;
wire x_28733;
wire x_28734;
wire x_28735;
wire x_28736;
wire x_28737;
wire x_28738;
wire x_28739;
wire x_28740;
wire x_28741;
wire x_28742;
wire x_28743;
wire x_28744;
wire x_28745;
wire x_28746;
wire x_28747;
wire x_28748;
wire x_28749;
wire x_28750;
wire x_28751;
wire x_28752;
wire x_28753;
wire x_28754;
wire x_28755;
wire x_28756;
wire x_28757;
wire x_28758;
wire x_28759;
wire x_28760;
wire x_28761;
wire x_28762;
wire x_28763;
wire x_28764;
wire x_28765;
wire x_28766;
wire x_28767;
wire x_28768;
wire x_28769;
wire x_28770;
wire x_28771;
wire x_28772;
wire x_28773;
wire x_28774;
wire x_28775;
wire x_28776;
wire x_28777;
wire x_28778;
wire x_28779;
wire x_28780;
wire x_28781;
wire x_28782;
wire x_28783;
wire x_28784;
wire x_28785;
wire x_28786;
wire x_28787;
wire x_28788;
wire x_28789;
wire x_28790;
wire x_28791;
wire x_28792;
wire x_28793;
wire x_28794;
wire x_28795;
wire x_28796;
wire x_28797;
wire x_28798;
wire x_28799;
wire x_28800;
wire x_28801;
wire x_28802;
wire x_28803;
wire x_28804;
wire x_28805;
wire x_28806;
wire x_28807;
wire x_28808;
wire x_28809;
wire x_28810;
wire x_28811;
wire x_28812;
wire x_28813;
wire x_28814;
wire x_28815;
wire x_28816;
wire x_28817;
wire x_28818;
wire x_28819;
wire x_28820;
wire x_28821;
wire x_28822;
wire x_28823;
wire x_28824;
wire x_28825;
wire x_28826;
wire x_28827;
wire x_28828;
wire x_28829;
wire x_28830;
wire x_28831;
wire x_28832;
wire x_28833;
wire x_28834;
wire x_28835;
wire x_28836;
wire x_28837;
wire x_28838;
wire x_28839;
wire x_28840;
wire x_28841;
wire x_28842;
wire x_28843;
wire x_28844;
wire x_28845;
wire x_28846;
wire x_28847;
wire x_28848;
wire x_28849;
wire x_28850;
wire x_28851;
wire x_28852;
wire x_28853;
wire x_28854;
wire x_28855;
wire x_28856;
wire x_28857;
wire x_28858;
wire x_28859;
wire x_28860;
wire x_28861;
wire x_28862;
wire x_28863;
wire x_28864;
wire x_28865;
wire x_28866;
wire x_28867;
wire x_28868;
wire x_28869;
wire x_28870;
wire x_28871;
wire x_28872;
wire x_28873;
wire x_28874;
wire x_28875;
wire x_28876;
wire x_28877;
wire x_28878;
wire x_28879;
wire x_28880;
wire x_28881;
wire x_28882;
wire x_28883;
wire x_28884;
wire x_28885;
wire x_28886;
wire x_28887;
wire x_28888;
wire x_28889;
wire x_28890;
wire x_28891;
wire x_28892;
wire x_28893;
wire x_28894;
wire x_28895;
wire x_28896;
wire x_28897;
wire x_28898;
wire x_28899;
wire x_28900;
wire x_28901;
wire x_28902;
wire x_28903;
wire x_28904;
wire x_28905;
wire x_28906;
wire x_28907;
wire x_28908;
wire x_28909;
wire x_28910;
wire x_28911;
wire x_28912;
wire x_28913;
wire x_28914;
wire x_28915;
wire x_28916;
wire x_28917;
wire x_28918;
wire x_28919;
wire x_28920;
wire x_28921;
wire x_28922;
wire x_28923;
wire x_28924;
wire x_28925;
wire x_28926;
wire x_28927;
wire x_28928;
wire x_28929;
wire x_28930;
wire x_28931;
wire x_28932;
wire x_28933;
wire x_28934;
wire x_28935;
wire x_28936;
wire x_28937;
wire x_28938;
wire x_28939;
wire x_28940;
wire x_28941;
wire x_28942;
wire x_28943;
wire x_28944;
wire x_28945;
wire x_28946;
wire x_28947;
wire x_28948;
wire x_28949;
wire x_28950;
wire x_28951;
wire x_28952;
wire x_28953;
wire x_28954;
wire x_28955;
wire x_28956;
wire x_28957;
wire x_28958;
wire x_28959;
wire x_28960;
wire x_28961;
wire x_28962;
wire x_28963;
wire x_28964;
wire x_28965;
wire x_28966;
wire x_28967;
wire x_28968;
wire x_28969;
wire x_28970;
wire x_28971;
wire x_28972;
wire x_28973;
wire x_28974;
wire x_28975;
wire x_28976;
wire x_28977;
wire x_28978;
wire x_28979;
wire x_28980;
wire x_28981;
wire x_28982;
wire x_28983;
wire x_28984;
wire x_28985;
wire x_28986;
wire x_28987;
wire x_28988;
wire x_28989;
wire x_28990;
wire x_28991;
wire x_28992;
wire x_28993;
wire x_28994;
wire x_28995;
wire x_28996;
wire x_28997;
wire x_28998;
wire x_28999;
wire x_29000;
wire x_29001;
wire x_29002;
wire x_29003;
wire x_29004;
wire x_29005;
wire x_29006;
wire x_29007;
wire x_29008;
wire x_29009;
wire x_29010;
wire x_29011;
wire x_29012;
wire x_29013;
wire x_29014;
wire x_29015;
wire x_29016;
wire x_29017;
wire x_29018;
wire x_29019;
wire x_29020;
wire x_29021;
wire x_29022;
wire x_29023;
wire x_29024;
wire x_29025;
wire x_29026;
wire x_29027;
wire x_29028;
wire x_29029;
wire x_29030;
wire x_29031;
wire x_29032;
wire x_29033;
wire x_29034;
wire x_29035;
wire x_29036;
wire x_29037;
wire x_29038;
wire x_29039;
wire x_29040;
wire x_29041;
wire x_29042;
wire x_29043;
wire x_29044;
wire x_29045;
wire x_29046;
wire x_29047;
wire x_29048;
wire x_29049;
wire x_29050;
wire x_29051;
wire x_29052;
wire x_29053;
wire x_29054;
wire x_29055;
wire x_29056;
wire x_29057;
wire x_29058;
wire x_29059;
wire x_29060;
wire x_29061;
wire x_29062;
wire x_29063;
wire x_29064;
wire x_29065;
wire x_29066;
wire x_29067;
wire x_29068;
wire x_29069;
wire x_29070;
wire x_29071;
wire x_29072;
wire x_29073;
wire x_29074;
wire x_29075;
wire x_29076;
wire x_29077;
wire x_29078;
wire x_29079;
wire x_29080;
wire x_29081;
wire x_29082;
wire x_29083;
wire x_29084;
wire x_29085;
wire x_29086;
wire x_29087;
wire x_29088;
wire x_29089;
wire x_29090;
wire x_29091;
wire x_29092;
wire x_29093;
wire x_29094;
wire x_29095;
wire x_29096;
wire x_29097;
wire x_29098;
wire x_29099;
wire x_29100;
wire x_29101;
wire x_29102;
wire x_29103;
wire x_29104;
wire x_29105;
wire x_29106;
wire x_29107;
wire x_29108;
wire x_29109;
wire x_29110;
wire x_29111;
wire x_29112;
wire x_29113;
wire x_29114;
wire x_29115;
wire x_29116;
wire x_29117;
wire x_29118;
wire x_29119;
wire x_29120;
wire x_29121;
wire x_29122;
wire x_29123;
wire x_29124;
wire x_29125;
wire x_29126;
wire x_29127;
wire x_29128;
wire x_29129;
wire x_29130;
wire x_29131;
wire x_29132;
wire x_29133;
wire x_29134;
wire x_29135;
wire x_29136;
wire x_29137;
wire x_29138;
wire x_29139;
wire x_29140;
wire x_29141;
wire x_29142;
wire x_29143;
wire x_29144;
wire x_29145;
wire x_29146;
wire x_29147;
wire x_29148;
wire x_29149;
wire x_29150;
wire x_29151;
wire x_29152;
wire x_29153;
wire x_29154;
wire x_29155;
wire x_29156;
wire x_29157;
wire x_29158;
wire x_29159;
wire x_29160;
wire x_29161;
wire x_29162;
wire x_29163;
wire x_29164;
wire x_29165;
wire x_29166;
wire x_29167;
wire x_29168;
wire x_29169;
wire x_29170;
wire x_29171;
wire x_29172;
wire x_29173;
wire x_29174;
wire x_29175;
wire x_29176;
wire x_29177;
wire x_29178;
wire x_29179;
wire x_29180;
wire x_29181;
wire x_29182;
wire x_29183;
wire x_29184;
wire x_29185;
wire x_29186;
wire x_29187;
wire x_29188;
wire x_29189;
wire x_29190;
wire x_29191;
wire x_29192;
wire x_29193;
wire x_29194;
wire x_29195;
wire x_29196;
wire x_29197;
wire x_29198;
wire x_29199;
wire x_29200;
wire x_29201;
wire x_29202;
wire x_29203;
wire x_29204;
wire x_29205;
wire x_29206;
wire x_29207;
wire x_29208;
wire x_29209;
wire x_29210;
wire x_29211;
wire x_29212;
wire x_29213;
wire x_29214;
wire x_29215;
wire x_29216;
wire x_29217;
wire x_29218;
wire x_29219;
wire x_29220;
wire x_29221;
wire x_29222;
wire x_29223;
wire x_29224;
wire x_29225;
wire x_29226;
wire x_29227;
wire x_29228;
wire x_29229;
wire x_29230;
wire x_29231;
wire x_29232;
wire x_29233;
wire x_29234;
wire x_29235;
wire x_29236;
wire x_29237;
wire x_29238;
wire x_29239;
wire x_29240;
wire x_29241;
wire x_29242;
wire x_29243;
wire x_29244;
wire x_29245;
wire x_29246;
wire x_29247;
wire x_29248;
wire x_29249;
wire x_29250;
wire x_29251;
wire x_29252;
wire x_29253;
wire x_29254;
wire x_29255;
wire x_29256;
wire x_29257;
wire x_29258;
wire x_29259;
wire x_29260;
wire x_29261;
wire x_29262;
wire x_29263;
wire x_29264;
wire x_29265;
wire x_29266;
wire x_29267;
wire x_29268;
wire x_29269;
wire x_29270;
wire x_29271;
wire x_29272;
wire x_29273;
wire x_29274;
wire x_29275;
wire x_29276;
wire x_29277;
wire x_29278;
wire x_29279;
wire x_29280;
wire x_29281;
wire x_29282;
wire x_29283;
wire x_29284;
wire x_29285;
wire x_29286;
wire x_29287;
wire x_29288;
wire x_29289;
wire x_29290;
wire x_29291;
wire x_29292;
wire x_29293;
wire x_29294;
wire x_29295;
wire x_29296;
wire x_29297;
wire x_29298;
wire x_29299;
wire x_29300;
wire x_29301;
wire x_29302;
wire x_29303;
wire x_29304;
wire x_29305;
wire x_29306;
wire x_29307;
wire x_29308;
wire x_29309;
wire x_29310;
wire x_29311;
wire x_29312;
wire x_29313;
wire x_29314;
wire x_29315;
wire x_29316;
wire x_29317;
wire x_29318;
wire x_29319;
wire x_29320;
wire x_29321;
wire x_29322;
wire x_29323;
wire x_29324;
wire x_29325;
wire x_29326;
wire x_29327;
wire x_29328;
wire x_29329;
wire x_29330;
wire x_29331;
wire x_29332;
wire x_29333;
wire x_29334;
wire x_29335;
wire x_29336;
wire x_29337;
wire x_29338;
wire x_29339;
wire x_29340;
wire x_29341;
wire x_29342;
wire x_29343;
wire x_29344;
wire x_29345;
wire x_29346;
wire x_29347;
wire x_29348;
wire x_29349;
wire x_29350;
wire x_29351;
wire x_29352;
wire x_29353;
wire x_29354;
wire x_29355;
wire x_29356;
wire x_29357;
wire x_29358;
wire x_29359;
wire x_29360;
wire x_29361;
wire x_29362;
wire x_29363;
wire x_29364;
wire x_29365;
wire x_29366;
wire x_29367;
wire x_29368;
wire x_29369;
wire x_29370;
wire x_29371;
wire x_29372;
wire x_29373;
wire x_29374;
wire x_29375;
wire x_29376;
wire x_29377;
wire x_29378;
wire x_29379;
wire x_29380;
wire x_29381;
wire x_29382;
wire x_29383;
wire x_29384;
wire x_29385;
wire x_29386;
wire x_29387;
wire x_29388;
wire x_29389;
wire x_29390;
wire x_29391;
wire x_29392;
wire x_29393;
wire x_29394;
wire x_29395;
wire x_29396;
wire x_29397;
wire x_29398;
wire x_29399;
wire x_29400;
wire x_29401;
wire x_29402;
wire x_29403;
wire x_29404;
wire x_29405;
wire x_29406;
wire x_29407;
wire x_29408;
wire x_29409;
wire x_29410;
wire x_29411;
wire x_29412;
wire x_29413;
wire x_29414;
wire x_29415;
wire x_29416;
wire x_29417;
wire x_29418;
wire x_29419;
wire x_29420;
wire x_29421;
wire x_29422;
wire x_29423;
wire x_29424;
wire x_29425;
wire x_29426;
wire x_29427;
wire x_29428;
wire x_29429;
wire x_29430;
wire x_29431;
wire x_29432;
wire x_29433;
wire x_29434;
wire x_29435;
wire x_29436;
wire x_29437;
wire x_29438;
wire x_29439;
wire x_29440;
wire x_29441;
wire x_29442;
wire x_29443;
wire x_29444;
wire x_29445;
wire x_29446;
wire x_29447;
wire x_29448;
wire x_29449;
wire x_29450;
wire x_29451;
wire x_29452;
wire x_29453;
wire x_29454;
wire x_29455;
wire x_29456;
wire x_29457;
wire x_29458;
wire x_29459;
wire x_29460;
wire x_29461;
wire x_29462;
wire x_29463;
wire x_29464;
wire x_29465;
wire x_29466;
wire x_29467;
wire x_29468;
wire x_29469;
wire x_29470;
wire x_29471;
wire x_29472;
wire x_29473;
wire x_29474;
wire x_29475;
wire x_29476;
wire x_29477;
wire x_29478;
wire x_29479;
wire x_29480;
wire x_29481;
wire x_29482;
wire x_29483;
wire x_29484;
wire x_29485;
wire x_29486;
wire x_29487;
wire x_29488;
wire x_29489;
wire x_29490;
wire x_29491;
wire x_29492;
wire x_29493;
wire x_29494;
wire x_29495;
wire x_29496;
wire x_29497;
wire x_29498;
wire x_29499;
wire x_29500;
wire x_29501;
wire x_29502;
wire x_29503;
wire x_29504;
wire x_29505;
wire x_29506;
wire x_29507;
wire x_29508;
wire x_29509;
wire x_29510;
wire x_29511;
wire x_29512;
wire x_29513;
wire x_29514;
wire x_29515;
wire x_29516;
wire x_29517;
wire x_29518;
wire x_29519;
wire x_29520;
wire x_29521;
wire x_29522;
wire x_29523;
wire x_29524;
wire x_29525;
wire x_29526;
wire x_29527;
wire x_29528;
wire x_29529;
wire x_29530;
wire x_29531;
wire x_29532;
wire x_29533;
wire x_29534;
wire x_29535;
wire x_29536;
wire x_29537;
wire x_29538;
wire x_29539;
wire x_29540;
wire x_29541;
wire x_29542;
wire x_29543;
wire x_29544;
wire x_29545;
wire x_29546;
wire x_29547;
wire x_29548;
wire x_29549;
wire x_29550;
wire x_29551;
wire x_29552;
wire x_29553;
wire x_29554;
wire x_29555;
wire x_29556;
wire x_29557;
wire x_29558;
wire x_29559;
wire x_29560;
wire x_29561;
wire x_29562;
wire x_29563;
wire x_29564;
wire x_29565;
wire x_29566;
wire x_29567;
wire x_29568;
wire x_29569;
wire x_29570;
wire x_29571;
wire x_29572;
wire x_29573;
wire x_29574;
wire x_29575;
wire x_29576;
wire x_29577;
wire x_29578;
wire x_29579;
wire x_29580;
wire x_29581;
wire x_29582;
wire x_29583;
wire x_29584;
wire x_29585;
wire x_29586;
wire x_29587;
wire x_29588;
wire x_29589;
wire x_29590;
wire x_29591;
wire x_29592;
wire x_29593;
wire x_29594;
wire x_29595;
wire x_29596;
wire x_29597;
wire x_29598;
wire x_29599;
wire x_29600;
wire x_29601;
wire x_29602;
wire x_29603;
wire x_29604;
wire x_29605;
wire x_29606;
wire x_29607;
wire x_29608;
wire x_29609;
wire x_29610;
wire x_29611;
wire x_29612;
wire x_29613;
wire x_29614;
wire x_29615;
wire x_29616;
wire x_29617;
wire x_29618;
wire x_29619;
wire x_29620;
wire x_29621;
wire x_29622;
wire x_29623;
wire x_29624;
wire x_29625;
wire x_29626;
wire x_29627;
wire x_29628;
wire x_29629;
wire x_29630;
wire x_29631;
wire x_29632;
wire x_29633;
wire x_29634;
wire x_29635;
wire x_29636;
wire x_29637;
wire x_29638;
wire x_29639;
wire x_29640;
wire x_29641;
wire x_29642;
wire x_29643;
wire x_29644;
wire x_29645;
wire x_29646;
wire x_29647;
wire x_29648;
wire x_29649;
wire x_29650;
wire x_29651;
wire x_29652;
wire x_29653;
wire x_29654;
wire x_29655;
wire x_29656;
wire x_29657;
wire x_29658;
wire x_29659;
wire x_29660;
wire x_29661;
wire x_29662;
wire x_29663;
wire x_29664;
wire x_29665;
wire x_29666;
wire x_29667;
wire x_29668;
wire x_29669;
wire x_29670;
wire x_29671;
wire x_29672;
wire x_29673;
wire x_29674;
wire x_29675;
wire x_29676;
wire x_29677;
wire x_29678;
wire x_29679;
wire x_29680;
wire x_29681;
wire x_29682;
wire x_29683;
wire x_29684;
wire x_29685;
wire x_29686;
wire x_29687;
wire x_29688;
wire x_29689;
wire x_29690;
wire x_29691;
wire x_29692;
wire x_29693;
wire x_29694;
wire x_29695;
wire x_29696;
wire x_29697;
wire x_29698;
wire x_29699;
wire x_29700;
wire x_29701;
wire x_29702;
wire x_29703;
wire x_29704;
wire x_29705;
wire x_29706;
wire x_29707;
wire x_29708;
wire x_29709;
wire x_29710;
wire x_29711;
wire x_29712;
wire x_29713;
wire x_29714;
wire x_29715;
wire x_29716;
wire x_29717;
wire x_29718;
wire x_29719;
wire x_29720;
wire x_29721;
wire x_29722;
wire x_29723;
wire x_29724;
wire x_29725;
wire x_29726;
wire x_29727;
wire x_29728;
wire x_29729;
wire x_29730;
wire x_29731;
wire x_29732;
wire x_29733;
wire x_29734;
wire x_29735;
wire x_29736;
wire x_29737;
wire x_29738;
wire x_29739;
wire x_29740;
wire x_29741;
wire x_29742;
wire x_29743;
wire x_29744;
wire x_29745;
wire x_29746;
wire x_29747;
wire x_29748;
wire x_29749;
wire x_29750;
wire x_29751;
wire x_29752;
wire x_29753;
wire x_29754;
wire x_29755;
wire x_29756;
wire x_29757;
wire x_29758;
wire x_29759;
wire x_29760;
wire x_29761;
wire x_29762;
wire x_29763;
wire x_29764;
wire x_29765;
wire x_29766;
wire x_29767;
wire x_29768;
wire x_29769;
wire x_29770;
wire x_29771;
wire x_29772;
wire x_29773;
wire x_29774;
wire x_29775;
wire x_29776;
wire x_29777;
wire x_29778;
wire x_29779;
wire x_29780;
wire x_29781;
wire x_29782;
wire x_29783;
wire x_29784;
wire x_29785;
wire x_29786;
wire x_29787;
wire x_29788;
wire x_29789;
wire x_29790;
wire x_29791;
wire x_29792;
wire x_29793;
wire x_29794;
wire x_29795;
wire x_29796;
wire x_29797;
wire x_29798;
wire x_29799;
wire x_29800;
wire x_29801;
wire x_29802;
wire x_29803;
wire x_29804;
wire x_29805;
wire x_29806;
wire x_29807;
wire x_29808;
wire x_29809;
wire x_29810;
wire x_29811;
wire x_29812;
wire x_29813;
wire x_29814;
wire x_29815;
wire x_29816;
wire x_29817;
wire x_29818;
wire x_29819;
wire x_29820;
wire x_29821;
wire x_29822;
wire x_29823;
wire x_29824;
wire x_29825;
wire x_29826;
wire x_29827;
wire x_29828;
wire x_29829;
wire x_29830;
wire x_29831;
wire x_29832;
wire x_29833;
wire x_29834;
wire x_29835;
wire x_29836;
wire x_29837;
wire x_29838;
wire x_29839;
wire x_29840;
wire x_29841;
wire x_29842;
wire x_29843;
wire x_29844;
wire x_29845;
wire x_29846;
wire x_29847;
wire x_29848;
wire x_29849;
wire x_29850;
wire x_29851;
wire x_29852;
wire x_29853;
wire x_29854;
wire x_29855;
wire x_29856;
wire x_29857;
wire x_29858;
wire x_29859;
wire x_29860;
wire x_29861;
wire x_29862;
wire x_29863;
wire x_29864;
wire x_29865;
wire x_29866;
wire x_29867;
wire x_29868;
wire x_29869;
wire x_29870;
wire x_29871;
wire x_29872;
wire x_29873;
wire x_29874;
wire x_29875;
wire x_29876;
wire x_29877;
wire x_29878;
wire x_29879;
wire x_29880;
wire x_29881;
wire x_29882;
wire x_29883;
wire x_29884;
wire x_29885;
wire x_29886;
wire x_29887;
wire x_29888;
wire x_29889;
wire x_29890;
wire x_29891;
wire x_29892;
wire x_29893;
wire x_29894;
wire x_29895;
wire x_29896;
wire x_29897;
wire x_29898;
wire x_29899;
wire x_29900;
wire x_29901;
wire x_29902;
wire x_29903;
wire x_29904;
wire x_29905;
wire x_29906;
wire x_29907;
wire x_29908;
wire x_29909;
wire x_29910;
wire x_29911;
wire x_29912;
wire x_29913;
wire x_29914;
wire x_29915;
wire x_29916;
wire x_29917;
wire x_29918;
wire x_29919;
wire x_29920;
wire x_29921;
wire x_29922;
wire x_29923;
wire x_29924;
wire x_29925;
wire x_29926;
wire x_29927;
wire x_29928;
wire x_29929;
wire x_29930;
wire x_29931;
wire x_29932;
wire x_29933;
wire x_29934;
wire x_29935;
wire x_29936;
wire x_29937;
wire x_29938;
wire x_29939;
wire x_29940;
wire x_29941;
wire x_29942;
wire x_29943;
wire x_29944;
wire x_29945;
wire x_29946;
wire x_29947;
wire x_29948;
wire x_29949;
wire x_29950;
wire x_29951;
wire x_29952;
wire x_29953;
wire x_29954;
wire x_29955;
wire x_29956;
wire x_29957;
wire x_29958;
wire x_29959;
wire x_29960;
wire x_29961;
wire x_29962;
wire x_29963;
wire x_29964;
wire x_29965;
wire x_29966;
wire x_29967;
wire x_29968;
wire x_29969;
wire x_29970;
wire x_29971;
wire x_29972;
wire x_29973;
wire x_29974;
wire x_29975;
wire x_29976;
wire x_29977;
wire x_29978;
wire x_29979;
wire x_29980;
wire x_29981;
wire x_29982;
wire x_29983;
wire x_29984;
wire x_29985;
wire x_29986;
wire x_29987;
wire x_29988;
wire x_29989;
wire x_29990;
wire x_29991;
wire x_29992;
wire x_29993;
wire x_29994;
wire x_29995;
wire x_29996;
wire x_29997;
wire x_29998;
wire x_29999;
wire x_30000;
wire x_30001;
wire x_30002;
wire x_30003;
wire x_30004;
wire x_30005;
wire x_30006;
wire x_30007;
wire x_30008;
wire x_30009;
wire x_30010;
wire x_30011;
wire x_30012;
wire x_30013;
wire x_30014;
wire x_30015;
wire x_30016;
wire x_30017;
wire x_30018;
wire x_30019;
wire x_30020;
wire x_30021;
wire x_30022;
wire x_30023;
wire x_30024;
wire x_30025;
wire x_30026;
wire x_30027;
wire x_30028;
wire x_30029;
wire x_30030;
wire x_30031;
wire x_30032;
wire x_30033;
wire x_30034;
wire x_30035;
wire x_30036;
wire x_30037;
wire x_30038;
wire x_30039;
wire x_30040;
wire x_30041;
wire x_30042;
wire x_30043;
wire x_30044;
wire x_30045;
wire x_30046;
wire x_30047;
wire x_30048;
wire x_30049;
wire x_30050;
wire x_30051;
wire x_30052;
wire x_30053;
wire x_30054;
wire x_30055;
wire x_30056;
wire x_30057;
wire x_30058;
wire x_30059;
wire x_30060;
wire x_30061;
wire x_30062;
wire x_30063;
wire x_30064;
wire x_30065;
wire x_30066;
wire x_30067;
wire x_30068;
wire x_30069;
wire x_30070;
wire x_30071;
wire x_30072;
wire x_30073;
wire x_30074;
wire x_30075;
wire x_30076;
wire x_30077;
wire x_30078;
wire x_30079;
wire x_30080;
wire x_30081;
wire x_30082;
wire x_30083;
wire x_30084;
wire x_30085;
wire x_30086;
wire x_30087;
wire x_30088;
wire x_30089;
wire x_30090;
wire x_30091;
wire x_30092;
wire x_30093;
wire x_30094;
wire x_30095;
wire x_30096;
wire x_30097;
wire x_30098;
wire x_30099;
wire x_30100;
wire x_30101;
wire x_30102;
wire x_30103;
wire x_30104;
wire x_30105;
wire x_30106;
wire x_30107;
wire x_30108;
wire x_30109;
wire x_30110;
wire x_30111;
wire x_30112;
wire x_30113;
wire x_30114;
wire x_30115;
wire x_30116;
wire x_30117;
wire x_30118;
wire x_30119;
wire x_30120;
wire x_30121;
wire x_30122;
wire x_30123;
wire x_30124;
wire x_30125;
wire x_30126;
wire x_30127;
wire x_30128;
wire x_30129;
wire x_30130;
wire x_30131;
wire x_30132;
wire x_30133;
wire x_30134;
wire x_30135;
wire x_30136;
wire x_30137;
wire x_30138;
wire x_30139;
wire x_30140;
wire x_30141;
wire x_30142;
wire x_30143;
wire x_30144;
wire x_30145;
wire x_30146;
wire x_30147;
wire x_30148;
wire x_30149;
wire x_30150;
wire x_30151;
wire x_30152;
wire x_30153;
wire x_30154;
wire x_30155;
wire x_30156;
wire x_30157;
wire x_30158;
wire x_30159;
wire x_30160;
wire x_30161;
wire x_30162;
wire x_30163;
wire x_30164;
wire x_30165;
wire x_30166;
wire x_30167;
wire x_30168;
wire x_30169;
wire x_30170;
wire x_30171;
wire x_30172;
wire x_30173;
wire x_30174;
wire x_30175;
wire x_30176;
wire x_30177;
wire x_30178;
wire x_30179;
wire x_30180;
wire x_30181;
wire x_30182;
wire x_30183;
wire x_30184;
wire x_30185;
wire x_30186;
wire x_30187;
wire x_30188;
wire x_30189;
wire x_30190;
wire x_30191;
wire x_30192;
wire x_30193;
wire x_30194;
wire x_30195;
wire x_30196;
wire x_30197;
wire x_30198;
wire x_30199;
wire x_30200;
wire x_30201;
wire x_30202;
wire x_30203;
wire x_30204;
wire x_30205;
wire x_30206;
wire x_30207;
wire x_30208;
wire x_30209;
wire x_30210;
wire x_30211;
wire x_30212;
wire x_30213;
wire x_30214;
wire x_30215;
wire x_30216;
wire x_30217;
wire x_30218;
wire x_30219;
wire x_30220;
wire x_30221;
wire x_30222;
wire x_30223;
wire x_30224;
wire x_30225;
wire x_30226;
wire x_30227;
wire x_30228;
wire x_30229;
wire x_30230;
wire x_30231;
wire x_30232;
wire x_30233;
wire x_30234;
wire x_30235;
wire x_30236;
wire x_30237;
wire x_30238;
wire x_30239;
wire x_30240;
wire x_30241;
wire x_30242;
wire x_30243;
wire x_30244;
wire x_30245;
wire x_30246;
wire x_30247;
wire x_30248;
wire x_30249;
wire x_30250;
wire x_30251;
wire x_30252;
wire x_30253;
wire x_30254;
wire x_30255;
wire x_30256;
wire x_30257;
wire x_30258;
wire x_30259;
wire x_30260;
wire x_30261;
wire x_30262;
wire x_30263;
wire x_30264;
wire x_30265;
wire x_30266;
wire x_30267;
wire x_30268;
wire x_30269;
wire x_30270;
wire x_30271;
wire x_30272;
wire x_30273;
wire x_30274;
wire x_30275;
wire x_30276;
wire x_30277;
wire x_30278;
wire x_30279;
wire x_30280;
wire x_30281;
wire x_30282;
wire x_30283;
wire x_30284;
wire x_30285;
wire x_30286;
wire x_30287;
wire x_30288;
wire x_30289;
wire x_30290;
wire x_30291;
wire x_30292;
wire x_30293;
wire x_30294;
wire x_30295;
wire x_30296;
wire x_30297;
wire x_30298;
wire x_30299;
wire x_30300;
wire x_30301;
wire x_30302;
wire x_30303;
wire x_30304;
wire x_30305;
wire x_30306;
wire x_30307;
wire x_30308;
wire x_30309;
wire x_30310;
wire x_30311;
wire x_30312;
wire x_30313;
wire x_30314;
wire x_30315;
wire x_30316;
wire x_30317;
wire x_30318;
wire x_30319;
wire x_30320;
wire x_30321;
wire x_30322;
wire x_30323;
wire x_30324;
wire x_30325;
wire x_30326;
wire x_30327;
wire x_30328;
wire x_30329;
wire x_30330;
wire x_30331;
wire x_30332;
wire x_30333;
wire x_30334;
wire x_30335;
wire x_30336;
wire x_30337;
wire x_30338;
wire x_30339;
wire x_30340;
wire x_30341;
wire x_30342;
wire x_30343;
wire x_30344;
wire x_30345;
wire x_30346;
wire x_30347;
wire x_30348;
wire x_30349;
wire x_30350;
wire x_30351;
wire x_30352;
wire x_30353;
wire x_30354;
wire x_30355;
wire x_30356;
wire x_30357;
wire x_30358;
wire x_30359;
wire x_30360;
wire x_30361;
wire x_30362;
wire x_30363;
wire x_30364;
wire x_30365;
wire x_30366;
wire x_30367;
wire x_30368;
wire x_30369;
wire x_30370;
wire x_30371;
wire x_30372;
wire x_30373;
wire x_30374;
wire x_30375;
wire x_30376;
wire x_30377;
wire x_30378;
wire x_30379;
wire x_30380;
wire x_30381;
wire x_30382;
wire x_30383;
wire x_30384;
wire x_30385;
wire x_30386;
wire x_30387;
wire x_30388;
wire x_30389;
wire x_30390;
wire x_30391;
wire x_30392;
wire x_30393;
wire x_30394;
wire x_30395;
wire x_30396;
wire x_30397;
wire x_30398;
wire x_30399;
wire x_30400;
wire x_30401;
wire x_30402;
wire x_30403;
wire x_30404;
wire x_30405;
wire x_30406;
wire x_30407;
wire x_30408;
wire x_30409;
wire x_30410;
wire x_30411;
wire x_30412;
wire x_30413;
wire x_30414;
wire x_30415;
wire x_30416;
wire x_30417;
wire x_30418;
wire x_30419;
wire x_30420;
wire x_30421;
wire x_30422;
wire x_30423;
wire x_30424;
wire x_30425;
wire x_30426;
wire x_30427;
wire x_30428;
wire x_30429;
wire x_30430;
wire x_30431;
wire x_30432;
wire x_30433;
wire x_30434;
wire x_30435;
wire x_30436;
wire x_30437;
wire x_30438;
wire x_30439;
wire x_30440;
wire x_30441;
wire x_30442;
wire x_30443;
wire x_30444;
wire x_30445;
wire x_30446;
wire x_30447;
wire x_30448;
wire x_30449;
wire x_30450;
wire x_30451;
wire x_30452;
wire x_30453;
wire x_30454;
wire x_30455;
wire x_30456;
wire x_30457;
wire x_30458;
wire x_30459;
wire x_30460;
wire x_30461;
wire x_30462;
wire x_30463;
wire x_30464;
wire x_30465;
wire x_30466;
wire x_30467;
wire x_30468;
wire x_30469;
wire x_30470;
wire x_30471;
wire x_30472;
wire x_30473;
wire x_30474;
wire x_30475;
wire x_30476;
wire x_30477;
wire x_30478;
wire x_30479;
wire x_30480;
wire x_30481;
wire x_30482;
wire x_30483;
wire x_30484;
wire x_30485;
wire x_30486;
wire x_30487;
wire x_30488;
wire x_30489;
wire x_30490;
wire x_30491;
wire x_30492;
wire x_30493;
wire x_30494;
wire x_30495;
wire x_30496;
wire x_30497;
wire x_30498;
wire x_30499;
wire x_30500;
wire x_30501;
wire x_30502;
wire x_30503;
wire x_30504;
wire x_30505;
wire x_30506;
wire x_30507;
wire x_30508;
wire x_30509;
wire x_30510;
wire x_30511;
wire x_30512;
wire x_30513;
wire x_30514;
wire x_30515;
wire x_30516;
wire x_30517;
wire x_30518;
wire x_30519;
wire x_30520;
wire x_30521;
wire x_30522;
wire x_30523;
wire x_30524;
wire x_30525;
wire x_30526;
wire x_30527;
wire x_30528;
wire x_30529;
wire x_30530;
wire x_30531;
wire x_30532;
wire x_30533;
wire x_30534;
wire x_30535;
wire x_30536;
wire x_30537;
wire x_30538;
wire x_30539;
wire x_30540;
wire x_30541;
wire x_30542;
wire x_30543;
wire x_30544;
wire x_30545;
wire x_30546;
wire x_30547;
wire x_30548;
wire x_30549;
wire x_30550;
wire x_30551;
wire x_30552;
wire x_30553;
wire x_30554;
wire x_30555;
wire x_30556;
wire x_30557;
wire x_30558;
wire x_30559;
wire x_30560;
wire x_30561;
wire x_30562;
wire x_30563;
wire x_30564;
wire x_30565;
wire x_30566;
wire x_30567;
wire x_30568;
wire x_30569;
wire x_30570;
wire x_30571;
wire x_30572;
wire x_30573;
wire x_30574;
wire x_30575;
wire x_30576;
wire x_30577;
wire x_30578;
wire x_30579;
wire x_30580;
wire x_30581;
wire x_30582;
wire x_30583;
wire x_30584;
wire x_30585;
wire x_30586;
wire x_30587;
wire x_30588;
wire x_30589;
wire x_30590;
wire x_30591;
wire x_30592;
wire x_30593;
wire x_30594;
wire x_30595;
wire x_30596;
wire x_30597;
wire x_30598;
wire x_30599;
wire x_30600;
wire x_30601;
wire x_30602;
wire x_30603;
wire x_30604;
wire x_30605;
wire x_30606;
wire x_30607;
wire x_30608;
wire x_30609;
wire x_30610;
wire x_30611;
wire x_30612;
wire x_30613;
wire x_30614;
wire x_30615;
wire x_30616;
wire x_30617;
wire x_30618;
wire x_30619;
wire x_30620;
wire x_30621;
wire x_30622;
wire x_30623;
wire x_30624;
wire x_30625;
wire x_30626;
wire x_30627;
wire x_30628;
wire x_30629;
wire x_30630;
wire x_30631;
wire x_30632;
wire x_30633;
wire x_30634;
wire x_30635;
wire x_30636;
wire x_30637;
wire x_30638;
wire x_30639;
wire x_30640;
wire x_30641;
wire x_30642;
wire x_30643;
wire x_30644;
wire x_30645;
wire x_30646;
wire x_30647;
wire x_30648;
wire x_30649;
wire x_30650;
wire x_30651;
wire x_30652;
wire x_30653;
wire x_30654;
wire x_30655;
wire x_30656;
wire x_30657;
wire x_30658;
wire x_30659;
wire x_30660;
wire x_30661;
wire x_30662;
wire x_30663;
wire x_30664;
wire x_30665;
wire x_30666;
wire x_30667;
wire x_30668;
wire x_30669;
wire x_30670;
wire x_30671;
wire x_30672;
wire x_30673;
wire x_30674;
wire x_30675;
wire x_30676;
wire x_30677;
wire x_30678;
wire x_30679;
wire x_30680;
wire x_30681;
wire x_30682;
wire x_30683;
wire x_30684;
wire x_30685;
wire x_30686;
wire x_30687;
wire x_30688;
wire x_30689;
wire x_30690;
wire x_30691;
wire x_30692;
wire x_30693;
wire x_30694;
wire x_30695;
wire x_30696;
wire x_30697;
wire x_30698;
wire x_30699;
wire x_30700;
wire x_30701;
wire x_30702;
wire x_30703;
wire x_30704;
wire x_30705;
wire x_30706;
wire x_30707;
wire x_30708;
wire x_30709;
wire x_30710;
wire x_30711;
wire x_30712;
wire x_30713;
wire x_30714;
wire x_30715;
wire x_30716;
wire x_30717;
wire x_30718;
wire x_30719;
wire x_30720;
wire x_30721;
wire x_30722;
wire x_30723;
wire x_30724;
wire x_30725;
wire x_30726;
wire x_30727;
wire x_30728;
wire x_30729;
wire x_30730;
wire x_30731;
wire x_30732;
wire x_30733;
wire x_30734;
wire x_30735;
wire x_30736;
wire x_30737;
wire x_30738;
wire x_30739;
wire x_30740;
wire x_30741;
wire x_30742;
wire x_30743;
wire x_30744;
wire x_30745;
wire x_30746;
wire x_30747;
wire x_30748;
wire x_30749;
wire x_30750;
wire x_30751;
wire x_30752;
wire x_30753;
wire x_30754;
wire x_30755;
wire x_30756;
wire x_30757;
wire x_30758;
wire x_30759;
wire x_30760;
wire x_30761;
wire x_30762;
wire x_30763;
wire x_30764;
wire x_30765;
wire x_30766;
wire x_30767;
wire x_30768;
wire x_30769;
wire x_30770;
wire x_30771;
wire x_30772;
wire x_30773;
wire x_30774;
wire x_30775;
wire x_30776;
wire x_30777;
wire x_30778;
wire x_30779;
wire x_30780;
wire x_30781;
wire x_30782;
wire x_30783;
wire x_30784;
wire x_30785;
wire x_30786;
wire x_30787;
wire x_30788;
wire x_30789;
wire x_30790;
wire x_30791;
wire x_30792;
wire x_30793;
wire x_30794;
wire x_30795;
wire x_30796;
wire x_30797;
wire x_30798;
wire x_30799;
wire x_30800;
wire x_30801;
wire x_30802;
wire x_30803;
wire x_30804;
wire x_30805;
wire x_30806;
wire x_30807;
wire x_30808;
wire x_30809;
wire x_30810;
wire x_30811;
wire x_30812;
wire x_30813;
wire x_30814;
wire x_30815;
wire x_30816;
wire x_30817;
wire x_30818;
wire x_30819;
wire x_30820;
wire x_30821;
wire x_30822;
wire x_30823;
wire x_30824;
wire x_30825;
wire x_30826;
wire x_30827;
wire x_30828;
wire x_30829;
wire x_30830;
wire x_30831;
wire x_30832;
wire x_30833;
wire x_30834;
wire x_30835;
wire x_30836;
wire x_30837;
wire x_30838;
wire x_30839;
wire x_30840;
wire x_30841;
wire x_30842;
wire x_30843;
wire x_30844;
wire x_30845;
wire x_30846;
wire x_30847;
wire x_30848;
wire x_30849;
wire x_30850;
wire x_30851;
wire x_30852;
wire x_30853;
wire x_30854;
wire x_30855;
wire x_30856;
wire x_30857;
wire x_30858;
wire x_30859;
wire x_30860;
wire x_30861;
wire x_30862;
wire x_30863;
wire x_30864;
wire x_30865;
wire x_30866;
wire x_30867;
wire x_30868;
wire x_30869;
wire x_30870;
wire x_30871;
wire x_30872;
wire x_30873;
wire x_30874;
wire x_30875;
wire x_30876;
wire x_30877;
wire x_30878;
wire x_30879;
wire x_30880;
wire x_30881;
wire x_30882;
wire x_30883;
wire x_30884;
wire x_30885;
wire x_30886;
wire x_30887;
wire x_30888;
wire x_30889;
wire x_30890;
wire x_30891;
wire x_30892;
wire x_30893;
wire x_30894;
wire x_30895;
wire x_30896;
wire x_30897;
wire x_30898;
wire x_30899;
wire x_30900;
wire x_30901;
wire x_30902;
wire x_30903;
wire x_30904;
wire x_30905;
wire x_30906;
wire x_30907;
wire x_30908;
wire x_30909;
wire x_30910;
wire x_30911;
wire x_30912;
wire x_30913;
wire x_30914;
wire x_30915;
wire x_30916;
wire x_30917;
wire x_30918;
wire x_30919;
wire x_30920;
wire x_30921;
wire x_30922;
wire x_30923;
wire x_30924;
wire x_30925;
wire x_30926;
wire x_30927;
wire x_30928;
wire x_30929;
wire x_30930;
wire x_30931;
wire x_30932;
wire x_30933;
wire x_30934;
wire x_30935;
wire x_30936;
wire x_30937;
wire x_30938;
wire x_30939;
wire x_30940;
wire x_30941;
wire x_30942;
wire x_30943;
wire x_30944;
wire x_30945;
wire x_30946;
wire x_30947;
wire x_30948;
wire x_30949;
wire x_30950;
wire x_30951;
wire x_30952;
wire x_30953;
wire x_30954;
wire x_30955;
wire x_30956;
wire x_30957;
wire x_30958;
wire x_30959;
wire x_30960;
wire x_30961;
wire x_30962;
wire x_30963;
wire x_30964;
wire x_30965;
wire x_30966;
wire x_30967;
wire x_30968;
wire x_30969;
wire x_30970;
wire x_30971;
wire x_30972;
wire x_30973;
wire x_30974;
wire x_30975;
wire x_30976;
wire x_30977;
wire x_30978;
wire x_30979;
wire x_30980;
wire x_30981;
wire x_30982;
wire x_30983;
wire x_30984;
wire x_30985;
wire x_30986;
wire x_30987;
wire x_30988;
wire x_30989;
wire x_30990;
wire x_30991;
wire x_30992;
wire x_30993;
wire x_30994;
wire x_30995;
wire x_30996;
wire x_30997;
wire x_30998;
wire x_30999;
wire x_31000;
wire x_31001;
wire x_31002;
wire x_31003;
wire x_31004;
wire x_31005;
wire x_31006;
wire x_31007;
wire x_31008;
wire x_31009;
wire x_31010;
wire x_31011;
wire x_31012;
wire x_31013;
wire x_31014;
wire x_31015;
wire x_31016;
wire x_31017;
wire x_31018;
wire x_31019;
wire x_31020;
wire x_31021;
wire x_31022;
wire x_31023;
wire x_31024;
wire x_31025;
wire x_31026;
wire x_31027;
wire x_31028;
wire x_31029;
wire x_31030;
wire x_31031;
wire x_31032;
wire x_31033;
wire x_31034;
wire x_31035;
wire x_31036;
wire x_31037;
wire x_31038;
wire x_31039;
wire x_31040;
wire x_31041;
wire x_31042;
wire x_31043;
wire x_31044;
wire x_31045;
wire x_31046;
wire x_31047;
wire x_31048;
wire x_31049;
wire x_31050;
wire x_31051;
wire x_31052;
wire x_31053;
wire x_31054;
wire x_31055;
wire x_31056;
wire x_31057;
wire x_31058;
wire x_31059;
wire x_31060;
wire x_31061;
wire x_31062;
wire x_31063;
wire x_31064;
wire x_31065;
wire x_31066;
wire x_31067;
wire x_31068;
wire x_31069;
wire x_31070;
wire x_31071;
wire x_31072;
wire x_31073;
wire x_31074;
wire x_31075;
wire x_31076;
wire x_31077;
wire x_31078;
wire x_31079;
wire x_31080;
wire x_31081;
wire x_31082;
wire x_31083;
wire x_31084;
wire x_31085;
wire x_31086;
wire x_31087;
wire x_31088;
wire x_31089;
wire x_31090;
wire x_31091;
wire x_31092;
wire x_31093;
wire x_31094;
wire x_31095;
wire x_31096;
wire x_31097;
wire x_31098;
wire x_31099;
wire x_31100;
wire x_31101;
wire x_31102;
wire x_31103;
wire x_31104;
wire x_31105;
wire x_31106;
wire x_31107;
wire x_31108;
wire x_31109;
wire x_31110;
wire x_31111;
wire x_31112;
wire x_31113;
wire x_31114;
wire x_31115;
wire x_31116;
wire x_31117;
wire x_31118;
wire x_31119;
wire x_31120;
wire x_31121;
wire x_31122;
wire x_31123;
wire x_31124;
wire x_31125;
wire x_31126;
wire x_31127;
wire x_31128;
wire x_31129;
wire x_31130;
wire x_31131;
wire x_31132;
wire x_31133;
wire x_31134;
wire x_31135;
wire x_31136;
wire x_31137;
wire x_31138;
wire x_31139;
wire x_31140;
wire x_31141;
wire x_31142;
wire x_31143;
wire x_31144;
wire x_31145;
wire x_31146;
wire x_31147;
wire x_31148;
wire x_31149;
wire x_31150;
wire x_31151;
wire x_31152;
wire x_31153;
wire x_31154;
wire x_31155;
wire x_31156;
wire x_31157;
wire x_31158;
wire x_31159;
wire x_31160;
wire x_31161;
wire x_31162;
wire x_31163;
wire x_31164;
wire x_31165;
wire x_31166;
wire x_31167;
wire x_31168;
wire x_31169;
wire x_31170;
wire x_31171;
wire x_31172;
wire x_31173;
wire x_31174;
wire x_31175;
wire x_31176;
wire x_31177;
wire x_31178;
wire x_31179;
wire x_31180;
wire x_31181;
wire x_31182;
wire x_31183;
wire x_31184;
wire x_31185;
wire x_31186;
wire x_31187;
wire x_31188;
wire x_31189;
wire x_31190;
wire x_31191;
wire x_31192;
wire x_31193;
wire x_31194;
wire x_31195;
wire x_31196;
wire x_31197;
wire x_31198;
wire x_31199;
wire x_31200;
wire x_31201;
wire x_31202;
wire x_31203;
wire x_31204;
wire x_31205;
wire x_31206;
wire x_31207;
wire x_31208;
wire x_31209;
wire x_31210;
wire x_31211;
wire x_31212;
wire x_31213;
wire x_31214;
wire x_31215;
wire x_31216;
wire x_31217;
wire x_31218;
wire x_31219;
wire x_31220;
wire x_31221;
wire x_31222;
wire x_31223;
wire x_31224;
wire x_31225;
wire x_31226;
wire x_31227;
wire x_31228;
wire x_31229;
wire x_31230;
wire x_31231;
wire x_31232;
wire x_31233;
wire x_31234;
wire x_31235;
wire x_31236;
wire x_31237;
wire x_31238;
wire x_31239;
wire x_31240;
wire x_31241;
wire x_31242;
wire x_31243;
wire x_31244;
wire x_31245;
wire x_31246;
wire x_31247;
wire x_31248;
wire x_31249;
wire x_31250;
wire x_31251;
wire x_31252;
wire x_31253;
wire x_31254;
wire x_31255;
wire x_31256;
wire x_31257;
wire x_31258;
wire x_31259;
wire x_31260;
wire x_31261;
wire x_31262;
wire x_31263;
wire x_31264;
wire x_31265;
wire x_31266;
wire x_31267;
wire x_31268;
wire x_31269;
wire x_31270;
wire x_31271;
wire x_31272;
wire x_31273;
wire x_31274;
wire x_31275;
wire x_31276;
wire x_31277;
wire x_31278;
wire x_31279;
wire x_31280;
wire x_31281;
wire x_31282;
wire x_31283;
wire x_31284;
wire x_31285;
wire x_31286;
wire x_31287;
wire x_31288;
wire x_31289;
wire x_31290;
wire x_31291;
wire x_31292;
wire x_31293;
wire x_31294;
wire x_31295;
wire x_31296;
wire x_31297;
wire x_31298;
wire x_31299;
wire x_31300;
wire x_31301;
wire x_31302;
wire x_31303;
wire x_31304;
wire x_31305;
wire x_31306;
wire x_31307;
wire x_31308;
wire x_31309;
wire x_31310;
wire x_31311;
wire x_31312;
wire x_31313;
wire x_31314;
wire x_31315;
wire x_31316;
wire x_31317;
wire x_31318;
wire x_31319;
wire x_31320;
wire x_31321;
wire x_31322;
wire x_31323;
wire x_31324;
wire x_31325;
wire x_31326;
wire x_31327;
wire x_31328;
wire x_31329;
wire x_31330;
wire x_31331;
wire x_31332;
wire x_31333;
wire x_31334;
wire x_31335;
wire x_31336;
wire x_31337;
wire x_31338;
wire x_31339;
wire x_31340;
wire x_31341;
wire x_31342;
wire x_31343;
wire x_31344;
wire x_31345;
wire x_31346;
wire x_31347;
wire x_31348;
wire x_31349;
wire x_31350;
wire x_31351;
wire x_31352;
wire x_31353;
wire x_31354;
wire x_31355;
wire x_31356;
wire x_31357;
wire x_31358;
wire x_31359;
wire x_31360;
wire x_31361;
wire x_31362;
wire x_31363;
wire x_31364;
wire x_31365;
wire x_31366;
wire x_31367;
wire x_31368;
wire x_31369;
wire x_31370;
wire x_31371;
wire x_31372;
wire x_31373;
wire x_31374;
wire x_31375;
wire x_31376;
wire x_31377;
wire x_31378;
wire x_31379;
wire x_31380;
wire x_31381;
wire x_31382;
wire x_31383;
wire x_31384;
wire x_31385;
wire x_31386;
wire x_31387;
wire x_31388;
wire x_31389;
wire x_31390;
wire x_31391;
wire x_31392;
wire x_31393;
wire x_31394;
wire x_31395;
wire x_31396;
wire x_31397;
wire x_31398;
wire x_31399;
wire x_31400;
wire x_31401;
wire x_31402;
wire x_31403;
wire x_31404;
wire x_31405;
wire x_31406;
wire x_31407;
wire x_31408;
wire x_31409;
wire x_31410;
wire x_31411;
wire x_31412;
wire x_31413;
wire x_31414;
wire x_31415;
wire x_31416;
wire x_31417;
wire x_31418;
wire x_31419;
wire x_31420;
wire x_31421;
wire x_31422;
wire x_31423;
wire x_31424;
wire x_31425;
wire x_31426;
wire x_31427;
wire x_31428;
wire x_31429;
wire x_31430;
wire x_31431;
wire x_31432;
wire x_31433;
wire x_31434;
wire x_31435;
wire x_31436;
wire x_31437;
wire x_31438;
wire x_31439;
wire x_31440;
wire x_31441;
wire x_31442;
wire x_31443;
wire x_31444;
wire x_31445;
wire x_31446;
wire x_31447;
wire x_31448;
wire x_31449;
wire x_31450;
wire x_31451;
wire x_31452;
wire x_31453;
wire x_31454;
wire x_31455;
wire x_31456;
wire x_31457;
wire x_31458;
wire x_31459;
wire x_31460;
wire x_31461;
wire x_31462;
wire x_31463;
wire x_31464;
wire x_31465;
wire x_31466;
wire x_31467;
wire x_31468;
wire x_31469;
wire x_31470;
wire x_31471;
wire x_31472;
wire x_31473;
wire x_31474;
wire x_31475;
wire x_31476;
wire x_31477;
wire x_31478;
wire x_31479;
wire x_31480;
wire x_31481;
wire x_31482;
wire x_31483;
wire x_31484;
wire x_31485;
wire x_31486;
wire x_31487;
wire x_31488;
wire x_31489;
wire x_31490;
wire x_31491;
wire x_31492;
wire x_31493;
wire x_31494;
wire x_31495;
wire x_31496;
wire x_31497;
wire x_31498;
wire x_31499;
wire x_31500;
wire x_31501;
wire x_31502;
wire x_31503;
wire x_31504;
wire x_31505;
wire x_31506;
wire x_31507;
wire x_31508;
wire x_31509;
wire x_31510;
wire x_31511;
wire x_31512;
wire x_31513;
wire x_31514;
wire x_31515;
wire x_31516;
wire x_31517;
wire x_31518;
wire x_31519;
wire x_31520;
wire x_31521;
wire x_31522;
wire x_31523;
wire x_31524;
wire x_31525;
wire x_31526;
wire x_31527;
wire x_31528;
wire x_31529;
wire x_31530;
wire x_31531;
wire x_31532;
wire x_31533;
wire x_31534;
wire x_31535;
wire x_31536;
wire x_31537;
wire x_31538;
wire x_31539;
wire x_31540;
wire x_31541;
wire x_31542;
wire x_31543;
wire x_31544;
wire x_31545;
wire x_31546;
wire x_31547;
wire x_31548;
wire x_31549;
wire x_31550;
wire x_31551;
wire x_31552;
wire x_31553;
wire x_31554;
wire x_31555;
wire x_31556;
wire x_31557;
wire x_31558;
wire x_31559;
wire x_31560;
wire x_31561;
wire x_31562;
wire x_31563;
wire x_31564;
wire x_31565;
wire x_31566;
wire x_31567;
wire x_31568;
wire x_31569;
wire x_31570;
wire x_31571;
wire x_31572;
wire x_31573;
wire x_31574;
wire x_31575;
wire x_31576;
wire x_31577;
wire x_31578;
wire x_31579;
wire x_31580;
wire x_31581;
wire x_31582;
wire x_31583;
wire x_31584;
wire x_31585;
wire x_31586;
wire x_31587;
wire x_31588;
wire x_31589;
wire x_31590;
wire x_31591;
wire x_31592;
wire x_31593;
wire x_31594;
wire x_31595;
wire x_31596;
wire x_31597;
wire x_31598;
wire x_31599;
wire x_31600;
wire x_31601;
wire x_31602;
wire x_31603;
wire x_31604;
wire x_31605;
wire x_31606;
wire x_31607;
wire x_31608;
wire x_31609;
wire x_31610;
wire x_31611;
wire x_31612;
wire x_31613;
wire x_31614;
wire x_31615;
wire x_31616;
wire x_31617;
wire x_31618;
wire x_31619;
wire x_31620;
wire x_31621;
wire x_31622;
wire x_31623;
wire x_31624;
wire x_31625;
wire x_31626;
wire x_31627;
wire x_31628;
wire x_31629;
wire x_31630;
wire x_31631;
wire x_31632;
wire x_31633;
wire x_31634;
wire x_31635;
wire x_31636;
wire x_31637;
wire x_31638;
wire x_31639;
wire x_31640;
wire x_31641;
wire x_31642;
wire x_31643;
wire x_31644;
wire x_31645;
wire x_31646;
wire x_31647;
wire x_31648;
wire x_31649;
wire x_31650;
wire x_31651;
wire x_31652;
wire x_31653;
wire x_31654;
wire x_31655;
wire x_31656;
wire x_31657;
wire x_31658;
wire x_31659;
wire x_31660;
wire x_31661;
wire x_31662;
wire x_31663;
wire x_31664;
wire x_31665;
wire x_31666;
wire x_31667;
wire x_31668;
wire x_31669;
wire x_31670;
wire x_31671;
wire x_31672;
wire x_31673;
wire x_31674;
wire x_31675;
wire x_31676;
wire x_31677;
wire x_31678;
wire x_31679;
wire x_31680;
wire x_31681;
wire x_31682;
wire x_31683;
wire x_31684;
wire x_31685;
wire x_31686;
wire x_31687;
wire x_31688;
wire x_31689;
wire x_31690;
wire x_31691;
wire x_31692;
wire x_31693;
wire x_31694;
wire x_31695;
wire x_31696;
wire x_31697;
wire x_31698;
wire x_31699;
wire x_31700;
wire x_31701;
wire x_31702;
wire x_31703;
wire x_31704;
wire x_31705;
wire x_31706;
wire x_31707;
wire x_31708;
wire x_31709;
wire x_31710;
wire x_31711;
wire x_31712;
wire x_31713;
wire x_31714;
wire x_31715;
wire x_31716;
wire x_31717;
wire x_31718;
wire x_31719;
wire x_31720;
wire x_31721;
wire x_31722;
wire x_31723;
wire x_31724;
wire x_31725;
wire x_31726;
wire x_31727;
wire x_31728;
wire x_31729;
wire x_31730;
wire x_31731;
wire x_31732;
wire x_31733;
wire x_31734;
wire x_31735;
wire x_31736;
wire x_31737;
wire x_31738;
wire x_31739;
wire x_31740;
wire x_31741;
wire x_31742;
wire x_31743;
wire x_31744;
wire x_31745;
wire x_31746;
wire x_31747;
wire x_31748;
wire x_31749;
wire x_31750;
wire x_31751;
wire x_31752;
wire x_31753;
wire x_31754;
wire x_31755;
wire x_31756;
wire x_31757;
wire x_31758;
wire x_31759;
wire x_31760;
wire x_31761;
wire x_31762;
wire x_31763;
wire x_31764;
wire x_31765;
wire x_31766;
wire x_31767;
wire x_31768;
wire x_31769;
wire x_31770;
wire x_31771;
wire x_31772;
wire x_31773;
wire x_31774;
wire x_31775;
wire x_31776;
wire x_31777;
wire x_31778;
wire x_31779;
wire x_31780;
wire x_31781;
wire x_31782;
wire x_31783;
wire x_31784;
wire x_31785;
wire x_31786;
wire x_31787;
wire x_31788;
wire x_31789;
wire x_31790;
wire x_31791;
wire x_31792;
wire x_31793;
wire x_31794;
wire x_31795;
wire x_31796;
wire x_31797;
wire x_31798;
wire x_31799;
wire x_31800;
wire x_31801;
wire x_31802;
wire x_31803;
wire x_31804;
wire x_31805;
wire x_31806;
wire x_31807;
wire x_31808;
wire x_31809;
wire x_31810;
wire x_31811;
wire x_31812;
wire x_31813;
wire x_31814;
wire x_31815;
wire x_31816;
wire x_31817;
wire x_31818;
wire x_31819;
wire x_31820;
wire x_31821;
wire x_31822;
wire x_31823;
wire x_31824;
wire x_31825;
wire x_31826;
wire x_31827;
wire x_31828;
wire x_31829;
wire x_31830;
wire x_31831;
wire x_31832;
wire x_31833;
wire x_31834;
wire x_31835;
wire x_31836;
wire x_31837;
wire x_31838;
wire x_31839;
wire x_31840;
wire x_31841;
wire x_31842;
wire x_31843;
wire x_31844;
wire x_31845;
wire x_31846;
wire x_31847;
wire x_31848;
wire x_31849;
wire x_31850;
wire x_31851;
wire x_31852;
wire x_31853;
wire x_31854;
wire x_31855;
wire x_31856;
wire x_31857;
wire x_31858;
wire x_31859;
wire x_31860;
wire x_31861;
wire x_31862;
wire x_31863;
wire x_31864;
wire x_31865;
wire x_31866;
wire x_31867;
wire x_31868;
wire x_31869;
wire x_31870;
wire x_31871;
wire x_31872;
wire x_31873;
wire x_31874;
wire x_31875;
wire x_31876;
wire x_31877;
wire x_31878;
wire x_31879;
wire x_31880;
wire x_31881;
wire x_31882;
wire x_31883;
wire x_31884;
wire x_31885;
wire x_31886;
wire x_31887;
wire x_31888;
wire x_31889;
wire x_31890;
wire x_31891;
wire x_31892;
wire x_31893;
wire x_31894;
wire x_31895;
wire x_31896;
wire x_31897;
wire x_31898;
wire x_31899;
wire x_31900;
wire x_31901;
wire x_31902;
wire x_31903;
wire x_31904;
wire x_31905;
wire x_31906;
wire x_31907;
wire x_31908;
wire x_31909;
wire x_31910;
wire x_31911;
wire x_31912;
wire x_31913;
wire x_31914;
wire x_31915;
wire x_31916;
wire x_31917;
wire x_31918;
wire x_31919;
wire x_31920;
wire x_31921;
wire x_31922;
wire x_31923;
wire x_31924;
wire x_31925;
wire x_31926;
wire x_31927;
wire x_31928;
wire x_31929;
wire x_31930;
wire x_31931;
wire x_31932;
wire x_31933;
wire x_31934;
wire x_31935;
wire x_31936;
wire x_31937;
wire x_31938;
wire x_31939;
wire x_31940;
wire x_31941;
wire x_31942;
wire x_31943;
wire x_31944;
wire x_31945;
wire x_31946;
wire x_31947;
wire x_31948;
wire x_31949;
wire x_31950;
wire x_31951;
wire x_31952;
wire x_31953;
wire x_31954;
wire x_31955;
wire x_31956;
wire x_31957;
wire x_31958;
wire x_31959;
wire x_31960;
wire x_31961;
wire x_31962;
wire x_31963;
wire x_31964;
wire x_31965;
wire x_31966;
wire x_31967;
wire x_31968;
wire x_31969;
wire x_31970;
wire x_31971;
wire x_31972;
wire x_31973;
wire x_31974;
wire x_31975;
wire x_31976;
wire x_31977;
wire x_31978;
wire x_31979;
wire x_31980;
wire x_31981;
wire x_31982;
wire x_31983;
wire x_31984;
wire x_31985;
wire x_31986;
wire x_31987;
wire x_31988;
wire x_31989;
wire x_31990;
wire x_31991;
wire x_31992;
wire x_31993;
wire x_31994;
wire x_31995;
wire x_31996;
wire x_31997;
wire x_31998;
wire x_31999;
wire x_32000;
wire x_32001;
wire x_32002;
wire x_32003;
wire x_32004;
wire x_32005;
wire x_32006;
wire x_32007;
wire x_32008;
wire x_32009;
wire x_32010;
wire x_32011;
wire x_32012;
wire x_32013;
wire x_32014;
wire x_32015;
wire x_32016;
wire x_32017;
wire x_32018;
wire x_32019;
wire x_32020;
wire x_32021;
wire x_32022;
wire x_32023;
wire x_32024;
wire x_32025;
wire x_32026;
wire x_32027;
wire x_32028;
wire x_32029;
wire x_32030;
wire x_32031;
wire x_32032;
wire x_32033;
wire x_32034;
wire x_32035;
wire x_32036;
wire x_32037;
wire x_32038;
wire x_32039;
wire x_32040;
wire x_32041;
wire x_32042;
wire x_32043;
wire x_32044;
wire x_32045;
wire x_32046;
wire x_32047;
wire x_32048;
wire x_32049;
wire x_32050;
wire x_32051;
wire x_32052;
wire x_32053;
wire x_32054;
wire x_32055;
wire x_32056;
wire x_32057;
wire x_32058;
wire x_32059;
wire x_32060;
wire x_32061;
wire x_32062;
wire x_32063;
wire x_32064;
wire x_32065;
wire x_32066;
wire x_32067;
wire x_32068;
wire x_32069;
wire x_32070;
wire x_32071;
wire x_32072;
wire x_32073;
wire x_32074;
wire x_32075;
wire x_32076;
wire x_32077;
wire x_32078;
wire x_32079;
wire x_32080;
wire x_32081;
wire x_32082;
wire x_32083;
wire x_32084;
wire x_32085;
wire x_32086;
wire x_32087;
wire x_32088;
wire x_32089;
wire x_32090;
wire x_32091;
wire x_32092;
wire x_32093;
wire x_32094;
wire x_32095;
wire x_32096;
wire x_32097;
wire x_32098;
wire x_32099;
wire x_32100;
wire x_32101;
wire x_32102;
wire x_32103;
wire x_32104;
wire x_32105;
wire x_32106;
wire x_32107;
wire x_32108;
wire x_32109;
wire x_32110;
wire x_32111;
wire x_32112;
wire x_32113;
wire x_32114;
wire x_32115;
wire x_32116;
wire x_32117;
wire x_32118;
wire x_32119;
wire x_32120;
wire x_32121;
wire x_32122;
wire x_32123;
wire x_32124;
wire x_32125;
wire x_32126;
wire x_32127;
wire x_32128;
wire x_32129;
wire x_32130;
wire x_32131;
wire x_32132;
wire x_32133;
wire x_32134;
wire x_32135;
wire x_32136;
wire x_32137;
wire x_32138;
wire x_32139;
wire x_32140;
wire x_32141;
wire x_32142;
wire x_32143;
wire x_32144;
wire x_32145;
wire x_32146;
wire x_32147;
wire x_32148;
wire x_32149;
wire x_32150;
wire x_32151;
wire x_32152;
wire x_32153;
wire x_32154;
wire x_32155;
wire x_32156;
wire x_32157;
wire x_32158;
wire x_32159;
wire x_32160;
wire x_32161;
wire x_32162;
wire x_32163;
wire x_32164;
wire x_32165;
wire x_32166;
wire x_32167;
wire x_32168;
wire x_32169;
wire x_32170;
wire x_32171;
wire x_32172;
wire x_32173;
wire x_32174;
wire x_32175;
wire x_32176;
wire x_32177;
wire x_32178;
wire x_32179;
wire x_32180;
wire x_32181;
wire x_32182;
wire x_32183;
wire x_32184;
wire x_32185;
wire x_32186;
wire x_32187;
wire x_32188;
wire x_32189;
wire x_32190;
wire x_32191;
wire x_32192;
wire x_32193;
wire x_32194;
wire x_32195;
wire x_32196;
wire x_32197;
wire x_32198;
wire x_32199;
wire x_32200;
wire x_32201;
wire x_32202;
wire x_32203;
wire x_32204;
wire x_32205;
wire x_32206;
wire x_32207;
wire x_32208;
wire x_32209;
wire x_32210;
wire x_32211;
wire x_32212;
wire x_32213;
wire x_32214;
wire x_32215;
wire x_32216;
wire x_32217;
wire x_32218;
wire x_32219;
wire x_32220;
wire x_32221;
wire x_32222;
wire x_32223;
wire x_32224;
wire x_32225;
wire x_32226;
wire x_32227;
wire x_32228;
wire x_32229;
wire x_32230;
wire x_32231;
wire x_32232;
wire x_32233;
wire x_32234;
wire x_32235;
wire x_32236;
wire x_32237;
wire x_32238;
wire x_32239;
wire x_32240;
wire x_32241;
wire x_32242;
wire x_32243;
wire x_32244;
wire x_32245;
wire x_32246;
wire x_32247;
wire x_32248;
wire x_32249;
wire x_32250;
wire x_32251;
wire x_32252;
wire x_32253;
wire x_32254;
wire x_32255;
wire x_32256;
wire x_32257;
wire x_32258;
wire x_32259;
wire x_32260;
wire x_32261;
wire x_32262;
wire x_32263;
wire x_32264;
wire x_32265;
wire x_32266;
wire x_32267;
wire x_32268;
wire x_32269;
wire x_32270;
wire x_32271;
wire x_32272;
wire x_32273;
wire x_32274;
wire x_32275;
wire x_32276;
wire x_32277;
wire x_32278;
wire x_32279;
wire x_32280;
wire x_32281;
wire x_32282;
wire x_32283;
wire x_32284;
wire x_32285;
wire x_32286;
wire x_32287;
wire x_32288;
wire x_32289;
wire x_32290;
wire x_32291;
wire x_32292;
wire x_32293;
wire x_32294;
wire x_32295;
wire x_32296;
wire x_32297;
wire x_32298;
wire x_32299;
wire x_32300;
wire x_32301;
wire x_32302;
wire x_32303;
wire x_32304;
wire x_32305;
wire x_32306;
wire x_32307;
wire x_32308;
wire x_32309;
wire x_32310;
wire x_32311;
wire x_32312;
wire x_32313;
wire x_32314;
wire x_32315;
wire x_32316;
wire x_32317;
wire x_32318;
wire x_32319;
wire x_32320;
wire x_32321;
wire x_32322;
wire x_32323;
wire x_32324;
wire x_32325;
wire x_32326;
wire x_32327;
wire x_32328;
wire x_32329;
wire x_32330;
wire x_32331;
wire x_32332;
wire x_32333;
wire x_32334;
wire x_32335;
wire x_32336;
wire x_32337;
wire x_32338;
wire x_32339;
wire x_32340;
wire x_32341;
wire x_32342;
wire x_32343;
wire x_32344;
wire x_32345;
wire x_32346;
wire x_32347;
wire x_32348;
wire x_32349;
wire x_32350;
wire x_32351;
wire x_32352;
wire x_32353;
wire x_32354;
wire x_32355;
wire x_32356;
wire x_32357;
wire x_32358;
wire x_32359;
wire x_32360;
wire x_32361;
wire x_32362;
wire x_32363;
wire x_32364;
wire x_32365;
wire x_32366;
wire x_32367;
wire x_32368;
wire x_32369;
wire x_32370;
wire x_32371;
wire x_32372;
wire x_32373;
wire x_32374;
wire x_32375;
wire x_32376;
wire x_32377;
wire x_32378;
wire x_32379;
wire x_32380;
wire x_32381;
wire x_32382;
wire x_32383;
wire x_32384;
wire x_32385;
wire x_32386;
wire x_32387;
wire x_32388;
wire x_32389;
wire x_32390;
wire x_32391;
wire x_32392;
wire x_32393;
wire x_32394;
wire x_32395;
wire x_32396;
wire x_32397;
wire x_32398;
wire x_32399;
wire x_32400;
wire x_32401;
wire x_32402;
wire x_32403;
wire x_32404;
wire x_32405;
wire x_32406;
wire x_32407;
wire x_32408;
wire x_32409;
wire x_32410;
wire x_32411;
wire x_32412;
wire x_32413;
wire x_32414;
wire x_32415;
wire x_32416;
wire x_32417;
wire x_32418;
wire x_32419;
wire x_32420;
wire x_32421;
wire x_32422;
wire x_32423;
wire x_32424;
wire x_32425;
wire x_32426;
wire x_32427;
wire x_32428;
wire x_32429;
wire x_32430;
wire x_32431;
wire x_32432;
wire x_32433;
wire x_32434;
wire x_32435;
wire x_32436;
wire x_32437;
wire x_32438;
wire x_32439;
wire x_32440;
wire x_32441;
wire x_32442;
wire x_32443;
wire x_32444;
wire x_32445;
wire x_32446;
wire x_32447;
wire x_32448;
wire x_32449;
wire x_32450;
wire x_32451;
wire x_32452;
wire x_32453;
wire x_32454;
wire x_32455;
wire x_32456;
wire x_32457;
wire x_32458;
wire x_32459;
wire x_32460;
wire x_32461;
wire x_32462;
wire x_32463;
wire x_32464;
wire x_32465;
wire x_32466;
wire x_32467;
wire x_32468;
wire x_32469;
wire x_32470;
wire x_32471;
wire x_32472;
wire x_32473;
wire x_32474;
wire x_32475;
wire x_32476;
wire x_32477;
wire x_32478;
wire x_32479;
wire x_32480;
wire x_32481;
wire x_32482;
wire x_32483;
wire x_32484;
wire x_32485;
wire x_32486;
wire x_32487;
wire x_32488;
wire x_32489;
wire x_32490;
wire x_32491;
wire x_32492;
wire x_32493;
wire x_32494;
wire x_32495;
wire x_32496;
wire x_32497;
wire x_32498;
wire x_32499;
wire x_32500;
wire x_32501;
wire x_32502;
wire x_32503;
wire x_32504;
wire x_32505;
wire x_32506;
wire x_32507;
wire x_32508;
wire x_32509;
wire x_32510;
wire x_32511;
wire x_32512;
wire x_32513;
wire x_32514;
wire x_32515;
wire x_32516;
wire x_32517;
wire x_32518;
wire x_32519;
wire x_32520;
wire x_32521;
wire x_32522;
wire x_32523;
wire x_32524;
wire x_32525;
wire x_32526;
wire x_32527;
wire x_32528;
wire x_32529;
wire x_32530;
wire x_32531;
wire x_32532;
wire x_32533;
wire x_32534;
wire x_32535;
wire x_32536;
wire x_32537;
wire x_32538;
wire x_32539;
wire x_32540;
wire x_32541;
wire x_32542;
wire x_32543;
wire x_32544;
wire x_32545;
wire x_32546;
wire x_32547;
wire x_32548;
wire x_32549;
wire x_32550;
wire x_32551;
wire x_32552;
wire x_32553;
wire x_32554;
wire x_32555;
wire x_32556;
wire x_32557;
wire x_32558;
wire x_32559;
wire x_32560;
wire x_32561;
wire x_32562;
wire x_32563;
wire x_32564;
wire x_32565;
wire x_32566;
wire x_32567;
wire x_32568;
wire x_32569;
wire x_32570;
wire x_32571;
wire x_32572;
wire x_32573;
wire x_32574;
wire x_32575;
wire x_32576;
wire x_32577;
wire x_32578;
wire x_32579;
wire x_32580;
wire x_32581;
wire x_32582;
wire x_32583;
wire x_32584;
wire x_32585;
wire x_32586;
wire x_32587;
wire x_32588;
wire x_32589;
wire x_32590;
wire x_32591;
wire x_32592;
wire x_32593;
wire x_32594;
wire x_32595;
wire x_32596;
wire x_32597;
wire x_32598;
wire x_32599;
wire x_32600;
wire x_32601;
wire x_32602;
wire x_32603;
wire x_32604;
wire x_32605;
wire x_32606;
wire x_32607;
wire x_32608;
wire x_32609;
wire x_32610;
wire x_32611;
wire x_32612;
wire x_32613;
wire x_32614;
wire x_32615;
wire x_32616;
wire x_32617;
wire x_32618;
wire x_32619;
wire x_32620;
wire x_32621;
wire x_32622;
wire x_32623;
wire x_32624;
wire x_32625;
wire x_32626;
wire x_32627;
wire x_32628;
wire x_32629;
wire x_32630;
wire x_32631;
wire x_32632;
wire x_32633;
wire x_32634;
wire x_32635;
wire x_32636;
wire x_32637;
wire x_32638;
wire x_32639;
wire x_32640;
wire x_32641;
wire x_32642;
wire x_32643;
wire x_32644;
wire x_32645;
wire x_32646;
wire x_32647;
wire x_32648;
wire x_32649;
wire x_32650;
wire x_32651;
wire x_32652;
wire x_32653;
wire x_32654;
wire x_32655;
wire x_32656;
wire x_32657;
wire x_32658;
wire x_32659;
wire x_32660;
wire x_32661;
wire x_32662;
wire x_32663;
wire x_32664;
wire x_32665;
wire x_32666;
wire x_32667;
wire x_32668;
wire x_32669;
wire x_32670;
wire x_32671;
wire x_32672;
wire x_32673;
wire x_32674;
wire x_32675;
wire x_32676;
wire x_32677;
wire x_32678;
wire x_32679;
wire x_32680;
wire x_32681;
wire x_32682;
wire x_32683;
wire x_32684;
wire x_32685;
wire x_32686;
wire x_32687;
wire x_32688;
wire x_32689;
wire x_32690;
wire x_32691;
wire x_32692;
wire x_32693;
wire x_32694;
wire x_32695;
wire x_32696;
wire x_32697;
wire x_32698;
wire x_32699;
wire x_32700;
wire x_32701;
wire x_32702;
wire x_32703;
wire x_32704;
wire x_32705;
wire x_32706;
wire x_32707;
wire x_32708;
wire x_32709;
wire x_32710;
wire x_32711;
wire x_32712;
wire x_32713;
wire x_32714;
wire x_32715;
wire x_32716;
wire x_32717;
wire x_32718;
wire x_32719;
wire x_32720;
wire x_32721;
wire x_32722;
wire x_32723;
wire x_32724;
wire x_32725;
wire x_32726;
wire x_32727;
wire x_32728;
wire x_32729;
wire x_32730;
wire x_32731;
wire x_32732;
wire x_32733;
wire x_32734;
wire x_32735;
wire x_32736;
wire x_32737;
wire x_32738;
wire x_32739;
wire x_32740;
wire x_32741;
wire x_32742;
wire x_32743;
wire x_32744;
wire x_32745;
wire x_32746;
wire x_32747;
wire x_32748;
wire x_32749;
wire x_32750;
wire x_32751;
wire x_32752;
wire x_32753;
wire x_32754;
wire x_32755;
wire x_32756;
wire x_32757;
wire x_32758;
wire x_32759;
wire x_32760;
wire x_32761;
wire x_32762;
wire x_32763;
wire x_32764;
wire x_32765;
wire x_32766;
wire x_32767;
wire x_32768;
wire x_32769;
wire x_32770;
wire x_32771;
wire x_32772;
wire x_32773;
wire x_32774;
wire x_32775;
wire x_32776;
wire x_32777;
wire x_32778;
wire x_32779;
wire x_32780;
wire x_32781;
wire x_32782;
wire x_32783;
wire x_32784;
wire x_32785;
wire x_32786;
wire x_32787;
wire x_32788;
wire x_32789;
wire x_32790;
wire x_32791;
wire x_32792;
wire x_32793;
wire x_32794;
wire x_32795;
wire x_32796;
wire x_32797;
wire x_32798;
wire x_32799;
wire x_32800;
wire x_32801;
wire x_32802;
wire x_32803;
wire x_32804;
wire x_32805;
wire x_32806;
wire x_32807;
wire x_32808;
wire x_32809;
wire x_32810;
wire x_32811;
wire x_32812;
wire x_32813;
wire x_32814;
wire x_32815;
wire x_32816;
wire x_32817;
wire x_32818;
wire x_32819;
wire x_32820;
wire x_32821;
wire x_32822;
wire x_32823;
wire x_32824;
wire x_32825;
wire x_32826;
wire x_32827;
wire x_32828;
wire x_32829;
wire x_32830;
wire x_32831;
wire x_32832;
wire x_32833;
wire x_32834;
wire x_32835;
wire x_32836;
wire x_32837;
wire x_32838;
wire x_32839;
wire x_32840;
wire x_32841;
wire x_32842;
wire x_32843;
wire x_32844;
wire x_32845;
wire x_32846;
wire x_32847;
wire x_32848;
wire x_32849;
wire x_32850;
wire x_32851;
wire x_32852;
wire x_32853;
wire x_32854;
wire x_32855;
wire x_32856;
wire x_32857;
wire x_32858;
wire x_32859;
wire x_32860;
wire x_32861;
wire x_32862;
wire x_32863;
wire x_32864;
wire x_32865;
wire x_32866;
wire x_32867;
wire x_32868;
wire x_32869;
wire x_32870;
wire x_32871;
wire x_32872;
wire x_32873;
wire x_32874;
wire x_32875;
wire x_32876;
wire x_32877;
wire x_32878;
wire x_32879;
wire x_32880;
wire x_32881;
wire x_32882;
wire x_32883;
wire x_32884;
wire x_32885;
wire x_32886;
wire x_32887;
wire x_32888;
wire x_32889;
wire x_32890;
wire x_32891;
wire x_32892;
wire x_32893;
wire x_32894;
wire x_32895;
wire x_32896;
wire x_32897;
wire x_32898;
wire x_32899;
wire x_32900;
wire x_32901;
wire x_32902;
wire x_32903;
wire x_32904;
wire x_32905;
wire x_32906;
wire x_32907;
wire x_32908;
wire x_32909;
wire x_32910;
wire x_32911;
wire x_32912;
wire x_32913;
wire x_32914;
wire x_32915;
wire x_32916;
wire x_32917;
wire x_32918;
wire x_32919;
wire x_32920;
wire x_32921;
wire x_32922;
wire x_32923;
wire x_32924;
wire x_32925;
wire x_32926;
wire x_32927;
wire x_32928;
wire x_32929;
wire x_32930;
wire x_32931;
wire x_32932;
wire x_32933;
wire x_32934;
wire x_32935;
wire x_32936;
wire x_32937;
wire x_32938;
wire x_32939;
wire x_32940;
wire x_32941;
wire x_32942;
wire x_32943;
wire x_32944;
wire x_32945;
wire x_32946;
wire x_32947;
wire x_32948;
wire x_32949;
wire x_32950;
wire x_32951;
wire x_32952;
wire x_32953;
wire x_32954;
wire x_32955;
wire x_32956;
wire x_32957;
wire x_32958;
wire x_32959;
wire x_32960;
wire x_32961;
wire x_32962;
wire x_32963;
wire x_32964;
wire x_32965;
wire x_32966;
wire x_32967;
wire x_32968;
wire x_32969;
wire x_32970;
wire x_32971;
wire x_32972;
wire x_32973;
wire x_32974;
wire x_32975;
wire x_32976;
wire x_32977;
wire x_32978;
wire x_32979;
wire x_32980;
wire x_32981;
wire x_32982;
wire x_32983;
wire x_32984;
wire x_32985;
wire x_32986;
wire x_32987;
wire x_32988;
wire x_32989;
wire x_32990;
wire x_32991;
wire x_32992;
wire x_32993;
wire x_32994;
wire x_32995;
wire x_32996;
wire x_32997;
wire x_32998;
wire x_32999;
wire x_33000;
wire x_33001;
wire x_33002;
wire x_33003;
wire x_33004;
wire x_33005;
wire x_33006;
wire x_33007;
wire x_33008;
wire x_33009;
wire x_33010;
wire x_33011;
wire x_33012;
wire x_33013;
wire x_33014;
wire x_33015;
wire x_33016;
wire x_33017;
wire x_33018;
wire x_33019;
wire x_33020;
wire x_33021;
wire x_33022;
wire x_33023;
wire x_33024;
wire x_33025;
wire x_33026;
wire x_33027;
wire x_33028;
wire x_33029;
wire x_33030;
wire x_33031;
wire x_33032;
wire x_33033;
wire x_33034;
wire x_33035;
wire x_33036;
wire x_33037;
wire x_33038;
wire x_33039;
wire x_33040;
wire x_33041;
wire x_33042;
wire x_33043;
wire x_33044;
wire x_33045;
wire x_33046;
wire x_33047;
wire x_33048;
wire x_33049;
wire x_33050;
wire x_33051;
wire x_33052;
wire x_33053;
wire x_33054;
wire x_33055;
wire x_33056;
wire x_33057;
wire x_33058;
wire x_33059;
wire x_33060;
wire x_33061;
wire x_33062;
wire x_33063;
wire x_33064;
wire x_33065;
wire x_33066;
wire x_33067;
wire x_33068;
wire x_33069;
wire x_33070;
wire x_33071;
wire x_33072;
wire x_33073;
wire x_33074;
wire x_33075;
wire x_33076;
wire x_33077;
wire x_33078;
wire x_33079;
wire x_33080;
wire x_33081;
wire x_33082;
wire x_33083;
wire x_33084;
wire x_33085;
wire x_33086;
wire x_33087;
wire x_33088;
wire x_33089;
wire x_33090;
wire x_33091;
wire x_33092;
wire x_33093;
wire x_33094;
wire x_33095;
wire x_33096;
wire x_33097;
wire x_33098;
wire x_33099;
wire x_33100;
wire x_33101;
wire x_33102;
wire x_33103;
wire x_33104;
wire x_33105;
wire x_33106;
wire x_33107;
wire x_33108;
wire x_33109;
wire x_33110;
wire x_33111;
wire x_33112;
wire x_33113;
wire x_33114;
wire x_33115;
wire x_33116;
wire x_33117;
wire x_33118;
wire x_33119;
wire x_33120;
wire x_33121;
wire x_33122;
wire x_33123;
wire x_33124;
wire x_33125;
wire x_33126;
wire x_33127;
wire x_33128;
wire x_33129;
wire x_33130;
wire x_33131;
wire x_33132;
wire x_33133;
wire x_33134;
wire x_33135;
wire x_33136;
wire x_33137;
wire x_33138;
wire x_33139;
wire x_33140;
wire x_33141;
wire x_33142;
wire x_33143;
wire x_33144;
wire x_33145;
wire x_33146;
wire x_33147;
wire x_33148;
wire x_33149;
wire x_33150;
wire x_33151;
wire x_33152;
wire x_33153;
wire x_33154;
wire x_33155;
wire x_33156;
wire x_33157;
wire x_33158;
wire x_33159;
wire x_33160;
wire x_33161;
wire x_33162;
wire x_33163;
wire x_33164;
wire x_33165;
wire x_33166;
wire x_33167;
wire x_33168;
wire x_33169;
wire x_33170;
wire x_33171;
wire x_33172;
wire x_33173;
wire x_33174;
wire x_33175;
wire x_33176;
wire x_33177;
wire x_33178;
wire x_33179;
wire x_33180;
wire x_33181;
wire x_33182;
wire x_33183;
wire x_33184;
wire x_33185;
wire x_33186;
wire x_33187;
wire x_33188;
wire x_33189;
wire x_33190;
wire x_33191;
wire x_33192;
wire x_33193;
wire x_33194;
wire x_33195;
wire x_33196;
wire x_33197;
wire x_33198;
wire x_33199;
wire x_33200;
wire x_33201;
wire x_33202;
wire x_33203;
wire x_33204;
wire x_33205;
wire x_33206;
wire x_33207;
wire x_33208;
wire x_33209;
wire x_33210;
wire x_33211;
wire x_33212;
wire x_33213;
wire x_33214;
wire x_33215;
wire x_33216;
wire x_33217;
wire x_33218;
wire x_33219;
wire x_33220;
wire x_33221;
wire x_33222;
wire x_33223;
wire x_33224;
wire x_33225;
wire x_33226;
wire x_33227;
wire x_33228;
wire x_33229;
wire x_33230;
wire x_33231;
wire x_33232;
wire x_33233;
wire x_33234;
wire x_33235;
wire x_33236;
wire x_33237;
wire x_33238;
wire x_33239;
wire x_33240;
wire x_33241;
wire x_33242;
wire x_33243;
wire x_33244;
wire x_33245;
wire x_33246;
wire x_33247;
wire x_33248;
wire x_33249;
wire x_33250;
wire x_33251;
wire x_33252;
wire x_33253;
wire x_33254;
wire x_33255;
wire x_33256;
wire x_33257;
wire x_33258;
wire x_33259;
wire x_33260;
wire x_33261;
wire x_33262;
wire x_33263;
wire x_33264;
wire x_33265;
wire x_33266;
wire x_33267;
wire x_33268;
wire x_33269;
wire x_33270;
wire x_33271;
wire x_33272;
wire x_33273;
wire x_33274;
wire x_33275;
wire x_33276;
wire x_33277;
wire x_33278;
wire x_33279;
wire x_33280;
wire x_33281;
wire x_33282;
wire x_33283;
wire x_33284;
wire x_33285;
wire x_33286;
wire x_33287;
wire x_33288;
wire x_33289;
wire x_33290;
wire x_33291;
wire x_33292;
wire x_33293;
wire x_33294;
wire x_33295;
wire x_33296;
wire x_33297;
wire x_33298;
wire x_33299;
wire x_33300;
wire x_33301;
wire x_33302;
wire x_33303;
wire x_33304;
wire x_33305;
wire x_33306;
wire x_33307;
wire x_33308;
wire x_33309;
wire x_33310;
wire x_33311;
wire x_33312;
wire x_33313;
wire x_33314;
wire x_33315;
wire x_33316;
wire x_33317;
wire x_33318;
wire x_33319;
wire x_33320;
wire x_33321;
wire x_33322;
wire x_33323;
wire x_33324;
wire x_33325;
wire x_33326;
wire x_33327;
wire x_33328;
wire x_33329;
wire x_33330;
wire x_33331;
wire x_33332;
wire x_33333;
wire x_33334;
wire x_33335;
wire x_33336;
wire x_33337;
wire x_33338;
wire x_33339;
wire x_33340;
wire x_33341;
wire x_33342;
wire x_33343;
wire x_33344;
wire x_33345;
wire x_33346;
wire x_33347;
wire x_33348;
wire x_33349;
wire x_33350;
wire x_33351;
wire x_33352;
wire x_33353;
wire x_33354;
wire x_33355;
wire x_33356;
wire x_33357;
wire x_33358;
wire x_33359;
wire x_33360;
wire x_33361;
wire x_33362;
wire x_33363;
wire x_33364;
wire x_33365;
wire x_33366;
wire x_33367;
wire x_33368;
wire x_33369;
wire x_33370;
wire x_33371;
wire x_33372;
wire x_33373;
wire x_33374;
wire x_33375;
wire x_33376;
wire x_33377;
wire x_33378;
wire x_33379;
wire x_33380;
wire x_33381;
wire x_33382;
wire x_33383;
wire x_33384;
wire x_33385;
wire x_33386;
wire x_33387;
wire x_33388;
wire x_33389;
wire x_33390;
wire x_33391;
wire x_33392;
wire x_33393;
wire x_33394;
wire x_33395;
wire x_33396;
wire x_33397;
wire x_33398;
wire x_33399;
wire x_33400;
wire x_33401;
wire x_33402;
wire x_33403;
wire x_33404;
wire x_33405;
wire x_33406;
wire x_33407;
wire x_33408;
wire x_33409;
wire x_33410;
wire x_33411;
wire x_33412;
wire x_33413;
wire x_33414;
wire x_33415;
wire x_33416;
wire x_33417;
wire x_33418;
wire x_33419;
wire x_33420;
wire x_33421;
wire x_33422;
wire x_33423;
wire x_33424;
wire x_33425;
wire x_33426;
wire x_33427;
wire x_33428;
wire x_33429;
wire x_33430;
wire x_33431;
wire x_33432;
wire x_33433;
wire x_33434;
wire x_33435;
wire x_33436;
wire x_33437;
wire x_33438;
wire x_33439;
wire x_33440;
wire x_33441;
wire x_33442;
wire x_33443;
wire x_33444;
wire x_33445;
wire x_33446;
wire x_33447;
wire x_33448;
wire x_33449;
wire x_33450;
wire x_33451;
wire x_33452;
wire x_33453;
wire x_33454;
wire x_33455;
wire x_33456;
wire x_33457;
wire x_33458;
wire x_33459;
wire x_33460;
wire x_33461;
wire x_33462;
wire x_33463;
wire x_33464;
wire x_33465;
wire x_33466;
wire x_33467;
wire x_33468;
wire x_33469;
wire x_33470;
wire x_33471;
wire x_33472;
wire x_33473;
wire x_33474;
wire x_33475;
wire x_33476;
wire x_33477;
wire x_33478;
wire x_33479;
wire x_33480;
wire x_33481;
wire x_33482;
wire x_33483;
wire x_33484;
wire x_33485;
wire x_33486;
wire x_33487;
wire x_33488;
wire x_33489;
wire x_33490;
wire x_33491;
wire x_33492;
wire x_33493;
wire x_33494;
wire x_33495;
wire x_33496;
wire x_33497;
wire x_33498;
wire x_33499;
wire x_33500;
wire x_33501;
wire x_33502;
wire x_33503;
wire x_33504;
wire x_33505;
wire x_33506;
wire x_33507;
wire x_33508;
wire x_33509;
wire x_33510;
wire x_33511;
wire x_33512;
wire x_33513;
wire x_33514;
wire x_33515;
wire x_33516;
wire x_33517;
wire x_33518;
wire x_33519;
wire x_33520;
wire x_33521;
wire x_33522;
wire x_33523;
wire x_33524;
wire x_33525;
wire x_33526;
wire x_33527;
wire x_33528;
wire x_33529;
wire x_33530;
wire x_33531;
wire x_33532;
wire x_33533;
wire x_33534;
wire x_33535;
wire x_33536;
wire x_33537;
wire x_33538;
wire x_33539;
wire x_33540;
wire x_33541;
wire x_33542;
wire x_33543;
wire x_33544;
wire x_33545;
wire x_33546;
wire x_33547;
wire x_33548;
wire x_33549;
wire x_33550;
wire x_33551;
wire x_33552;
wire x_33553;
wire x_33554;
wire x_33555;
wire x_33556;
wire x_33557;
wire x_33558;
wire x_33559;
wire x_33560;
wire x_33561;
wire x_33562;
wire x_33563;
wire x_33564;
wire x_33565;
wire x_33566;
wire x_33567;
wire x_33568;
wire x_33569;
wire x_33570;
wire x_33571;
wire x_33572;
wire x_33573;
wire x_33574;
wire x_33575;
wire x_33576;
wire x_33577;
wire x_33578;
wire x_33579;
wire x_33580;
wire x_33581;
wire x_33582;
wire x_33583;
wire x_33584;
wire x_33585;
wire x_33586;
wire x_33587;
wire x_33588;
wire x_33589;
wire x_33590;
wire x_33591;
wire x_33592;
wire x_33593;
wire x_33594;
wire x_33595;
wire x_33596;
wire x_33597;
wire x_33598;
wire x_33599;
wire x_33600;
wire x_33601;
wire x_33602;
wire x_33603;
wire x_33604;
wire x_33605;
wire x_33606;
wire x_33607;
wire x_33608;
wire x_33609;
wire x_33610;
wire x_33611;
wire x_33612;
wire x_33613;
wire x_33614;
wire x_33615;
wire x_33616;
wire x_33617;
wire x_33618;
wire x_33619;
wire x_33620;
wire x_33621;
wire x_33622;
wire x_33623;
wire x_33624;
wire x_33625;
wire x_33626;
wire x_33627;
wire x_33628;
wire x_33629;
wire x_33630;
wire x_33631;
wire x_33632;
wire x_33633;
wire x_33634;
wire x_33635;
wire x_33636;
wire x_33637;
wire x_33638;
wire x_33639;
wire x_33640;
wire x_33641;
wire x_33642;
wire x_33643;
wire x_33644;
wire x_33645;
wire x_33646;
wire x_33647;
wire x_33648;
wire x_33649;
wire x_33650;
wire x_33651;
wire x_33652;
wire x_33653;
wire x_33654;
wire x_33655;
wire x_33656;
wire x_33657;
wire x_33658;
wire x_33659;
wire x_33660;
wire x_33661;
wire x_33662;
wire x_33663;
wire x_33664;
wire x_33665;
wire x_33666;
wire x_33667;
wire x_33668;
wire x_33669;
wire x_33670;
wire x_33671;
wire x_33672;
wire x_33673;
wire x_33674;
wire x_33675;
wire x_33676;
wire x_33677;
wire x_33678;
wire x_33679;
wire x_33680;
wire x_33681;
wire x_33682;
wire x_33683;
wire x_33684;
wire x_33685;
wire x_33686;
wire x_33687;
wire x_33688;
wire x_33689;
wire x_33690;
wire x_33691;
wire x_33692;
wire x_33693;
wire x_33694;
wire x_33695;
wire x_33696;
wire x_33697;
wire x_33698;
wire x_33699;
wire x_33700;
wire x_33701;
wire x_33702;
wire x_33703;
wire x_33704;
wire x_33705;
wire x_33706;
wire x_33707;
wire x_33708;
wire x_33709;
wire x_33710;
wire x_33711;
wire x_33712;
wire x_33713;
wire x_33714;
wire x_33715;
wire x_33716;
wire x_33717;
wire x_33718;
wire x_33719;
wire x_33720;
wire x_33721;
wire x_33722;
wire x_33723;
wire x_33724;
wire x_33725;
wire x_33726;
wire x_33727;
wire x_33728;
wire x_33729;
wire x_33730;
wire x_33731;
wire x_33732;
wire x_33733;
wire x_33734;
wire x_33735;
wire x_33736;
wire x_33737;
wire x_33738;
wire x_33739;
wire x_33740;
wire x_33741;
wire x_33742;
wire x_33743;
wire x_33744;
wire x_33745;
wire x_33746;
wire x_33747;
wire x_33748;
wire x_33749;
wire x_33750;
wire x_33751;
wire x_33752;
wire x_33753;
wire x_33754;
wire x_33755;
wire x_33756;
wire x_33757;
wire x_33758;
wire x_33759;
wire x_33760;
wire x_33761;
wire x_33762;
wire x_33763;
wire x_33764;
wire x_33765;
wire x_33766;
wire x_33767;
wire x_33768;
wire x_33769;
wire x_33770;
wire x_33771;
wire x_33772;
wire x_33773;
wire x_33774;
wire x_33775;
wire x_33776;
wire x_33777;
wire x_33778;
wire x_33779;
wire x_33780;
wire x_33781;
wire x_33782;
wire x_33783;
wire x_33784;
wire x_33785;
wire x_33786;
wire x_33787;
wire x_33788;
wire x_33789;
wire x_33790;
wire x_33791;
wire x_33792;
wire x_33793;
wire x_33794;
wire x_33795;
wire x_33796;
wire x_33797;
wire x_33798;
wire x_33799;
wire x_33800;
wire x_33801;
wire x_33802;
wire x_33803;
wire x_33804;
wire x_33805;
wire x_33806;
wire x_33807;
wire x_33808;
wire x_33809;
wire x_33810;
wire x_33811;
wire x_33812;
wire x_33813;
wire x_33814;
wire x_33815;
wire x_33816;
wire x_33817;
wire x_33818;
wire x_33819;
wire x_33820;
wire x_33821;
wire x_33822;
wire x_33823;
wire x_33824;
wire x_33825;
wire x_33826;
wire x_33827;
wire x_33828;
wire x_33829;
wire x_33830;
wire x_33831;
wire x_33832;
wire x_33833;
wire x_33834;
wire x_33835;
wire x_33836;
wire x_33837;
wire x_33838;
wire x_33839;
wire x_33840;
wire x_33841;
wire x_33842;
wire x_33843;
wire x_33844;
wire x_33845;
wire x_33846;
wire x_33847;
wire x_33848;
wire x_33849;
wire x_33850;
wire x_33851;
wire x_33852;
wire x_33853;
wire x_33854;
wire x_33855;
wire x_33856;
wire x_33857;
wire x_33858;
wire x_33859;
wire x_33860;
wire x_33861;
wire x_33862;
wire x_33863;
wire x_33864;
wire x_33865;
wire x_33866;
wire x_33867;
wire x_33868;
wire x_33869;
wire x_33870;
wire x_33871;
wire x_33872;
wire x_33873;
wire x_33874;
wire x_33875;
wire x_33876;
wire x_33877;
wire x_33878;
wire x_33879;
wire x_33880;
wire x_33881;
wire x_33882;
wire x_33883;
wire x_33884;
wire x_33885;
wire x_33886;
wire x_33887;
wire x_33888;
wire x_33889;
wire x_33890;
wire x_33891;
wire x_33892;
wire x_33893;
wire x_33894;
wire x_33895;
wire x_33896;
wire x_33897;
wire x_33898;
wire x_33899;
wire x_33900;
wire x_33901;
wire x_33902;
wire x_33903;
wire x_33904;
wire x_33905;
wire x_33906;
wire x_33907;
wire x_33908;
wire x_33909;
wire x_33910;
wire x_33911;
wire x_33912;
wire x_33913;
wire x_33914;
wire x_33915;
wire x_33916;
wire x_33917;
wire x_33918;
wire x_33919;
wire x_33920;
wire x_33921;
wire x_33922;
wire x_33923;
wire x_33924;
wire x_33925;
wire x_33926;
wire x_33927;
wire x_33928;
wire x_33929;
wire x_33930;
wire x_33931;
wire x_33932;
wire x_33933;
wire x_33934;
wire x_33935;
wire x_33936;
wire x_33937;
wire x_33938;
wire x_33939;
wire x_33940;
wire x_33941;
wire x_33942;
wire x_33943;
wire x_33944;
wire x_33945;
wire x_33946;
wire x_33947;
wire x_33948;
wire x_33949;
wire x_33950;
wire x_33951;
wire x_33952;
wire x_33953;
wire x_33954;
wire x_33955;
wire x_33956;
wire x_33957;
wire x_33958;
wire x_33959;
wire x_33960;
wire x_33961;
wire x_33962;
wire x_33963;
wire x_33964;
wire x_33965;
wire x_33966;
wire x_33967;
wire x_33968;
wire x_33969;
wire x_33970;
wire x_33971;
wire x_33972;
wire x_33973;
wire x_33974;
wire x_33975;
wire x_33976;
wire x_33977;
wire x_33978;
wire x_33979;
wire x_33980;
wire x_33981;
wire x_33982;
wire x_33983;
wire x_33984;
wire x_33985;
wire x_33986;
wire x_33987;
wire x_33988;
wire x_33989;
wire x_33990;
wire x_33991;
wire x_33992;
wire x_33993;
wire x_33994;
wire x_33995;
wire x_33996;
wire x_33997;
wire x_33998;
wire x_33999;
wire x_34000;
wire x_34001;
wire x_34002;
wire x_34003;
wire x_34004;
wire x_34005;
wire x_34006;
wire x_34007;
wire x_34008;
wire x_34009;
wire x_34010;
wire x_34011;
wire x_34012;
wire x_34013;
wire x_34014;
wire x_34015;
wire x_34016;
wire x_34017;
wire x_34018;
wire x_34019;
wire x_34020;
wire x_34021;
wire x_34022;
wire x_34023;
wire x_34024;
wire x_34025;
wire x_34026;
wire x_34027;
wire x_34028;
wire x_34029;
wire x_34030;
wire x_34031;
wire x_34032;
wire x_34033;
wire x_34034;
wire x_34035;
wire x_34036;
wire x_34037;
wire x_34038;
wire x_34039;
wire x_34040;
wire x_34041;
wire x_34042;
wire x_34043;
wire x_34044;
wire x_34045;
wire x_34046;
wire x_34047;
wire x_34048;
wire x_34049;
wire x_34050;
wire x_34051;
wire x_34052;
wire x_34053;
wire x_34054;
wire x_34055;
wire x_34056;
wire x_34057;
wire x_34058;
wire x_34059;
wire x_34060;
wire x_34061;
wire x_34062;
wire x_34063;
wire x_34064;
wire x_34065;
wire x_34066;
wire x_34067;
wire x_34068;
wire x_34069;
wire x_34070;
wire x_34071;
wire x_34072;
wire x_34073;
wire x_34074;
wire x_34075;
wire x_34076;
wire x_34077;
wire x_34078;
wire x_34079;
wire x_34080;
wire x_34081;
wire x_34082;
wire x_34083;
wire x_34084;
wire x_34085;
wire x_34086;
wire x_34087;
wire x_34088;
wire x_34089;
wire x_34090;
wire x_34091;
wire x_34092;
wire x_34093;
wire x_34094;
wire x_34095;
wire x_34096;
wire x_34097;
wire x_34098;
wire x_34099;
wire x_34100;
wire x_34101;
wire x_34102;
wire x_34103;
wire x_34104;
wire x_34105;
wire x_34106;
wire x_34107;
wire x_34108;
wire x_34109;
wire x_34110;
wire x_34111;
wire x_34112;
wire x_34113;
wire x_34114;
wire x_34115;
wire x_34116;
wire x_34117;
wire x_34118;
wire x_34119;
wire x_34120;
wire x_34121;
wire x_34122;
wire x_34123;
wire x_34124;
wire x_34125;
wire x_34126;
wire x_34127;
wire x_34128;
wire x_34129;
wire x_34130;
wire x_34131;
wire x_34132;
wire x_34133;
wire x_34134;
wire x_34135;
wire x_34136;
wire x_34137;
wire x_34138;
wire x_34139;
wire x_34140;
wire x_34141;
wire x_34142;
wire x_34143;
wire x_34144;
wire x_34145;
wire x_34146;
wire x_34147;
wire x_34148;
wire x_34149;
wire x_34150;
wire x_34151;
wire x_34152;
wire x_34153;
wire x_34154;
wire x_34155;
wire x_34156;
wire x_34157;
wire x_34158;
wire x_34159;
wire x_34160;
wire x_34161;
wire x_34162;
wire x_34163;
wire x_34164;
wire x_34165;
wire x_34166;
wire x_34167;
wire x_34168;
wire x_34169;
wire x_34170;
wire x_34171;
wire x_34172;
wire x_34173;
wire x_34174;
wire x_34175;
wire x_34176;
wire x_34177;
wire x_34178;
wire x_34179;
wire x_34180;
wire x_34181;
wire x_34182;
wire x_34183;
wire x_34184;
wire x_34185;
wire x_34186;
wire x_34187;
wire x_34188;
wire x_34189;
wire x_34190;
wire x_34191;
wire x_34192;
wire x_34193;
wire x_34194;
wire x_34195;
wire x_34196;
wire x_34197;
wire x_34198;
wire x_34199;
wire x_34200;
wire x_34201;
wire x_34202;
wire x_34203;
wire x_34204;
wire x_34205;
wire x_34206;
wire x_34207;
wire x_34208;
wire x_34209;
wire x_34210;
wire x_34211;
wire x_34212;
wire x_34213;
wire x_34214;
wire x_34215;
wire x_34216;
wire x_34217;
wire x_34218;
wire x_34219;
wire x_34220;
wire x_34221;
wire x_34222;
wire x_34223;
wire x_34224;
wire x_34225;
wire x_34226;
wire x_34227;
wire x_34228;
wire x_34229;
wire x_34230;
wire x_34231;
wire x_34232;
wire x_34233;
wire x_34234;
wire x_34235;
wire x_34236;
wire x_34237;
wire x_34238;
wire x_34239;
wire x_34240;
wire x_34241;
wire x_34242;
wire x_34243;
wire x_34244;
wire x_34245;
wire x_34246;
wire x_34247;
wire x_34248;
wire x_34249;
wire x_34250;
wire x_34251;
wire x_34252;
wire x_34253;
wire x_34254;
wire x_34255;
wire x_34256;
wire x_34257;
wire x_34258;
wire x_34259;
wire x_34260;
wire x_34261;
wire x_34262;
wire x_34263;
wire x_34264;
wire x_34265;
wire x_34266;
wire x_34267;
wire x_34268;
wire x_34269;
wire x_34270;
wire x_34271;
wire x_34272;
wire x_34273;
wire x_34274;
wire x_34275;
wire x_34276;
wire x_34277;
wire x_34278;
wire x_34279;
wire x_34280;
wire x_34281;
wire x_34282;
wire x_34283;
wire x_34284;
wire x_34285;
wire x_34286;
wire x_34287;
wire x_34288;
wire x_34289;
wire x_34290;
wire x_34291;
wire x_34292;
wire x_34293;
wire x_34294;
wire x_34295;
wire x_34296;
wire x_34297;
wire x_34298;
wire x_34299;
wire x_34300;
wire x_34301;
wire x_34302;
wire x_34303;
wire x_34304;
wire x_34305;
wire x_34306;
wire x_34307;
wire x_34308;
wire x_34309;
wire x_34310;
wire x_34311;
wire x_34312;
wire x_34313;
wire x_34314;
wire x_34315;
wire x_34316;
wire x_34317;
wire x_34318;
wire x_34319;
wire x_34320;
wire x_34321;
wire x_34322;
wire x_34323;
wire x_34324;
wire x_34325;
wire x_34326;
wire x_34327;
wire x_34328;
wire x_34329;
wire x_34330;
wire x_34331;
wire x_34332;
wire x_34333;
wire x_34334;
wire x_34335;
wire x_34336;
wire x_34337;
wire x_34338;
wire x_34339;
wire x_34340;
wire x_34341;
wire x_34342;
wire x_34343;
wire x_34344;
wire x_34345;
wire x_34346;
wire x_34347;
wire x_34348;
wire x_34349;
wire x_34350;
wire x_34351;
wire x_34352;
wire x_34353;
wire x_34354;
wire x_34355;
wire x_34356;
wire x_34357;
wire x_34358;
wire x_34359;
wire x_34360;
wire x_34361;
wire x_34362;
wire x_34363;
wire x_34364;
wire x_34365;
wire x_34366;
wire x_34367;
wire x_34368;
wire x_34369;
wire x_34370;
wire x_34371;
wire x_34372;
wire x_34373;
wire x_34374;
wire x_34375;
wire x_34376;
wire x_34377;
wire x_34378;
wire x_34379;
wire x_34380;
wire x_34381;
wire x_34382;
wire x_34383;
wire x_34384;
wire x_34385;
wire x_34386;
wire x_34387;
wire x_34388;
wire x_34389;
wire x_34390;
wire x_34391;
wire x_34392;
wire x_34393;
wire x_34394;
wire x_34395;
wire x_34396;
wire x_34397;
wire x_34398;
wire x_34399;
wire x_34400;
wire x_34401;
wire x_34402;
wire x_34403;
wire x_34404;
wire x_34405;
wire x_34406;
wire x_34407;
wire x_34408;
wire x_34409;
wire x_34410;
wire x_34411;
wire x_34412;
wire x_34413;
wire x_34414;
wire x_34415;
wire x_34416;
wire x_34417;
wire x_34418;
wire x_34419;
wire x_34420;
wire x_34421;
wire x_34422;
wire x_34423;
wire x_34424;
wire x_34425;
wire x_34426;
wire x_34427;
wire x_34428;
wire x_34429;
wire x_34430;
wire x_34431;
wire x_34432;
wire x_34433;
wire x_34434;
wire x_34435;
wire x_34436;
wire x_34437;
wire x_34438;
wire x_34439;
wire x_34440;
wire x_34441;
wire x_34442;
wire x_34443;
wire x_34444;
wire x_34445;
wire x_34446;
wire x_34447;
wire x_34448;
wire x_34449;
wire x_34450;
wire x_34451;
wire x_34452;
wire x_34453;
wire x_34454;
wire x_34455;
wire x_34456;
wire x_34457;
wire x_34458;
wire x_34459;
wire x_34460;
wire x_34461;
wire x_34462;
wire x_34463;
wire x_34464;
wire x_34465;
wire x_34466;
wire x_34467;
wire x_34468;
wire x_34469;
wire x_34470;
wire x_34471;
wire x_34472;
wire x_34473;
wire x_34474;
wire x_34475;
wire x_34476;
wire x_34477;
wire x_34478;
wire x_34479;
wire x_34480;
wire x_34481;
wire x_34482;
wire x_34483;
wire x_34484;
wire x_34485;
wire x_34486;
wire x_34487;
wire x_34488;
wire x_34489;
wire x_34490;
wire x_34491;
wire x_34492;
wire x_34493;
wire x_34494;
wire x_34495;
wire x_34496;
wire x_34497;
wire x_34498;
wire x_34499;
wire x_34500;
wire x_34501;
wire x_34502;
wire x_34503;
wire x_34504;
wire x_34505;
wire x_34506;
wire x_34507;
wire x_34508;
wire x_34509;
wire x_34510;
wire x_34511;
wire x_34512;
wire x_34513;
wire x_34514;
wire x_34515;
wire x_34516;
wire x_34517;
wire x_34518;
wire x_34519;
wire x_34520;
wire x_34521;
wire x_34522;
wire x_34523;
wire x_34524;
wire x_34525;
wire x_34526;
wire x_34527;
wire x_34528;
wire x_34529;
wire x_34530;
wire x_34531;
wire x_34532;
wire x_34533;
wire x_34534;
wire x_34535;
wire x_34536;
wire x_34537;
wire x_34538;
wire x_34539;
wire x_34540;
wire x_34541;
wire x_34542;
wire x_34543;
wire x_34544;
wire x_34545;
wire x_34546;
wire x_34547;
wire x_34548;
wire x_34549;
wire x_34550;
wire x_34551;
wire x_34552;
wire x_34553;
wire x_34554;
wire x_34555;
wire x_34556;
wire x_34557;
wire x_34558;
wire x_34559;
wire x_34560;
wire x_34561;
wire x_34562;
wire x_34563;
wire x_34564;
wire x_34565;
wire x_34566;
wire x_34567;
wire x_34568;
wire x_34569;
wire x_34570;
wire x_34571;
wire x_34572;
wire x_34573;
wire x_34574;
wire x_34575;
wire x_34576;
wire x_34577;
wire x_34578;
wire x_34579;
wire x_34580;
wire x_34581;
wire x_34582;
wire x_34583;
wire x_34584;
wire x_34585;
wire x_34586;
wire x_34587;
wire x_34588;
wire x_34589;
wire x_34590;
wire x_34591;
wire x_34592;
wire x_34593;
wire x_34594;
wire x_34595;
wire x_34596;
wire x_34597;
wire x_34598;
wire x_34599;
wire x_34600;
wire x_34601;
wire x_34602;
wire x_34603;
wire x_34604;
wire x_34605;
wire x_34606;
wire x_34607;
wire x_34608;
wire x_34609;
wire x_34610;
wire x_34611;
wire x_34612;
wire x_34613;
wire x_34614;
wire x_34615;
wire x_34616;
wire x_34617;
wire x_34618;
wire x_34619;
wire x_34620;
wire x_34621;
wire x_34622;
wire x_34623;
wire x_34624;
wire x_34625;
wire x_34626;
wire x_34627;
wire x_34628;
wire x_34629;
wire x_34630;
wire x_34631;
wire x_34632;
wire x_34633;
wire x_34634;
wire x_34635;
wire x_34636;
wire x_34637;
wire x_34638;
wire x_34639;
wire x_34640;
wire x_34641;
wire x_34642;
wire x_34643;
wire x_34644;
wire x_34645;
wire x_34646;
wire x_34647;
wire x_34648;
wire x_34649;
wire x_34650;
wire x_34651;
wire x_34652;
wire x_34653;
wire x_34654;
wire x_34655;
wire x_34656;
wire x_34657;
wire x_34658;
wire x_34659;
wire x_34660;
wire x_34661;
wire x_34662;
wire x_34663;
wire x_34664;
wire x_34665;
wire x_34666;
wire x_34667;
wire x_34668;
wire x_34669;
wire x_34670;
wire x_34671;
wire x_34672;
wire x_34673;
wire x_34674;
wire x_34675;
wire x_34676;
wire x_34677;
wire x_34678;
wire x_34679;
wire x_34680;
wire x_34681;
wire x_34682;
wire x_34683;
wire x_34684;
wire x_34685;
wire x_34686;
wire x_34687;
wire x_34688;
wire x_34689;
wire x_34690;
wire x_34691;
wire x_34692;
wire x_34693;
wire x_34694;
wire x_34695;
wire x_34696;
wire x_34697;
wire x_34698;
wire x_34699;
wire x_34700;
wire x_34701;
wire x_34702;
wire x_34703;
wire x_34704;
wire x_34705;
wire x_34706;
wire x_34707;
wire x_34708;
wire x_34709;
wire x_34710;
wire x_34711;
wire x_34712;
wire x_34713;
wire x_34714;
wire x_34715;
wire x_34716;
wire x_34717;
wire x_34718;
wire x_34719;
wire x_34720;
wire x_34721;
wire x_34722;
wire x_34723;
wire x_34724;
wire x_34725;
wire x_34726;
wire x_34727;
wire x_34728;
wire x_34729;
wire x_34730;
wire x_34731;
wire x_34732;
wire x_34733;
wire x_34734;
wire x_34735;
wire x_34736;
wire x_34737;
wire x_34738;
wire x_34739;
wire x_34740;
wire x_34741;
wire x_34742;
wire x_34743;
wire x_34744;
wire x_34745;
wire x_34746;
wire x_34747;
wire x_34748;
wire x_34749;
wire x_34750;
wire x_34751;
wire x_34752;
wire x_34753;
wire x_34754;
wire x_34755;
wire x_34756;
wire x_34757;
wire x_34758;
wire x_34759;
wire x_34760;
wire x_34761;
wire x_34762;
wire x_34763;
wire x_34764;
wire x_34765;
wire x_34766;
wire x_34767;
wire x_34768;
wire x_34769;
wire x_34770;
wire x_34771;
wire x_34772;
wire x_34773;
wire x_34774;
wire x_34775;
wire x_34776;
wire x_34777;
wire x_34778;
wire x_34779;
wire x_34780;
wire x_34781;
wire x_34782;
wire x_34783;
wire x_34784;
wire x_34785;
wire x_34786;
wire x_34787;
wire x_34788;
wire x_34789;
wire x_34790;
wire x_34791;
wire x_34792;
wire x_34793;
wire x_34794;
wire x_34795;
wire x_34796;
wire x_34797;
wire x_34798;
wire x_34799;
wire x_34800;
wire x_34801;
wire x_34802;
wire x_34803;
wire x_34804;
wire x_34805;
wire x_34806;
wire x_34807;
wire x_34808;
wire x_34809;
wire x_34810;
wire x_34811;
wire x_34812;
wire x_34813;
wire x_34814;
wire x_34815;
wire x_34816;
wire x_34817;
wire x_34818;
wire x_34819;
wire x_34820;
wire x_34821;
wire x_34822;
wire x_34823;
wire x_34824;
wire x_34825;
wire x_34826;
wire x_34827;
wire x_34828;
wire x_34829;
wire x_34830;
wire x_34831;
wire x_34832;
wire x_34833;
wire x_34834;
wire x_34835;
wire x_34836;
wire x_34837;
wire x_34838;
wire x_34839;
wire x_34840;
wire x_34841;
wire x_34842;
wire x_34843;
wire x_34844;
wire x_34845;
wire x_34846;
wire x_34847;
wire x_34848;
wire x_34849;
wire x_34850;
wire x_34851;
wire x_34852;
wire x_34853;
wire x_34854;
wire x_34855;
wire x_34856;
wire x_34857;
wire x_34858;
wire x_34859;
wire x_34860;
wire x_34861;
wire x_34862;
wire x_34863;
wire x_34864;
wire x_34865;
wire x_34866;
wire x_34867;
wire x_34868;
wire x_34869;
wire x_34870;
wire x_34871;
wire x_34872;
wire x_34873;
wire x_34874;
wire x_34875;
wire x_34876;
wire x_34877;
wire x_34878;
wire x_34879;
wire x_34880;
wire x_34881;
wire x_34882;
wire x_34883;
wire x_34884;
wire x_34885;
wire x_34886;
wire x_34887;
wire x_34888;
wire x_34889;
wire x_34890;
wire x_34891;
wire x_34892;
wire x_34893;
wire x_34894;
wire x_34895;
wire x_34896;
wire x_34897;
wire x_34898;
wire x_34899;
wire x_34900;
wire x_34901;
wire x_34902;
wire x_34903;
wire x_34904;
wire x_34905;
wire x_34906;
wire x_34907;
wire x_34908;
wire x_34909;
wire x_34910;
wire x_34911;
wire x_34912;
wire x_34913;
wire x_34914;
wire x_34915;
wire x_34916;
wire x_34917;
wire x_34918;
wire x_34919;
wire x_34920;
wire x_34921;
wire x_34922;
wire x_34923;
wire x_34924;
wire x_34925;
wire x_34926;
wire x_34927;
wire x_34928;
wire x_34929;
wire x_34930;
wire x_34931;
wire x_34932;
wire x_34933;
wire x_34934;
wire x_34935;
wire x_34936;
wire x_34937;
wire x_34938;
wire x_34939;
wire x_34940;
wire x_34941;
wire x_34942;
wire x_34943;
wire x_34944;
wire x_34945;
wire x_34946;
wire x_34947;
wire x_34948;
wire x_34949;
wire x_34950;
wire x_34951;
wire x_34952;
wire x_34953;
wire x_34954;
wire x_34955;
wire x_34956;
wire x_34957;
wire x_34958;
wire x_34959;
wire x_34960;
wire x_34961;
wire x_34962;
wire x_34963;
wire x_34964;
wire x_34965;
wire x_34966;
wire x_34967;
wire x_34968;
wire x_34969;
wire x_34970;
wire x_34971;
wire x_34972;
wire x_34973;
wire x_34974;
wire x_34975;
wire x_34976;
wire x_34977;
wire x_34978;
wire x_34979;
wire x_34980;
wire x_34981;
wire x_34982;
wire x_34983;
wire x_34984;
wire x_34985;
wire x_34986;
wire x_34987;
wire x_34988;
wire x_34989;
wire x_34990;
wire x_34991;
wire x_34992;
wire x_34993;
wire x_34994;
wire x_34995;
wire x_34996;
wire x_34997;
wire x_34998;
wire x_34999;
wire x_35000;
wire x_35001;
wire x_35002;
wire x_35003;
wire x_35004;
wire x_35005;
wire x_35006;
wire x_35007;
wire x_35008;
wire x_35009;
wire x_35010;
wire x_35011;
wire x_35012;
wire x_35013;
wire x_35014;
wire x_35015;
wire x_35016;
wire x_35017;
wire x_35018;
wire x_35019;
wire x_35020;
wire x_35021;
wire x_35022;
wire x_35023;
wire x_35024;
wire x_35025;
wire x_35026;
wire x_35027;
wire x_35028;
wire x_35029;
wire x_35030;
wire x_35031;
wire x_35032;
wire x_35033;
wire x_35034;
wire x_35035;
wire x_35036;
wire x_35037;
wire x_35038;
wire x_35039;
wire x_35040;
wire x_35041;
wire x_35042;
wire x_35043;
wire x_35044;
wire x_35045;
wire x_35046;
wire x_35047;
wire x_35048;
wire x_35049;
wire x_35050;
wire x_35051;
wire x_35052;
wire x_35053;
wire x_35054;
wire x_35055;
wire x_35056;
wire x_35057;
wire x_35058;
wire x_35059;
wire x_35060;
wire x_35061;
wire x_35062;
wire x_35063;
wire x_35064;
wire x_35065;
wire x_35066;
wire x_35067;
wire x_35068;
wire x_35069;
wire x_35070;
wire x_35071;
wire x_35072;
wire x_35073;
wire x_35074;
wire x_35075;
wire x_35076;
wire x_35077;
wire x_35078;
wire x_35079;
wire x_35080;
wire x_35081;
wire x_35082;
wire x_35083;
wire x_35084;
wire x_35085;
wire x_35086;
wire x_35087;
wire x_35088;
wire x_35089;
wire x_35090;
wire x_35091;
wire x_35092;
wire x_35093;
wire x_35094;
wire x_35095;
wire x_35096;
wire x_35097;
wire x_35098;
wire x_35099;
wire x_35100;
wire x_35101;
wire x_35102;
wire x_35103;
wire x_35104;
wire x_35105;
wire x_35106;
wire x_35107;
wire x_35108;
wire x_35109;
wire x_35110;
wire x_35111;
wire x_35112;
wire x_35113;
wire x_35114;
wire x_35115;
wire x_35116;
wire x_35117;
wire x_35118;
wire x_35119;
wire x_35120;
wire x_35121;
wire x_35122;
wire x_35123;
wire x_35124;
wire x_35125;
wire x_35126;
wire x_35127;
wire x_35128;
wire x_35129;
wire x_35130;
wire x_35131;
wire x_35132;
wire x_35133;
wire x_35134;
wire x_35135;
wire x_35136;
wire x_35137;
wire x_35138;
wire x_35139;
wire x_35140;
wire x_35141;
wire x_35142;
wire x_35143;
wire x_35144;
wire x_35145;
wire x_35146;
wire x_35147;
wire x_35148;
wire x_35149;
wire x_35150;
wire x_35151;
wire x_35152;
wire x_35153;
wire x_35154;
wire x_35155;
wire x_35156;
wire x_35157;
wire x_35158;
wire x_35159;
wire x_35160;
wire x_35161;
wire x_35162;
wire x_35163;
wire x_35164;
wire x_35165;
wire x_35166;
wire x_35167;
wire x_35168;
wire x_35169;
wire x_35170;
wire x_35171;
wire x_35172;
wire x_35173;
wire x_35174;
wire x_35175;
wire x_35176;
wire x_35177;
wire x_35178;
wire x_35179;
wire x_35180;
wire x_35181;
wire x_35182;
wire x_35183;
wire x_35184;
wire x_35185;
wire x_35186;
wire x_35187;
wire x_35188;
wire x_35189;
wire x_35190;
wire x_35191;
wire x_35192;
wire x_35193;
wire x_35194;
wire x_35195;
wire x_35196;
wire x_35197;
wire x_35198;
wire x_35199;
wire x_35200;
wire x_35201;
wire x_35202;
wire x_35203;
wire x_35204;
wire x_35205;
wire x_35206;
wire x_35207;
wire x_35208;
wire x_35209;
wire x_35210;
wire x_35211;
wire x_35212;
wire x_35213;
wire x_35214;
wire x_35215;
wire x_35216;
wire x_35217;
wire x_35218;
wire x_35219;
wire x_35220;
wire x_35221;
wire x_35222;
wire x_35223;
wire x_35224;
wire x_35225;
wire x_35226;
wire x_35227;
wire x_35228;
wire x_35229;
wire x_35230;
wire x_35231;
wire x_35232;
wire x_35233;
wire x_35234;
wire x_35235;
wire x_35236;
wire x_35237;
wire x_35238;
wire x_35239;
wire x_35240;
wire x_35241;
wire x_35242;
wire x_35243;
wire x_35244;
wire x_35245;
wire x_35246;
wire x_35247;
wire x_35248;
wire x_35249;
wire x_35250;
wire x_35251;
wire x_35252;
wire x_35253;
wire x_35254;
wire x_35255;
wire x_35256;
wire x_35257;
wire x_35258;
wire x_35259;
wire x_35260;
wire x_35261;
wire x_35262;
wire x_35263;
wire x_35264;
wire x_35265;
wire x_35266;
wire x_35267;
wire x_35268;
wire x_35269;
wire x_35270;
wire x_35271;
wire x_35272;
wire x_35273;
wire x_35274;
wire x_35275;
wire x_35276;
wire x_35277;
wire x_35278;
wire x_35279;
wire x_35280;
wire x_35281;
wire x_35282;
wire x_35283;
wire x_35284;
wire x_35285;
wire x_35286;
wire x_35287;
wire x_35288;
wire x_35289;
wire x_35290;
wire x_35291;
wire x_35292;
wire x_35293;
wire x_35294;
wire x_35295;
wire x_35296;
wire x_35297;
wire x_35298;
wire x_35299;
wire x_35300;
wire x_35301;
wire x_35302;
wire x_35303;
wire x_35304;
wire x_35305;
wire x_35306;
wire x_35307;
wire x_35308;
wire x_35309;
wire x_35310;
wire x_35311;
wire x_35312;
wire x_35313;
wire x_35314;
wire x_35315;
wire x_35316;
wire x_35317;
wire x_35318;
wire x_35319;
wire x_35320;
wire x_35321;
wire x_35322;
wire x_35323;
wire x_35324;
wire x_35325;
wire x_35326;
wire x_35327;
wire x_35328;
wire x_35329;
wire x_35330;
wire x_35331;
wire x_35332;
wire x_35333;
wire x_35334;
wire x_35335;
wire x_35336;
wire x_35337;
wire x_35338;
wire x_35339;
wire x_35340;
wire x_35341;
wire x_35342;
wire x_35343;
wire x_35344;
wire x_35345;
wire x_35346;
wire x_35347;
wire x_35348;
wire x_35349;
wire x_35350;
wire x_35351;
wire x_35352;
wire x_35353;
wire x_35354;
wire x_35355;
wire x_35356;
wire x_35357;
wire x_35358;
wire x_35359;
wire x_35360;
wire x_35361;
wire x_35362;
wire x_35363;
wire x_35364;
wire x_35365;
wire x_35366;
wire x_35367;
wire x_35368;
wire x_35369;
wire x_35370;
wire x_35371;
wire x_35372;
wire x_35373;
wire x_35374;
wire x_35375;
wire x_35376;
wire x_35377;
wire x_35378;
wire x_35379;
wire x_35380;
wire x_35381;
wire x_35382;
wire x_35383;
wire x_35384;
wire x_35385;
wire x_35386;
wire x_35387;
wire x_35388;
wire x_35389;
wire x_35390;
wire x_35391;
wire x_35392;
wire x_35393;
wire x_35394;
wire x_35395;
wire x_35396;
wire x_35397;
wire x_35398;
wire x_35399;
wire x_35400;
wire x_35401;
wire x_35402;
wire x_35403;
wire x_35404;
wire x_35405;
wire x_35406;
wire x_35407;
wire x_35408;
wire x_35409;
wire x_35410;
wire x_35411;
wire x_35412;
wire x_35413;
wire x_35414;
wire x_35415;
wire x_35416;
wire x_35417;
wire x_35418;
wire x_35419;
wire x_35420;
wire x_35421;
wire x_35422;
wire x_35423;
wire x_35424;
wire x_35425;
wire x_35426;
wire x_35427;
wire x_35428;
wire x_35429;
wire x_35430;
wire x_35431;
wire x_35432;
wire x_35433;
wire x_35434;
wire x_35435;
wire x_35436;
wire x_35437;
wire x_35438;
wire x_35439;
wire x_35440;
wire x_35441;
wire x_35442;
wire x_35443;
wire x_35444;
wire x_35445;
wire x_35446;
wire x_35447;
wire x_35448;
wire x_35449;
wire x_35450;
wire x_35451;
wire x_35452;
wire x_35453;
wire x_35454;
wire x_35455;
wire x_35456;
wire x_35457;
wire x_35458;
wire x_35459;
wire x_35460;
wire x_35461;
wire x_35462;
wire x_35463;
wire x_35464;
wire x_35465;
wire x_35466;
wire x_35467;
wire x_35468;
wire x_35469;
wire x_35470;
wire x_35471;
wire x_35472;
wire x_35473;
wire x_35474;
wire x_35475;
wire x_35476;
wire x_35477;
wire x_35478;
wire x_35479;
wire x_35480;
wire x_35481;
wire x_35482;
wire x_35483;
wire x_35484;
wire x_35485;
wire x_35486;
wire x_35487;
wire x_35488;
wire x_35489;
wire x_35490;
wire x_35491;
wire x_35492;
wire x_35493;
wire x_35494;
wire x_35495;
wire x_35496;
wire x_35497;
wire x_35498;
wire x_35499;
wire x_35500;
wire x_35501;
wire x_35502;
wire x_35503;
wire x_35504;
wire x_35505;
wire x_35506;
wire x_35507;
wire x_35508;
wire x_35509;
wire x_35510;
wire x_35511;
wire x_35512;
wire x_35513;
wire x_35514;
wire x_35515;
wire x_35516;
wire x_35517;
wire x_35518;
wire x_35519;
wire x_35520;
wire x_35521;
wire x_35522;
wire x_35523;
wire x_35524;
wire x_35525;
wire x_35526;
wire x_35527;
wire x_35528;
wire x_35529;
wire x_35530;
wire x_35531;
wire x_35532;
wire x_35533;
wire x_35534;
wire x_35535;
wire x_35536;
wire x_35537;
wire x_35538;
wire x_35539;
wire x_35540;
wire x_35541;
wire x_35542;
wire x_35543;
wire x_35544;
wire x_35545;
wire x_35546;
wire x_35547;
wire x_35548;
wire x_35549;
wire x_35550;
wire x_35551;
wire x_35552;
wire x_35553;
wire x_35554;
wire x_35555;
wire x_35556;
wire x_35557;
wire x_35558;
wire x_35559;
wire x_35560;
wire x_35561;
wire x_35562;
wire x_35563;
wire x_35564;
wire x_35565;
wire x_35566;
wire x_35567;
wire x_35568;
wire x_35569;
wire x_35570;
wire x_35571;
wire x_35572;
wire x_35573;
wire x_35574;
wire x_35575;
wire x_35576;
wire x_35577;
wire x_35578;
wire x_35579;
wire x_35580;
wire x_35581;
wire x_35582;
wire x_35583;
wire x_35584;
wire x_35585;
wire x_35586;
wire x_35587;
wire x_35588;
wire x_35589;
wire x_35590;
wire x_35591;
wire x_35592;
wire x_35593;
wire x_35594;
wire x_35595;
wire x_35596;
wire x_35597;
wire x_35598;
wire x_35599;
wire x_35600;
wire x_35601;
wire x_35602;
wire x_35603;
wire x_35604;
wire x_35605;
wire x_35606;
wire x_35607;
wire x_35608;
wire x_35609;
wire x_35610;
wire x_35611;
wire x_35612;
wire x_35613;
wire x_35614;
wire x_35615;
wire x_35616;
wire x_35617;
wire x_35618;
wire x_35619;
wire x_35620;
wire x_35621;
wire x_35622;
wire x_35623;
wire x_35624;
wire x_35625;
wire x_35626;
wire x_35627;
wire x_35628;
wire x_35629;
wire x_35630;
wire x_35631;
wire x_35632;
wire x_35633;
wire x_35634;
wire x_35635;
wire x_35636;
wire x_35637;
wire x_35638;
wire x_35639;
wire x_35640;
wire x_35641;
wire x_35642;
wire x_35643;
wire x_35644;
wire x_35645;
wire x_35646;
wire x_35647;
wire x_35648;
wire x_35649;
wire x_35650;
wire x_35651;
wire x_35652;
wire x_35653;
wire x_35654;
wire x_35655;
wire x_35656;
wire x_35657;
wire x_35658;
wire x_35659;
wire x_35660;
wire x_35661;
wire x_35662;
wire x_35663;
wire x_35664;
wire x_35665;
wire x_35666;
wire x_35667;
wire x_35668;
wire x_35669;
wire x_35670;
wire x_35671;
wire x_35672;
wire x_35673;
wire x_35674;
wire x_35675;
wire x_35676;
wire x_35677;
wire x_35678;
wire x_35679;
wire x_35680;
wire x_35681;
wire x_35682;
wire x_35683;
wire x_35684;
wire x_35685;
wire x_35686;
wire x_35687;
wire x_35688;
wire x_35689;
wire x_35690;
wire x_35691;
wire x_35692;
wire x_35693;
wire x_35694;
wire x_35695;
wire x_35696;
wire x_35697;
wire x_35698;
wire x_35699;
wire x_35700;
wire x_35701;
wire x_35702;
wire x_35703;
wire x_35704;
wire x_35705;
wire x_35706;
wire x_35707;
wire x_35708;
wire x_35709;
wire x_35710;
wire x_35711;
wire x_35712;
wire x_35713;
wire x_35714;
wire x_35715;
wire x_35716;
wire x_35717;
wire x_35718;
wire x_35719;
wire x_35720;
wire x_35721;
wire x_35722;
wire x_35723;
wire x_35724;
wire x_35725;
wire x_35726;
wire x_35727;
wire x_35728;
wire x_35729;
wire x_35730;
wire x_35731;
wire x_35732;
wire x_35733;
wire x_35734;
wire x_35735;
wire x_35736;
wire x_35737;
wire x_35738;
wire x_35739;
wire x_35740;
wire x_35741;
wire x_35742;
wire x_35743;
wire x_35744;
wire x_35745;
wire x_35746;
wire x_35747;
wire x_35748;
wire x_35749;
wire x_35750;
wire x_35751;
wire x_35752;
wire x_35753;
wire x_35754;
wire x_35755;
wire x_35756;
wire x_35757;
wire x_35758;
wire x_35759;
wire x_35760;
wire x_35761;
wire x_35762;
wire x_35763;
wire x_35764;
wire x_35765;
wire x_35766;
wire x_35767;
wire x_35768;
wire x_35769;
wire x_35770;
wire x_35771;
wire x_35772;
wire x_35773;
wire x_35774;
wire x_35775;
wire x_35776;
wire x_35777;
wire x_35778;
wire x_35779;
wire x_35780;
wire x_35781;
wire x_35782;
wire x_35783;
wire x_35784;
wire x_35785;
wire x_35786;
wire x_35787;
wire x_35788;
wire x_35789;
wire x_35790;
wire x_35791;
wire x_35792;
wire x_35793;
wire x_35794;
wire x_35795;
wire x_35796;
wire x_35797;
wire x_35798;
wire x_35799;
wire x_35800;
wire x_35801;
wire x_35802;
wire x_35803;
wire x_35804;
wire x_35805;
wire x_35806;
wire x_35807;
wire x_35808;
wire x_35809;
wire x_35810;
wire x_35811;
wire x_35812;
wire x_35813;
wire x_35814;
wire x_35815;
wire x_35816;
wire x_35817;
wire x_35818;
wire x_35819;
wire x_35820;
wire x_35821;
wire x_35822;
wire x_35823;
wire x_35824;
wire x_35825;
wire x_35826;
wire x_35827;
wire x_35828;
wire x_35829;
wire x_35830;
wire x_35831;
wire x_35832;
wire x_35833;
wire x_35834;
wire x_35835;
wire x_35836;
wire x_35837;
wire x_35838;
wire x_35839;
wire x_35840;
wire x_35841;
wire x_35842;
wire x_35843;
wire x_35844;
wire x_35845;
wire x_35846;
wire x_35847;
wire x_35848;
wire x_35849;
wire x_35850;
wire x_35851;
wire x_35852;
wire x_35853;
wire x_35854;
wire x_35855;
wire x_35856;
wire x_35857;
wire x_35858;
wire x_35859;
wire x_35860;
wire x_35861;
wire x_35862;
wire x_35863;
wire x_35864;
wire x_35865;
wire x_35866;
wire x_35867;
wire x_35868;
wire x_35869;
wire x_35870;
wire x_35871;
wire x_35872;
wire x_35873;
wire x_35874;
wire x_35875;
wire x_35876;
wire x_35877;
wire x_35878;
wire x_35879;
wire x_35880;
wire x_35881;
wire x_35882;
wire x_35883;
wire x_35884;
wire x_35885;
wire x_35886;
wire x_35887;
wire x_35888;
wire x_35889;
wire x_35890;
wire x_35891;
wire x_35892;
wire x_35893;
wire x_35894;
wire x_35895;
wire x_35896;
wire x_35897;
wire x_35898;
wire x_35899;
wire x_35900;
wire x_35901;
wire x_35902;
wire x_35903;
wire x_35904;
wire x_35905;
wire x_35906;
wire x_35907;
wire x_35908;
wire x_35909;
wire x_35910;
wire x_35911;
wire x_35912;
wire x_35913;
wire x_35914;
wire x_35915;
wire x_35916;
wire x_35917;
wire x_35918;
wire x_35919;
wire x_35920;
wire x_35921;
wire x_35922;
wire x_35923;
wire x_35924;
wire x_35925;
wire x_35926;
wire x_35927;
wire x_35928;
wire x_35929;
wire x_35930;
wire x_35931;
wire x_35932;
wire x_35933;
wire x_35934;
wire x_35935;
wire x_35936;
wire x_35937;
wire x_35938;
wire x_35939;
wire x_35940;
wire x_35941;
wire x_35942;
wire x_35943;
wire x_35944;
wire x_35945;
wire x_35946;
wire x_35947;
wire x_35948;
wire x_35949;
wire x_35950;
wire x_35951;
wire x_35952;
wire x_35953;
wire x_35954;
wire x_35955;
wire x_35956;
wire x_35957;
wire x_35958;
wire x_35959;
wire x_35960;
wire x_35961;
wire x_35962;
wire x_35963;
wire x_35964;
wire x_35965;
wire x_35966;
wire x_35967;
wire x_35968;
wire x_35969;
wire x_35970;
wire x_35971;
wire x_35972;
wire x_35973;
wire x_35974;
wire x_35975;
wire x_35976;
wire x_35977;
wire x_35978;
wire x_35979;
wire x_35980;
wire x_35981;
wire x_35982;
wire x_35983;
wire x_35984;
wire x_35985;
wire x_35986;
wire x_35987;
wire x_35988;
wire x_35989;
wire x_35990;
wire x_35991;
wire x_35992;
wire x_35993;
wire x_35994;
wire x_35995;
wire x_35996;
wire x_35997;
wire x_35998;
wire x_35999;
wire x_36000;
wire x_36001;
wire x_36002;
wire x_36003;
wire x_36004;
wire x_36005;
wire x_36006;
wire x_36007;
wire x_36008;
wire x_36009;
wire x_36010;
wire x_36011;
wire x_36012;
wire x_36013;
wire x_36014;
wire x_36015;
wire x_36016;
wire x_36017;
wire x_36018;
wire x_36019;
wire x_36020;
wire x_36021;
wire x_36022;
wire x_36023;
wire x_36024;
wire x_36025;
wire x_36026;
wire x_36027;
wire x_36028;
wire x_36029;
wire x_36030;
wire x_36031;
wire x_36032;
wire x_36033;
wire x_36034;
wire x_36035;
wire x_36036;
wire x_36037;
wire x_36038;
wire x_36039;
wire x_36040;
wire x_36041;
wire x_36042;
wire x_36043;
wire x_36044;
wire x_36045;
wire x_36046;
wire x_36047;
wire x_36048;
wire x_36049;
wire x_36050;
wire x_36051;
wire x_36052;
wire x_36053;
wire x_36054;
wire x_36055;
wire x_36056;
wire x_36057;
wire x_36058;
wire x_36059;
wire x_36060;
wire x_36061;
wire x_36062;
wire x_36063;
wire x_36064;
wire x_36065;
wire x_36066;
wire x_36067;
wire x_36068;
wire x_36069;
wire x_36070;
wire x_36071;
wire x_36072;
wire x_36073;
wire x_36074;
wire x_36075;
wire x_36076;
wire x_36077;
wire x_36078;
wire x_36079;
wire x_36080;
wire x_36081;
wire x_36082;
wire x_36083;
wire x_36084;
wire x_36085;
wire x_36086;
wire x_36087;
wire x_36088;
wire x_36089;
wire x_36090;
wire x_36091;
wire x_36092;
wire x_36093;
wire x_36094;
wire x_36095;
wire x_36096;
wire x_36097;
wire x_36098;
wire x_36099;
wire x_36100;
wire x_36101;
wire x_36102;
wire x_36103;
wire x_36104;
wire x_36105;
wire x_36106;
wire x_36107;
wire x_36108;
wire x_36109;
wire x_36110;
wire x_36111;
wire x_36112;
wire x_36113;
wire x_36114;
wire x_36115;
wire x_36116;
wire x_36117;
wire x_36118;
wire x_36119;
wire x_36120;
wire x_36121;
wire x_36122;
wire x_36123;
wire x_36124;
wire x_36125;
wire x_36126;
wire x_36127;
wire x_36128;
wire x_36129;
wire x_36130;
wire x_36131;
wire x_36132;
wire x_36133;
wire x_36134;
wire x_36135;
wire x_36136;
wire x_36137;
wire x_36138;
wire x_36139;
wire x_36140;
wire x_36141;
wire x_36142;
wire x_36143;
wire x_36144;
wire x_36145;
wire x_36146;
wire x_36147;
wire x_36148;
wire x_36149;
wire x_36150;
wire x_36151;
wire x_36152;
wire x_36153;
wire x_36154;
wire x_36155;
wire x_36156;
wire x_36157;
wire x_36158;
wire x_36159;
wire x_36160;
wire x_36161;
wire x_36162;
wire x_36163;
wire x_36164;
wire x_36165;
wire x_36166;
wire x_36167;
wire x_36168;
wire x_36169;
wire x_36170;
wire x_36171;
wire x_36172;
wire x_36173;
wire x_36174;
wire x_36175;
wire x_36176;
wire x_36177;
wire x_36178;
wire x_36179;
wire x_36180;
wire x_36181;
wire x_36182;
wire x_36183;
wire x_36184;
wire x_36185;
wire x_36186;
wire x_36187;
wire x_36188;
wire x_36189;
wire x_36190;
wire x_36191;
wire x_36192;
wire x_36193;
wire x_36194;
wire x_36195;
wire x_36196;
wire x_36197;
wire x_36198;
wire x_36199;
wire x_36200;
wire x_36201;
wire x_36202;
wire x_36203;
wire x_36204;
wire x_36205;
wire x_36206;
wire x_36207;
wire x_36208;
wire x_36209;
wire x_36210;
wire x_36211;
wire x_36212;
wire x_36213;
wire x_36214;
wire x_36215;
wire x_36216;
wire x_36217;
wire x_36218;
wire x_36219;
wire x_36220;
wire x_36221;
wire x_36222;
wire x_36223;
wire x_36224;
wire x_36225;
wire x_36226;
wire x_36227;
wire x_36228;
wire x_36229;
wire x_36230;
wire x_36231;
wire x_36232;
wire x_36233;
wire x_36234;
wire x_36235;
wire x_36236;
wire x_36237;
wire x_36238;
wire x_36239;
wire x_36240;
wire x_36241;
wire x_36242;
wire x_36243;
wire x_36244;
wire x_36245;
wire x_36246;
wire x_36247;
wire x_36248;
wire x_36249;
wire x_36250;
wire x_36251;
wire x_36252;
wire x_36253;
wire x_36254;
wire x_36255;
wire x_36256;
wire x_36257;
wire x_36258;
wire x_36259;
wire x_36260;
wire x_36261;
wire x_36262;
wire x_36263;
wire x_36264;
wire x_36265;
wire x_36266;
wire x_36267;
wire x_36268;
wire x_36269;
wire x_36270;
wire x_36271;
wire x_36272;
wire x_36273;
wire x_36274;
wire x_36275;
wire x_36276;
wire x_36277;
wire x_36278;
wire x_36279;
wire x_36280;
wire x_36281;
wire x_36282;
wire x_36283;
wire x_36284;
wire x_36285;
wire x_36286;
wire x_36287;
wire x_36288;
wire x_36289;
wire x_36290;
wire x_36291;
wire x_36292;
wire x_36293;
wire x_36294;
wire x_36295;
wire x_36296;
wire x_36297;
wire x_36298;
wire x_36299;
wire x_36300;
wire x_36301;
wire x_36302;
wire x_36303;
wire x_36304;
wire x_36305;
wire x_36306;
wire x_36307;
wire x_36308;
wire x_36309;
wire x_36310;
wire x_36311;
wire x_36312;
wire x_36313;
wire x_36314;
wire x_36315;
wire x_36316;
wire x_36317;
wire x_36318;
wire x_36319;
wire x_36320;
wire x_36321;
wire x_36322;
wire x_36323;
wire x_36324;
wire x_36325;
wire x_36326;
wire x_36327;
wire x_36328;
wire x_36329;
wire x_36330;
wire x_36331;
wire x_36332;
wire x_36333;
wire x_36334;
wire x_36335;
wire x_36336;
wire x_36337;
wire x_36338;
wire x_36339;
wire x_36340;
wire x_36341;
wire x_36342;
wire x_36343;
wire x_36344;
wire x_36345;
wire x_36346;
wire x_36347;
wire x_36348;
wire x_36349;
wire x_36350;
wire x_36351;
wire x_36352;
wire x_36353;
wire x_36354;
wire x_36355;
wire x_36356;
wire x_36357;
wire x_36358;
wire x_36359;
wire x_36360;
wire x_36361;
wire x_36362;
wire x_36363;
wire x_36364;
wire x_36365;
wire x_36366;
wire x_36367;
wire x_36368;
wire x_36369;
wire x_36370;
wire x_36371;
wire x_36372;
wire x_36373;
wire x_36374;
wire x_36375;
wire x_36376;
wire x_36377;
wire x_36378;
wire x_36379;
wire x_36380;
wire x_36381;
wire x_36382;
wire x_36383;
wire x_36384;
wire x_36385;
wire x_36386;
wire x_36387;
wire x_36388;
wire x_36389;
wire x_36390;
wire x_36391;
wire x_36392;
wire x_36393;
wire x_36394;
wire x_36395;
wire x_36396;
wire x_36397;
wire x_36398;
wire x_36399;
wire x_36400;
wire x_36401;
wire x_36402;
wire x_36403;
wire x_36404;
wire x_36405;
wire x_36406;
wire x_36407;
wire x_36408;
wire x_36409;
wire x_36410;
wire x_36411;
wire x_36412;
wire x_36413;
wire x_36414;
wire x_36415;
wire x_36416;
wire x_36417;
wire x_36418;
wire x_36419;
wire x_36420;
wire x_36421;
wire x_36422;
wire x_36423;
wire x_36424;
wire x_36425;
wire x_36426;
wire x_36427;
wire x_36428;
wire x_36429;
wire x_36430;
wire x_36431;
wire x_36432;
wire x_36433;
wire x_36434;
wire x_36435;
wire x_36436;
wire x_36437;
wire x_36438;
wire x_36439;
wire x_36440;
wire x_36441;
wire x_36442;
wire x_36443;
wire x_36444;
wire x_36445;
wire x_36446;
wire x_36447;
wire x_36448;
wire x_36449;
wire x_36450;
wire x_36451;
wire x_36452;
wire x_36453;
wire x_36454;
wire x_36455;
wire x_36456;
wire x_36457;
wire x_36458;
wire x_36459;
wire x_36460;
wire x_36461;
wire x_36462;
wire x_36463;
wire x_36464;
wire x_36465;
wire x_36466;
wire x_36467;
wire x_36468;
wire x_36469;
wire x_36470;
wire x_36471;
wire x_36472;
wire x_36473;
wire x_36474;
wire x_36475;
wire x_36476;
wire x_36477;
wire x_36478;
wire x_36479;
wire x_36480;
wire x_36481;
wire x_36482;
wire x_36483;
wire x_36484;
wire x_36485;
wire x_36486;
wire x_36487;
wire x_36488;
wire x_36489;
wire x_36490;
wire x_36491;
wire x_36492;
wire x_36493;
wire x_36494;
wire x_36495;
wire x_36496;
wire x_36497;
wire x_36498;
wire x_36499;
wire x_36500;
wire x_36501;
wire x_36502;
wire x_36503;
wire x_36504;
wire x_36505;
wire x_36506;
wire x_36507;
wire x_36508;
wire x_36509;
wire x_36510;
wire x_36511;
wire x_36512;
wire x_36513;
wire x_36514;
wire x_36515;
wire x_36516;
wire x_36517;
wire x_36518;
wire x_36519;
wire x_36520;
wire x_36521;
wire x_36522;
wire x_36523;
wire x_36524;
wire x_36525;
wire x_36526;
wire x_36527;
wire x_36528;
wire x_36529;
wire x_36530;
wire x_36531;
wire x_36532;
wire x_36533;
wire x_36534;
wire x_36535;
wire x_36536;
wire x_36537;
wire x_36538;
wire x_36539;
wire x_36540;
wire x_36541;
wire x_36542;
wire x_36543;
wire x_36544;
wire x_36545;
wire x_36546;
wire x_36547;
wire x_36548;
wire x_36549;
wire x_36550;
wire x_36551;
wire x_36552;
wire x_36553;
wire x_36554;
wire x_36555;
wire x_36556;
wire x_36557;
wire x_36558;
wire x_36559;
wire x_36560;
wire x_36561;
wire x_36562;
wire x_36563;
wire x_36564;
wire x_36565;
wire x_36566;
wire x_36567;
wire x_36568;
wire x_36569;
wire x_36570;
wire x_36571;
wire x_36572;
wire x_36573;
wire x_36574;
wire x_36575;
wire x_36576;
wire x_36577;
wire x_36578;
wire x_36579;
wire x_36580;
wire x_36581;
wire x_36582;
wire x_36583;
wire x_36584;
wire x_36585;
wire x_36586;
wire x_36587;
wire x_36588;
wire x_36589;
wire x_36590;
wire x_36591;
wire x_36592;
wire x_36593;
wire x_36594;
wire x_36595;
wire x_36596;
wire x_36597;
wire x_36598;
wire x_36599;
wire x_36600;
wire x_36601;
wire x_36602;
wire x_36603;
wire x_36604;
wire x_36605;
wire x_36606;
wire x_36607;
wire x_36608;
wire x_36609;
wire x_36610;
wire x_36611;
wire x_36612;
wire x_36613;
wire x_36614;
wire x_36615;
wire x_36616;
wire x_36617;
wire x_36618;
wire x_36619;
wire x_36620;
wire x_36621;
wire x_36622;
wire x_36623;
wire x_36624;
wire x_36625;
wire x_36626;
wire x_36627;
wire x_36628;
wire x_36629;
wire x_36630;
wire x_36631;
wire x_36632;
wire x_36633;
wire x_36634;
wire x_36635;
wire x_36636;
wire x_36637;
wire x_36638;
wire x_36639;
wire x_36640;
wire x_36641;
wire x_36642;
wire x_36643;
wire x_36644;
wire x_36645;
wire x_36646;
wire x_36647;
wire x_36648;
wire x_36649;
wire x_36650;
wire x_36651;
wire x_36652;
wire x_36653;
wire x_36654;
wire x_36655;
wire x_36656;
wire x_36657;
wire x_36658;
wire x_36659;
wire x_36660;
wire x_36661;
wire x_36662;
wire x_36663;
wire x_36664;
wire x_36665;
wire x_36666;
wire x_36667;
wire x_36668;
wire x_36669;
wire x_36670;
wire x_36671;
wire x_36672;
wire x_36673;
wire x_36674;
wire x_36675;
wire x_36676;
wire x_36677;
wire x_36678;
wire x_36679;
wire x_36680;
wire x_36681;
wire x_36682;
wire x_36683;
wire x_36684;
wire x_36685;
wire x_36686;
wire x_36687;
wire x_36688;
wire x_36689;
wire x_36690;
wire x_36691;
wire x_36692;
wire x_36693;
wire x_36694;
wire x_36695;
wire x_36696;
wire x_36697;
wire x_36698;
wire x_36699;
wire x_36700;
wire x_36701;
wire x_36702;
wire x_36703;
wire x_36704;
wire x_36705;
wire x_36706;
wire x_36707;
wire x_36708;
wire x_36709;
wire x_36710;
wire x_36711;
wire x_36712;
wire x_36713;
wire x_36714;
wire x_36715;
wire x_36716;
wire x_36717;
wire x_36718;
wire x_36719;
wire x_36720;
wire x_36721;
wire x_36722;
wire x_36723;
wire x_36724;
wire x_36725;
wire x_36726;
wire x_36727;
wire x_36728;
wire x_36729;
wire x_36730;
wire x_36731;
wire x_36732;
wire x_36733;
wire x_36734;
wire x_36735;
wire x_36736;
wire x_36737;
wire x_36738;
wire x_36739;
wire x_36740;
wire x_36741;
wire x_36742;
wire x_36743;
wire x_36744;
wire x_36745;
wire x_36746;
wire x_36747;
wire x_36748;
wire x_36749;
wire x_36750;
wire x_36751;
wire x_36752;
wire x_36753;
wire x_36754;
wire x_36755;
wire x_36756;
wire x_36757;
wire x_36758;
wire x_36759;
wire x_36760;
wire x_36761;
wire x_36762;
wire x_36763;
wire x_36764;
wire x_36765;
wire x_36766;
wire x_36767;
wire x_36768;
wire x_36769;
wire x_36770;
wire x_36771;
wire x_36772;
wire x_36773;
wire x_36774;
wire x_36775;
wire x_36776;
wire x_36777;
wire x_36778;
wire x_36779;
wire x_36780;
wire x_36781;
wire x_36782;
wire x_36783;
wire x_36784;
wire x_36785;
wire x_36786;
wire x_36787;
wire x_36788;
wire x_36789;
wire x_36790;
wire x_36791;
wire x_36792;
wire x_36793;
wire x_36794;
wire x_36795;
wire x_36796;
wire x_36797;
wire x_36798;
wire x_36799;
wire x_36800;
wire x_36801;
wire x_36802;
wire x_36803;
wire x_36804;
wire x_36805;
wire x_36806;
wire x_36807;
wire x_36808;
wire x_36809;
wire x_36810;
wire x_36811;
wire x_36812;
wire x_36813;
wire x_36814;
wire x_36815;
wire x_36816;
wire x_36817;
wire x_36818;
wire x_36819;
wire x_36820;
wire x_36821;
wire x_36822;
wire x_36823;
wire x_36824;
wire x_36825;
wire x_36826;
wire x_36827;
wire x_36828;
wire x_36829;
wire x_36830;
wire x_36831;
wire x_36832;
wire x_36833;
wire x_36834;
wire x_36835;
wire x_36836;
wire x_36837;
wire x_36838;
wire x_36839;
wire x_36840;
wire x_36841;
wire x_36842;
wire x_36843;
wire x_36844;
wire x_36845;
wire x_36846;
wire x_36847;
wire x_36848;
wire x_36849;
wire x_36850;
wire x_36851;
wire x_36852;
wire x_36853;
wire x_36854;
wire x_36855;
wire x_36856;
wire x_36857;
wire x_36858;
wire x_36859;
wire x_36860;
wire x_36861;
wire x_36862;
wire x_36863;
wire x_36864;
wire x_36865;
wire x_36866;
wire x_36867;
wire x_36868;
wire x_36869;
wire x_36870;
wire x_36871;
wire x_36872;
wire x_36873;
wire x_36874;
wire x_36875;
wire x_36876;
wire x_36877;
wire x_36878;
wire x_36879;
wire x_36880;
wire x_36881;
wire x_36882;
wire x_36883;
wire x_36884;
wire x_36885;
wire x_36886;
wire x_36887;
wire x_36888;
wire x_36889;
wire x_36890;
wire x_36891;
wire x_36892;
wire x_36893;
wire x_36894;
wire x_36895;
wire x_36896;
wire x_36897;
wire x_36898;
wire x_36899;
wire x_36900;
wire x_36901;
wire x_36902;
wire x_36903;
wire x_36904;
wire x_36905;
wire x_36906;
wire x_36907;
wire x_36908;
wire x_36909;
wire x_36910;
wire x_36911;
wire x_36912;
wire x_36913;
wire x_36914;
wire x_36915;
wire x_36916;
wire x_36917;
wire x_36918;
wire x_36919;
wire x_36920;
wire x_36921;
wire x_36922;
wire x_36923;
wire x_36924;
wire x_36925;
wire x_36926;
wire x_36927;
wire x_36928;
wire x_36929;
wire x_36930;
wire x_36931;
wire x_36932;
wire x_36933;
wire x_36934;
wire x_36935;
wire x_36936;
wire x_36937;
wire x_36938;
wire x_36939;
wire x_36940;
wire x_36941;
wire x_36942;
wire x_36943;
wire x_36944;
wire x_36945;
wire x_36946;
wire x_36947;
wire x_36948;
wire x_36949;
wire x_36950;
wire x_36951;
wire x_36952;
wire x_36953;
wire x_36954;
wire x_36955;
wire x_36956;
wire x_36957;
wire x_36958;
wire x_36959;
wire x_36960;
wire x_36961;
wire x_36962;
wire x_36963;
wire x_36964;
wire x_36965;
wire x_36966;
wire x_36967;
wire x_36968;
wire x_36969;
wire x_36970;
wire x_36971;
wire x_36972;
wire x_36973;
wire x_36974;
wire x_36975;
wire x_36976;
wire x_36977;
wire x_36978;
wire x_36979;
wire x_36980;
wire x_36981;
wire x_36982;
wire x_36983;
wire x_36984;
wire x_36985;
wire x_36986;
wire x_36987;
wire x_36988;
wire x_36989;
wire x_36990;
wire x_36991;
wire x_36992;
wire x_36993;
wire x_36994;
wire x_36995;
wire x_36996;
wire x_36997;
wire x_36998;
wire x_36999;
wire x_37000;
wire x_37001;
wire x_37002;
wire x_37003;
wire x_37004;
wire x_37005;
wire x_37006;
wire x_37007;
wire x_37008;
wire x_37009;
wire x_37010;
wire x_37011;
wire x_37012;
wire x_37013;
wire x_37014;
wire x_37015;
wire x_37016;
wire x_37017;
wire x_37018;
wire x_37019;
wire x_37020;
wire x_37021;
wire x_37022;
wire x_37023;
wire x_37024;
wire x_37025;
wire x_37026;
wire x_37027;
wire x_37028;
wire x_37029;
wire x_37030;
wire x_37031;
wire x_37032;
wire x_37033;
wire x_37034;
wire x_37035;
wire x_37036;
wire x_37037;
wire x_37038;
wire x_37039;
wire x_37040;
wire x_37041;
wire x_37042;
wire x_37043;
wire x_37044;
wire x_37045;
wire x_37046;
wire x_37047;
wire x_37048;
wire x_37049;
wire x_37050;
wire x_37051;
wire x_37052;
wire x_37053;
wire x_37054;
wire x_37055;
wire x_37056;
wire x_37057;
wire x_37058;
wire x_37059;
wire x_37060;
wire x_37061;
wire x_37062;
wire x_37063;
wire x_37064;
wire x_37065;
wire x_37066;
wire x_37067;
wire x_37068;
wire x_37069;
wire x_37070;
wire x_37071;
wire x_37072;
wire x_37073;
wire x_37074;
wire x_37075;
wire x_37076;
wire x_37077;
wire x_37078;
wire x_37079;
wire x_37080;
wire x_37081;
wire x_37082;
wire x_37083;
wire x_37084;
wire x_37085;
wire x_37086;
wire x_37087;
wire x_37088;
wire x_37089;
wire x_37090;
wire x_37091;
wire x_37092;
wire x_37093;
wire x_37094;
wire x_37095;
wire x_37096;
wire x_37097;
wire x_37098;
wire x_37099;
wire x_37100;
wire x_37101;
wire x_37102;
wire x_37103;
wire x_37104;
wire x_37105;
wire x_37106;
wire x_37107;
wire x_37108;
wire x_37109;
wire x_37110;
wire x_37111;
wire x_37112;
wire x_37113;
wire x_37114;
wire x_37115;
wire x_37116;
wire x_37117;
wire x_37118;
wire x_37119;
wire x_37120;
wire x_37121;
wire x_37122;
wire x_37123;
wire x_37124;
wire x_37125;
wire x_37126;
wire x_37127;
wire x_37128;
wire x_37129;
wire x_37130;
wire x_37131;
wire x_37132;
wire x_37133;
wire x_37134;
wire x_37135;
wire x_37136;
wire x_37137;
wire x_37138;
wire x_37139;
wire x_37140;
wire x_37141;
wire x_37142;
wire x_37143;
wire x_37144;
wire x_37145;
wire x_37146;
wire x_37147;
wire x_37148;
wire x_37149;
wire x_37150;
wire x_37151;
wire x_37152;
wire x_37153;
wire x_37154;
wire x_37155;
wire x_37156;
wire x_37157;
wire x_37158;
wire x_37159;
wire x_37160;
wire x_37161;
wire x_37162;
wire x_37163;
wire x_37164;
wire x_37165;
wire x_37166;
wire x_37167;
wire x_37168;
wire x_37169;
wire x_37170;
wire x_37171;
wire x_37172;
wire x_37173;
wire x_37174;
wire x_37175;
wire x_37176;
wire x_37177;
wire x_37178;
wire x_37179;
wire x_37180;
wire x_37181;
wire x_37182;
wire x_37183;
wire x_37184;
wire x_37185;
wire x_37186;
wire x_37187;
wire x_37188;
wire x_37189;
wire x_37190;
wire x_37191;
wire x_37192;
wire x_37193;
wire x_37194;
wire x_37195;
wire x_37196;
wire x_37197;
wire x_37198;
wire x_37199;
wire x_37200;
wire x_37201;
wire x_37202;
wire x_37203;
wire x_37204;
wire x_37205;
wire x_37206;
wire x_37207;
wire x_37208;
wire x_37209;
wire x_37210;
wire x_37211;
wire x_37212;
wire x_37213;
wire x_37214;
wire x_37215;
wire x_37216;
wire x_37217;
wire x_37218;
wire x_37219;
wire x_37220;
wire x_37221;
wire x_37222;
wire x_37223;
wire x_37224;
wire x_37225;
wire x_37226;
wire x_37227;
wire x_37228;
wire x_37229;
wire x_37230;
wire x_37231;
wire x_37232;
wire x_37233;
wire x_37234;
wire x_37235;
wire x_37236;
wire x_37237;
wire x_37238;
wire x_37239;
wire x_37240;
wire x_37241;
wire x_37242;
wire x_37243;
wire x_37244;
wire x_37245;
wire x_37246;
wire x_37247;
wire x_37248;
wire x_37249;
wire x_37250;
wire x_37251;
wire x_37252;
wire x_37253;
wire x_37254;
wire x_37255;
wire x_37256;
wire x_37257;
wire x_37258;
wire x_37259;
wire x_37260;
wire x_37261;
wire x_37262;
wire x_37263;
wire x_37264;
wire x_37265;
wire x_37266;
wire x_37267;
wire x_37268;
wire x_37269;
wire x_37270;
wire x_37271;
wire x_37272;
wire x_37273;
wire x_37274;
wire x_37275;
wire x_37276;
wire x_37277;
wire x_37278;
wire x_37279;
wire x_37280;
wire x_37281;
wire x_37282;
wire x_37283;
wire x_37284;
wire x_37285;
wire x_37286;
wire x_37287;
wire x_37288;
wire x_37289;
wire x_37290;
wire x_37291;
wire x_37292;
wire x_37293;
wire x_37294;
wire x_37295;
wire x_37296;
wire x_37297;
wire x_37298;
wire x_37299;
wire x_37300;
wire x_37301;
wire x_37302;
wire x_37303;
wire x_37304;
wire x_37305;
wire x_37306;
wire x_37307;
wire x_37308;
wire x_37309;
wire x_37310;
wire x_37311;
wire x_37312;
wire x_37313;
wire x_37314;
wire x_37315;
wire x_37316;
wire x_37317;
wire x_37318;
wire x_37319;
wire x_37320;
wire x_37321;
wire x_37322;
wire x_37323;
wire x_37324;
wire x_37325;
wire x_37326;
wire x_37327;
wire x_37328;
wire x_37329;
wire x_37330;
wire x_37331;
wire x_37332;
wire x_37333;
wire x_37334;
wire x_37335;
wire x_37336;
wire x_37337;
wire x_37338;
wire x_37339;
wire x_37340;
wire x_37341;
wire x_37342;
wire x_37343;
wire x_37344;
wire x_37345;
wire x_37346;
wire x_37347;
wire x_37348;
wire x_37349;
wire x_37350;
wire x_37351;
wire x_37352;
wire x_37353;
wire x_37354;
wire x_37355;
wire x_37356;
wire x_37357;
wire x_37358;
wire x_37359;
wire x_37360;
wire x_37361;
wire x_37362;
wire x_37363;
wire x_37364;
wire x_37365;
wire x_37366;
wire x_37367;
wire x_37368;
wire x_37369;
wire x_37370;
wire x_37371;
wire x_37372;
wire x_37373;
wire x_37374;
wire x_37375;
wire x_37376;
wire x_37377;
wire x_37378;
wire x_37379;
wire x_37380;
wire x_37381;
wire x_37382;
wire x_37383;
wire x_37384;
wire x_37385;
wire x_37386;
wire x_37387;
wire x_37388;
wire x_37389;
wire x_37390;
wire x_37391;
wire x_37392;
wire x_37393;
wire x_37394;
wire x_37395;
wire x_37396;
wire x_37397;
wire x_37398;
wire x_37399;
wire x_37400;
wire x_37401;
wire x_37402;
wire x_37403;
wire x_37404;
wire x_37405;
wire x_37406;
wire x_37407;
wire x_37408;
wire x_37409;
wire x_37410;
wire x_37411;
wire x_37412;
wire x_37413;
wire x_37414;
wire x_37415;
wire x_37416;
wire x_37417;
wire x_37418;
wire x_37419;
wire x_37420;
wire x_37421;
wire x_37422;
wire x_37423;
wire x_37424;
wire x_37425;
wire x_37426;
wire x_37427;
wire x_37428;
wire x_37429;
wire x_37430;
wire x_37431;
wire x_37432;
wire x_37433;
wire x_37434;
wire x_37435;
wire x_37436;
wire x_37437;
wire x_37438;
wire x_37439;
wire x_37440;
wire x_37441;
wire x_37442;
wire x_37443;
wire x_37444;
wire x_37445;
wire x_37446;
wire x_37447;
wire x_37448;
wire x_37449;
wire x_37450;
wire x_37451;
wire x_37452;
wire x_37453;
wire x_37454;
wire x_37455;
wire x_37456;
wire x_37457;
wire x_37458;
wire x_37459;
wire x_37460;
wire x_37461;
wire x_37462;
wire x_37463;
wire x_37464;
wire x_37465;
wire x_37466;
wire x_37467;
wire x_37468;
wire x_37469;
wire x_37470;
wire x_37471;
wire x_37472;
wire x_37473;
wire x_37474;
wire x_37475;
wire x_37476;
wire x_37477;
wire x_37478;
wire x_37479;
wire x_37480;
wire x_37481;
wire x_37482;
wire x_37483;
wire x_37484;
wire x_37485;
wire x_37486;
wire x_37487;
wire x_37488;
wire x_37489;
wire x_37490;
wire x_37491;
wire x_37492;
wire x_37493;
wire x_37494;
wire x_37495;
wire x_37496;
wire x_37497;
wire x_37498;
wire x_37499;
wire x_37500;
wire x_37501;
wire x_37502;
wire x_37503;
wire x_37504;
wire x_37505;
wire x_37506;
wire x_37507;
wire x_37508;
wire x_37509;
wire x_37510;
wire x_37511;
wire x_37512;
wire x_37513;
wire x_37514;
wire x_37515;
wire x_37516;
wire x_37517;
wire x_37518;
wire x_37519;
wire x_37520;
wire x_37521;
wire x_37522;
wire x_37523;
wire x_37524;
wire x_37525;
wire x_37526;
wire x_37527;
wire x_37528;
wire x_37529;
wire x_37530;
wire x_37531;
wire x_37532;
wire x_37533;
wire x_37534;
wire x_37535;
wire x_37536;
wire x_37537;
wire x_37538;
wire x_37539;
wire x_37540;
wire x_37541;
wire x_37542;
wire x_37543;
wire x_37544;
wire x_37545;
wire x_37546;
wire x_37547;
wire x_37548;
wire x_37549;
wire x_37550;
wire x_37551;
wire x_37552;
wire x_37553;
wire x_37554;
wire x_37555;
wire x_37556;
wire x_37557;
wire x_37558;
wire x_37559;
wire x_37560;
wire x_37561;
wire x_37562;
wire x_37563;
wire x_37564;
wire x_37565;
wire x_37566;
wire x_37567;
wire x_37568;
wire x_37569;
wire x_37570;
wire x_37571;
wire x_37572;
wire x_37573;
wire x_37574;
wire x_37575;
wire x_37576;
wire x_37577;
wire x_37578;
wire x_37579;
wire x_37580;
wire x_37581;
wire x_37582;
wire x_37583;
wire x_37584;
wire x_37585;
wire x_37586;
wire x_37587;
wire x_37588;
wire x_37589;
wire x_37590;
wire x_37591;
wire x_37592;
wire x_37593;
wire x_37594;
wire x_37595;
wire x_37596;
wire x_37597;
wire x_37598;
wire x_37599;
wire x_37600;
wire x_37601;
wire x_37602;
wire x_37603;
wire x_37604;
wire x_37605;
wire x_37606;
wire x_37607;
wire x_37608;
wire x_37609;
wire x_37610;
wire x_37611;
wire x_37612;
wire x_37613;
wire x_37614;
wire x_37615;
wire x_37616;
wire x_37617;
wire x_37618;
wire x_37619;
wire x_37620;
wire x_37621;
wire x_37622;
wire x_37623;
wire x_37624;
wire x_37625;
wire x_37626;
wire x_37627;
wire x_37628;
wire x_37629;
wire x_37630;
wire x_37631;
wire x_37632;
wire x_37633;
wire x_37634;
wire x_37635;
wire x_37636;
wire x_37637;
wire x_37638;
wire x_37639;
wire x_37640;
wire x_37641;
wire x_37642;
wire x_37643;
wire x_37644;
wire x_37645;
wire x_37646;
wire x_37647;
wire x_37648;
wire x_37649;
wire x_37650;
wire x_37651;
wire x_37652;
wire x_37653;
wire x_37654;
wire x_37655;
wire x_37656;
wire x_37657;
wire x_37658;
wire x_37659;
wire x_37660;
wire x_37661;
wire x_37662;
wire x_37663;
wire x_37664;
wire x_37665;
wire x_37666;
wire x_37667;
wire x_37668;
wire x_37669;
wire x_37670;
wire x_37671;
wire x_37672;
wire x_37673;
wire x_37674;
wire x_37675;
wire x_37676;
wire x_37677;
wire x_37678;
wire x_37679;
wire x_37680;
wire x_37681;
wire x_37682;
wire x_37683;
wire x_37684;
wire x_37685;
wire x_37686;
wire x_37687;
wire x_37688;
wire x_37689;
wire x_37690;
wire x_37691;
wire x_37692;
wire x_37693;
wire x_37694;
wire x_37695;
wire x_37696;
wire x_37697;
wire x_37698;
wire x_37699;
wire x_37700;
wire x_37701;
wire x_37702;
wire x_37703;
wire x_37704;
wire x_37705;
wire x_37706;
wire x_37707;
wire x_37708;
wire x_37709;
wire x_37710;
wire x_37711;
wire x_37712;
wire x_37713;
wire x_37714;
wire x_37715;
wire x_37716;
wire x_37717;
wire x_37718;
wire x_37719;
wire x_37720;
wire x_37721;
wire x_37722;
wire x_37723;
wire x_37724;
wire x_37725;
wire x_37726;
wire x_37727;
wire x_37728;
wire x_37729;
wire x_37730;
wire x_37731;
wire x_37732;
wire x_37733;
wire x_37734;
wire x_37735;
wire x_37736;
wire x_37737;
wire x_37738;
wire x_37739;
wire x_37740;
wire x_37741;
wire x_37742;
wire x_37743;
wire x_37744;
wire x_37745;
wire x_37746;
wire x_37747;
wire x_37748;
wire x_37749;
wire x_37750;
wire x_37751;
wire x_37752;
wire x_37753;
wire x_37754;
wire x_37755;
wire x_37756;
wire x_37757;
wire x_37758;
wire x_37759;
wire x_37760;
wire x_37761;
wire x_37762;
wire x_37763;
wire x_37764;
wire x_37765;
wire x_37766;
wire x_37767;
wire x_37768;
wire x_37769;
wire x_37770;
wire x_37771;
wire x_37772;
wire x_37773;
wire x_37774;
wire x_37775;
wire x_37776;
wire x_37777;
wire x_37778;
wire x_37779;
wire x_37780;
wire x_37781;
wire x_37782;
wire x_37783;
wire x_37784;
wire x_37785;
wire x_37786;
wire x_37787;
wire x_37788;
wire x_37789;
wire x_37790;
wire x_37791;
wire x_37792;
wire x_37793;
wire x_37794;
wire x_37795;
wire x_37796;
wire x_37797;
wire x_37798;
wire x_37799;
wire x_37800;
wire x_37801;
wire x_37802;
wire x_37803;
wire x_37804;
wire x_37805;
wire x_37806;
wire x_37807;
wire x_37808;
wire x_37809;
wire x_37810;
wire x_37811;
wire x_37812;
wire x_37813;
wire x_37814;
wire x_37815;
wire x_37816;
wire x_37817;
wire x_37818;
wire x_37819;
wire x_37820;
wire x_37821;
wire x_37822;
wire x_37823;
wire x_37824;
wire x_37825;
wire x_37826;
wire x_37827;
wire x_37828;
wire x_37829;
wire x_37830;
wire x_37831;
wire x_37832;
wire x_37833;
wire x_37834;
wire x_37835;
wire x_37836;
wire x_37837;
wire x_37838;
wire x_37839;
wire x_37840;
wire x_37841;
wire x_37842;
wire x_37843;
wire x_37844;
wire x_37845;
wire x_37846;
wire x_37847;
wire x_37848;
wire x_37849;
wire x_37850;
wire x_37851;
wire x_37852;
wire x_37853;
wire x_37854;
wire x_37855;
wire x_37856;
wire x_37857;
wire x_37858;
wire x_37859;
wire x_37860;
wire x_37861;
wire x_37862;
wire x_37863;
wire x_37864;
wire x_37865;
wire x_37866;
wire x_37867;
wire x_37868;
wire x_37869;
wire x_37870;
wire x_37871;
wire x_37872;
wire x_37873;
wire x_37874;
wire x_37875;
wire x_37876;
wire x_37877;
wire x_37878;
wire x_37879;
wire x_37880;
wire x_37881;
wire x_37882;
wire x_37883;
wire x_37884;
wire x_37885;
wire x_37886;
wire x_37887;
wire x_37888;
wire x_37889;
wire x_37890;
wire x_37891;
wire x_37892;
wire x_37893;
wire x_37894;
wire x_37895;
wire x_37896;
wire x_37897;
wire x_37898;
wire x_37899;
wire x_37900;
wire x_37901;
wire x_37902;
wire x_37903;
wire x_37904;
wire x_37905;
wire x_37906;
wire x_37907;
wire x_37908;
wire x_37909;
wire x_37910;
wire x_37911;
wire x_37912;
wire x_37913;
wire x_37914;
wire x_37915;
wire x_37916;
wire x_37917;
wire x_37918;
wire x_37919;
wire x_37920;
wire x_37921;
wire x_37922;
wire x_37923;
wire x_37924;
wire x_37925;
wire x_37926;
wire x_37927;
wire x_37928;
wire x_37929;
wire x_37930;
wire x_37931;
wire x_37932;
wire x_37933;
wire x_37934;
wire x_37935;
wire x_37936;
wire x_37937;
wire x_37938;
wire x_37939;
wire x_37940;
wire x_37941;
wire x_37942;
wire x_37943;
wire x_37944;
wire x_37945;
wire x_37946;
wire x_37947;
wire x_37948;
wire x_37949;
wire x_37950;
wire x_37951;
wire x_37952;
wire x_37953;
wire x_37954;
wire x_37955;
wire x_37956;
wire x_37957;
wire x_37958;
wire x_37959;
wire x_37960;
wire x_37961;
wire x_37962;
wire x_37963;
wire x_37964;
wire x_37965;
wire x_37966;
wire x_37967;
wire x_37968;
wire x_37969;
wire x_37970;
wire x_37971;
wire x_37972;
wire x_37973;
wire x_37974;
wire x_37975;
wire x_37976;
wire x_37977;
wire x_37978;
wire x_37979;
wire x_37980;
wire x_37981;
wire x_37982;
wire x_37983;
wire x_37984;
wire x_37985;
wire x_37986;
wire x_37987;
wire x_37988;
wire x_37989;
wire x_37990;
wire x_37991;
wire x_37992;
wire x_37993;
wire x_37994;
wire x_37995;
wire x_37996;
wire x_37997;
wire x_37998;
wire x_37999;
wire x_38000;
wire x_38001;
wire x_38002;
wire x_38003;
wire x_38004;
wire x_38005;
wire x_38006;
wire x_38007;
wire x_38008;
wire x_38009;
wire x_38010;
wire x_38011;
wire x_38012;
wire x_38013;
wire x_38014;
wire x_38015;
wire x_38016;
wire x_38017;
wire x_38018;
wire x_38019;
wire x_38020;
wire x_38021;
wire x_38022;
wire x_38023;
wire x_38024;
wire x_38025;
wire x_38026;
wire x_38027;
wire x_38028;
wire x_38029;
wire x_38030;
wire x_38031;
wire x_38032;
wire x_38033;
wire x_38034;
wire x_38035;
wire x_38036;
wire x_38037;
wire x_38038;
wire x_38039;
wire x_38040;
wire x_38041;
wire x_38042;
wire x_38043;
wire x_38044;
wire x_38045;
wire x_38046;
wire x_38047;
wire x_38048;
wire x_38049;
wire x_38050;
wire x_38051;
wire x_38052;
wire x_38053;
wire x_38054;
wire x_38055;
wire x_38056;
wire x_38057;
wire x_38058;
wire x_38059;
wire x_38060;
wire x_38061;
wire x_38062;
wire x_38063;
wire x_38064;
wire x_38065;
wire x_38066;
wire x_38067;
wire x_38068;
wire x_38069;
wire x_38070;
wire x_38071;
wire x_38072;
wire x_38073;
wire x_38074;
wire x_38075;
wire x_38076;
wire x_38077;
wire x_38078;
wire x_38079;
wire x_38080;
wire x_38081;
wire x_38082;
wire x_38083;
wire x_38084;
wire x_38085;
wire x_38086;
wire x_38087;
wire x_38088;
wire x_38089;
wire x_38090;
wire x_38091;
wire x_38092;
wire x_38093;
wire x_38094;
wire x_38095;
wire x_38096;
wire x_38097;
wire x_38098;
wire x_38099;
wire x_38100;
wire x_38101;
wire x_38102;
wire x_38103;
wire x_38104;
wire x_38105;
wire x_38106;
wire x_38107;
wire x_38108;
wire x_38109;
wire x_38110;
wire x_38111;
wire x_38112;
wire x_38113;
wire x_38114;
wire x_38115;
wire x_38116;
wire x_38117;
wire x_38118;
wire x_38119;
wire x_38120;
wire x_38121;
wire x_38122;
wire x_38123;
wire x_38124;
wire x_38125;
wire x_38126;
wire x_38127;
wire x_38128;
wire x_38129;
wire x_38130;
wire x_38131;
wire x_38132;
wire x_38133;
wire x_38134;
wire x_38135;
wire x_38136;
wire x_38137;
wire x_38138;
wire x_38139;
wire x_38140;
wire x_38141;
wire x_38142;
wire x_38143;
wire x_38144;
wire x_38145;
wire x_38146;
wire x_38147;
wire x_38148;
wire x_38149;
wire x_38150;
wire x_38151;
wire x_38152;
wire x_38153;
wire x_38154;
wire x_38155;
wire x_38156;
wire x_38157;
wire x_38158;
wire x_38159;
wire x_38160;
wire x_38161;
wire x_38162;
wire x_38163;
wire x_38164;
wire x_38165;
wire x_38166;
wire x_38167;
wire x_38168;
wire x_38169;
wire x_38170;
wire x_38171;
wire x_38172;
wire x_38173;
wire x_38174;
wire x_38175;
wire x_38176;
wire x_38177;
wire x_38178;
wire x_38179;
wire x_38180;
wire x_38181;
wire x_38182;
wire x_38183;
wire x_38184;
wire x_38185;
wire x_38186;
wire x_38187;
wire x_38188;
wire x_38189;
wire x_38190;
wire x_38191;
wire x_38192;
wire x_38193;
wire x_38194;
wire x_38195;
wire x_38196;
wire x_38197;
wire x_38198;
wire x_38199;
wire x_38200;
wire x_38201;
wire x_38202;
wire x_38203;
wire x_38204;
wire x_38205;
wire x_38206;
wire x_38207;
wire x_38208;
wire x_38209;
wire x_38210;
wire x_38211;
wire x_38212;
wire x_38213;
wire x_38214;
wire x_38215;
wire x_38216;
wire x_38217;
wire x_38218;
wire x_38219;
wire x_38220;
wire x_38221;
wire x_38222;
wire x_38223;
wire x_38224;
wire x_38225;
wire x_38226;
wire x_38227;
wire x_38228;
wire x_38229;
wire x_38230;
wire x_38231;
wire x_38232;
wire x_38233;
wire x_38234;
wire x_38235;
wire x_38236;
wire x_38237;
wire x_38238;
wire x_38239;
wire x_38240;
wire x_38241;
wire x_38242;
wire x_38243;
wire x_38244;
wire x_38245;
wire x_38246;
wire x_38247;
wire x_38248;
wire x_38249;
wire x_38250;
wire x_38251;
wire x_38252;
wire x_38253;
wire x_38254;
wire x_38255;
wire x_38256;
wire x_38257;
wire x_38258;
wire x_38259;
wire x_38260;
wire x_38261;
wire x_38262;
wire x_38263;
wire x_38264;
wire x_38265;
wire x_38266;
wire x_38267;
wire x_38268;
wire x_38269;
wire x_38270;
wire x_38271;
wire x_38272;
wire x_38273;
wire x_38274;
wire x_38275;
wire x_38276;
wire x_38277;
wire x_38278;
wire x_38279;
wire x_38280;
wire x_38281;
wire x_38282;
wire x_38283;
wire x_38284;
wire x_38285;
wire x_38286;
wire x_38287;
wire x_38288;
wire x_38289;
wire x_38290;
wire x_38291;
wire x_38292;
wire x_38293;
wire x_38294;
wire x_38295;
wire x_38296;
wire x_38297;
wire x_38298;
wire x_38299;
wire x_38300;
wire x_38301;
wire x_38302;
wire x_38303;
wire x_38304;
wire x_38305;
wire x_38306;
wire x_38307;
wire x_38308;
wire x_38309;
wire x_38310;
wire x_38311;
wire x_38312;
wire x_38313;
wire x_38314;
wire x_38315;
wire x_38316;
wire x_38317;
wire x_38318;
wire x_38319;
wire x_38320;
wire x_38321;
wire x_38322;
wire x_38323;
wire x_38324;
wire x_38325;
wire x_38326;
wire x_38327;
wire x_38328;
wire x_38329;
wire x_38330;
wire x_38331;
wire x_38332;
wire x_38333;
wire x_38334;
wire x_38335;
wire x_38336;
wire x_38337;
wire x_38338;
wire x_38339;
wire x_38340;
wire x_38341;
wire x_38342;
wire x_38343;
wire x_38344;
wire x_38345;
wire x_38346;
wire x_38347;
wire x_38348;
wire x_38349;
wire x_38350;
wire x_38351;
wire x_38352;
wire x_38353;
wire x_38354;
wire x_38355;
wire x_38356;
wire x_38357;
wire x_38358;
wire x_38359;
wire x_38360;
wire x_38361;
wire x_38362;
wire x_38363;
wire x_38364;
wire x_38365;
wire x_38366;
wire x_38367;
wire x_38368;
wire x_38369;
wire x_38370;
wire x_38371;
wire x_38372;
wire x_38373;
wire x_38374;
wire x_38375;
wire x_38376;
wire x_38377;
wire x_38378;
wire x_38379;
wire x_38380;
wire x_38381;
wire x_38382;
wire x_38383;
wire x_38384;
wire x_38385;
wire x_38386;
wire x_38387;
wire x_38388;
wire x_38389;
wire x_38390;
wire x_38391;
wire x_38392;
wire x_38393;
wire x_38394;
wire x_38395;
wire x_38396;
wire x_38397;
wire x_38398;
wire x_38399;
wire x_38400;
wire x_38401;
wire x_38402;
wire x_38403;
wire x_38404;
wire x_38405;
wire x_38406;
wire x_38407;
wire x_38408;
wire x_38409;
wire x_38410;
wire x_38411;
wire x_38412;
wire x_38413;
wire x_38414;
wire x_38415;
wire x_38416;
wire x_38417;
wire x_38418;
wire x_38419;
wire x_38420;
wire x_38421;
wire x_38422;
wire x_38423;
wire x_38424;
wire x_38425;
wire x_38426;
wire x_38427;
wire x_38428;
wire x_38429;
wire x_38430;
wire x_38431;
wire x_38432;
wire x_38433;
wire x_38434;
wire x_38435;
wire x_38436;
wire x_38437;
wire x_38438;
wire x_38439;
wire x_38440;
wire x_38441;
wire x_38442;
wire x_38443;
wire x_38444;
wire x_38445;
wire x_38446;
wire x_38447;
wire x_38448;
wire x_38449;
wire x_38450;
wire x_38451;
wire x_38452;
wire x_38453;
wire x_38454;
wire x_38455;
wire x_38456;
wire x_38457;
wire x_38458;
wire x_38459;
wire x_38460;
wire x_38461;
wire x_38462;
wire x_38463;
wire x_38464;
wire x_38465;
wire x_38466;
wire x_38467;
wire x_38468;
wire x_38469;
wire x_38470;
wire x_38471;
wire x_38472;
wire x_38473;
wire x_38474;
wire x_38475;
wire x_38476;
wire x_38477;
wire x_38478;
wire x_38479;
wire x_38480;
wire x_38481;
wire x_38482;
wire x_38483;
wire x_38484;
wire x_38485;
wire x_38486;
wire x_38487;
wire x_38488;
wire x_38489;
wire x_38490;
wire x_38491;
wire x_38492;
wire x_38493;
wire x_38494;
wire x_38495;
wire x_38496;
wire x_38497;
wire x_38498;
wire x_38499;
wire x_38500;
wire x_38501;
wire x_38502;
wire x_38503;
wire x_38504;
wire x_38505;
wire x_38506;
wire x_38507;
wire x_38508;
wire x_38509;
wire x_38510;
wire x_38511;
wire x_38512;
wire x_38513;
wire x_38514;
wire x_38515;
wire x_38516;
wire x_38517;
wire x_38518;
wire x_38519;
wire x_38520;
wire x_38521;
wire x_38522;
wire x_38523;
wire x_38524;
wire x_38525;
wire x_38526;
wire x_38527;
wire x_38528;
wire x_38529;
wire x_38530;
wire x_38531;
wire x_38532;
wire x_38533;
wire x_38534;
wire x_38535;
wire x_38536;
wire x_38537;
wire x_38538;
wire x_38539;
wire x_38540;
wire x_38541;
wire x_38542;
wire x_38543;
wire x_38544;
wire x_38545;
wire x_38546;
wire x_38547;
wire x_38548;
wire x_38549;
wire x_38550;
wire x_38551;
wire x_38552;
wire x_38553;
wire x_38554;
wire x_38555;
wire x_38556;
wire x_38557;
wire x_38558;
wire x_38559;
wire x_38560;
wire x_38561;
wire x_38562;
wire x_38563;
wire x_38564;
wire x_38565;
wire x_38566;
wire x_38567;
wire x_38568;
wire x_38569;
wire x_38570;
wire x_38571;
wire x_38572;
wire x_38573;
wire x_38574;
wire x_38575;
wire x_38576;
wire x_38577;
wire x_38578;
wire x_38579;
wire x_38580;
wire x_38581;
wire x_38582;
wire x_38583;
wire x_38584;
wire x_38585;
wire x_38586;
wire x_38587;
wire x_38588;
wire x_38589;
wire x_38590;
wire x_38591;
wire x_38592;
wire x_38593;
wire x_38594;
wire x_38595;
wire x_38596;
wire x_38597;
wire x_38598;
wire x_38599;
wire x_38600;
wire x_38601;
wire x_38602;
wire x_38603;
wire x_38604;
wire x_38605;
wire x_38606;
wire x_38607;
wire x_38608;
wire x_38609;
wire x_38610;
wire x_38611;
wire x_38612;
wire x_38613;
wire x_38614;
wire x_38615;
wire x_38616;
wire x_38617;
wire x_38618;
wire x_38619;
wire x_38620;
wire x_38621;
wire x_38622;
wire x_38623;
wire x_38624;
wire x_38625;
wire x_38626;
wire x_38627;
wire x_38628;
wire x_38629;
wire x_38630;
wire x_38631;
wire x_38632;
wire x_38633;
wire x_38634;
wire x_38635;
wire x_38636;
wire x_38637;
wire x_38638;
wire x_38639;
wire x_38640;
wire x_38641;
wire x_38642;
wire x_38643;
wire x_38644;
wire x_38645;
wire x_38646;
wire x_38647;
wire x_38648;
wire x_38649;
wire x_38650;
wire x_38651;
wire x_38652;
wire x_38653;
wire x_38654;
wire x_38655;
wire x_38656;
wire x_38657;
wire x_38658;
wire x_38659;
wire x_38660;
wire x_38661;
wire x_38662;
wire x_38663;
wire x_38664;
wire x_38665;
wire x_38666;
wire x_38667;
wire x_38668;
wire x_38669;
wire x_38670;
wire x_38671;
wire x_38672;
wire x_38673;
wire x_38674;
wire x_38675;
wire x_38676;
wire x_38677;
wire x_38678;
wire x_38679;
wire x_38680;
wire x_38681;
wire x_38682;
wire x_38683;
wire x_38684;
wire x_38685;
wire x_38686;
wire x_38687;
wire x_38688;
wire x_38689;
wire x_38690;
wire x_38691;
wire x_38692;
wire x_38693;
wire x_38694;
wire x_38695;
wire x_38696;
wire x_38697;
wire x_38698;
wire x_38699;
wire x_38700;
wire x_38701;
wire x_38702;
wire x_38703;
wire x_38704;
wire x_38705;
wire x_38706;
wire x_38707;
wire x_38708;
wire x_38709;
wire x_38710;
wire x_38711;
wire x_38712;
wire x_38713;
wire x_38714;
wire x_38715;
wire x_38716;
wire x_38717;
wire x_38718;
wire x_38719;
wire x_38720;
wire x_38721;
wire x_38722;
wire x_38723;
wire x_38724;
wire x_38725;
wire x_38726;
wire x_38727;
wire x_38728;
wire x_38729;
wire x_38730;
wire x_38731;
wire x_38732;
wire x_38733;
wire x_38734;
wire x_38735;
wire x_38736;
wire x_38737;
wire x_38738;
wire x_38739;
wire x_38740;
wire x_38741;
wire x_38742;
wire x_38743;
wire x_38744;
wire x_38745;
wire x_38746;
wire x_38747;
wire x_38748;
wire x_38749;
wire x_38750;
wire x_38751;
wire x_38752;
wire x_38753;
wire x_38754;
wire x_38755;
wire x_38756;
wire x_38757;
wire x_38758;
wire x_38759;
wire x_38760;
wire x_38761;
wire x_38762;
wire x_38763;
wire x_38764;
wire x_38765;
wire x_38766;
wire x_38767;
wire x_38768;
wire x_38769;
wire x_38770;
wire x_38771;
wire x_38772;
wire x_38773;
wire x_38774;
wire x_38775;
wire x_38776;
wire x_38777;
wire x_38778;
wire x_38779;
wire x_38780;
wire x_38781;
wire x_38782;
wire x_38783;
wire x_38784;
wire x_38785;
wire x_38786;
wire x_38787;
wire x_38788;
wire x_38789;
wire x_38790;
wire x_38791;
wire x_38792;
wire x_38793;
wire x_38794;
wire x_38795;
wire x_38796;
wire x_38797;
wire x_38798;
wire x_38799;
wire x_38800;
wire x_38801;
wire x_38802;
wire x_38803;
wire x_38804;
wire x_38805;
wire x_38806;
wire x_38807;
wire x_38808;
wire x_38809;
wire x_38810;
wire x_38811;
wire x_38812;
wire x_38813;
wire x_38814;
wire x_38815;
wire x_38816;
wire x_38817;
wire x_38818;
wire x_38819;
wire x_38820;
wire x_38821;
wire x_38822;
wire x_38823;
wire x_38824;
wire x_38825;
wire x_38826;
wire x_38827;
wire x_38828;
wire x_38829;
wire x_38830;
wire x_38831;
wire x_38832;
wire x_38833;
wire x_38834;
wire x_38835;
wire x_38836;
wire x_38837;
wire x_38838;
wire x_38839;
wire x_38840;
wire x_38841;
wire x_38842;
wire x_38843;
wire x_38844;
wire x_38845;
wire x_38846;
wire x_38847;
wire x_38848;
wire x_38849;
wire x_38850;
wire x_38851;
wire x_38852;
wire x_38853;
wire x_38854;
wire x_38855;
wire x_38856;
wire x_38857;
wire x_38858;
wire x_38859;
wire x_38860;
wire x_38861;
wire x_38862;
wire x_38863;
wire x_38864;
wire x_38865;
wire x_38866;
wire x_38867;
wire x_38868;
wire x_38869;
wire x_38870;
wire x_38871;
wire x_38872;
wire x_38873;
wire x_38874;
wire x_38875;
wire x_38876;
wire x_38877;
wire x_38878;
wire x_38879;
wire x_38880;
wire x_38881;
wire x_38882;
wire x_38883;
wire x_38884;
wire x_38885;
wire x_38886;
wire x_38887;
wire x_38888;
wire x_38889;
wire x_38890;
wire x_38891;
wire x_38892;
wire x_38893;
wire x_38894;
wire x_38895;
wire x_38896;
wire x_38897;
wire x_38898;
wire x_38899;
wire x_38900;
wire x_38901;
wire x_38902;
wire x_38903;
wire x_38904;
wire x_38905;
wire x_38906;
wire x_38907;
wire x_38908;
wire x_38909;
wire x_38910;
wire x_38911;
wire x_38912;
wire x_38913;
wire x_38914;
wire x_38915;
wire x_38916;
wire x_38917;
wire x_38918;
wire x_38919;
wire x_38920;
wire x_38921;
wire x_38922;
wire x_38923;
wire x_38924;
wire x_38925;
wire x_38926;
wire x_38927;
wire x_38928;
wire x_38929;
wire x_38930;
wire x_38931;
wire x_38932;
wire x_38933;
wire x_38934;
wire x_38935;
wire x_38936;
wire x_38937;
wire x_38938;
wire x_38939;
wire x_38940;
wire x_38941;
wire x_38942;
wire x_38943;
wire x_38944;
wire x_38945;
wire x_38946;
wire x_38947;
wire x_38948;
wire x_38949;
wire x_38950;
wire x_38951;
wire x_38952;
wire x_38953;
wire x_38954;
wire x_38955;
wire x_38956;
wire x_38957;
wire x_38958;
wire x_38959;
wire x_38960;
wire x_38961;
wire x_38962;
wire x_38963;
wire x_38964;
wire x_38965;
wire x_38966;
wire x_38967;
wire x_38968;
wire x_38969;
wire x_38970;
wire x_38971;
wire x_38972;
wire x_38973;
wire x_38974;
wire x_38975;
wire x_38976;
wire x_38977;
wire x_38978;
wire x_38979;
wire x_38980;
wire x_38981;
wire x_38982;
wire x_38983;
wire x_38984;
wire x_38985;
wire x_38986;
wire x_38987;
wire x_38988;
wire x_38989;
wire x_38990;
wire x_38991;
wire x_38992;
wire x_38993;
wire x_38994;
wire x_38995;
wire x_38996;
wire x_38997;
wire x_38998;
wire x_38999;
wire x_39000;
wire x_39001;
wire x_39002;
wire x_39003;
wire x_39004;
wire x_39005;
wire x_39006;
wire x_39007;
wire x_39008;
wire x_39009;
wire x_39010;
wire x_39011;
wire x_39012;
wire x_39013;
wire x_39014;
wire x_39015;
wire x_39016;
wire x_39017;
wire x_39018;
wire x_39019;
wire x_39020;
wire x_39021;
wire x_39022;
wire x_39023;
wire x_39024;
wire x_39025;
wire x_39026;
wire x_39027;
wire x_39028;
wire x_39029;
wire x_39030;
wire x_39031;
wire x_39032;
wire x_39033;
wire x_39034;
wire x_39035;
wire x_39036;
wire x_39037;
wire x_39038;
wire x_39039;
wire x_39040;
wire x_39041;
wire x_39042;
wire x_39043;
wire x_39044;
wire x_39045;
wire x_39046;
wire x_39047;
wire x_39048;
wire x_39049;
wire x_39050;
wire x_39051;
wire x_39052;
wire x_39053;
wire x_39054;
wire x_39055;
wire x_39056;
wire x_39057;
wire x_39058;
wire x_39059;
wire x_39060;
wire x_39061;
wire x_39062;
wire x_39063;
wire x_39064;
wire x_39065;
wire x_39066;
wire x_39067;
wire x_39068;
wire x_39069;
wire x_39070;
wire x_39071;
wire x_39072;
wire x_39073;
wire x_39074;
wire x_39075;
wire x_39076;
wire x_39077;
wire x_39078;
wire x_39079;
wire x_39080;
wire x_39081;
wire x_39082;
wire x_39083;
wire x_39084;
wire x_39085;
wire x_39086;
wire x_39087;
wire x_39088;
wire x_39089;
wire x_39090;
wire x_39091;
wire x_39092;
wire x_39093;
wire x_39094;
wire x_39095;
wire x_39096;
wire x_39097;
wire x_39098;
wire x_39099;
wire x_39100;
wire x_39101;
wire x_39102;
wire x_39103;
wire x_39104;
wire x_39105;
wire x_39106;
wire x_39107;
wire x_39108;
wire x_39109;
wire x_39110;
wire x_39111;
wire x_39112;
wire x_39113;
wire x_39114;
wire x_39115;
wire x_39116;
wire x_39117;
wire x_39118;
wire x_39119;
wire x_39120;
wire x_39121;
wire x_39122;
wire x_39123;
wire x_39124;
wire x_39125;
wire x_39126;
wire x_39127;
wire x_39128;
wire x_39129;
wire x_39130;
wire x_39131;
wire x_39132;
wire x_39133;
wire x_39134;
wire x_39135;
wire x_39136;
wire x_39137;
wire x_39138;
wire x_39139;
wire x_39140;
wire x_39141;
wire x_39142;
wire x_39143;
wire x_39144;
wire x_39145;
wire x_39146;
wire x_39147;
wire x_39148;
wire x_39149;
wire x_39150;
wire x_39151;
wire x_39152;
wire x_39153;
wire x_39154;
wire x_39155;
wire x_39156;
wire x_39157;
wire x_39158;
wire x_39159;
wire x_39160;
wire x_39161;
wire x_39162;
wire x_39163;
wire x_39164;
wire x_39165;
wire x_39166;
wire x_39167;
wire x_39168;
wire x_39169;
wire x_39170;
wire x_39171;
wire x_39172;
wire x_39173;
wire x_39174;
wire x_39175;
wire x_39176;
wire x_39177;
wire x_39178;
wire x_39179;
wire x_39180;
wire x_39181;
wire x_39182;
wire x_39183;
wire x_39184;
wire x_39185;
wire x_39186;
wire x_39187;
wire x_39188;
wire x_39189;
wire x_39190;
wire x_39191;
wire x_39192;
wire x_39193;
wire x_39194;
wire x_39195;
wire x_39196;
wire x_39197;
wire x_39198;
wire x_39199;
wire x_39200;
wire x_39201;
wire x_39202;
wire x_39203;
wire x_39204;
wire x_39205;
wire x_39206;
wire x_39207;
wire x_39208;
wire x_39209;
wire x_39210;
wire x_39211;
wire x_39212;
wire x_39213;
wire x_39214;
wire x_39215;
wire x_39216;
wire x_39217;
wire x_39218;
wire x_39219;
wire x_39220;
wire x_39221;
wire x_39222;
wire x_39223;
wire x_39224;
wire x_39225;
wire x_39226;
wire x_39227;
wire x_39228;
wire x_39229;
wire x_39230;
wire x_39231;
wire x_39232;
wire x_39233;
wire x_39234;
wire x_39235;
wire x_39236;
wire x_39237;
wire x_39238;
wire x_39239;
wire x_39240;
wire x_39241;
wire x_39242;
wire x_39243;
wire x_39244;
wire x_39245;
wire x_39246;
wire x_39247;
wire x_39248;
wire x_39249;
wire x_39250;
wire x_39251;
wire x_39252;
wire x_39253;
wire x_39254;
wire x_39255;
wire x_39256;
wire x_39257;
wire x_39258;
wire x_39259;
wire x_39260;
wire x_39261;
wire x_39262;
wire x_39263;
wire x_39264;
wire x_39265;
wire x_39266;
wire x_39267;
wire x_39268;
wire x_39269;
wire x_39270;
wire x_39271;
wire x_39272;
wire x_39273;
wire x_39274;
wire x_39275;
wire x_39276;
wire x_39277;
wire x_39278;
wire x_39279;
wire x_39280;
wire x_39281;
wire x_39282;
wire x_39283;
wire x_39284;
wire x_39285;
wire x_39286;
wire x_39287;
wire x_39288;
wire x_39289;
wire x_39290;
wire x_39291;
wire x_39292;
wire x_39293;
wire x_39294;
wire x_39295;
wire x_39296;
wire x_39297;
wire x_39298;
wire x_39299;
wire x_39300;
wire x_39301;
wire x_39302;
wire x_39303;
wire x_39304;
wire x_39305;
wire x_39306;
wire x_39307;
wire x_39308;
wire x_39309;
wire x_39310;
wire x_39311;
wire x_39312;
wire x_39313;
wire x_39314;
wire x_39315;
wire x_39316;
wire x_39317;
wire x_39318;
wire x_39319;
wire x_39320;
wire x_39321;
wire x_39322;
wire x_39323;
wire x_39324;
wire x_39325;
wire x_39326;
wire x_39327;
wire x_39328;
wire x_39329;
wire x_39330;
wire x_39331;
wire x_39332;
wire x_39333;
wire x_39334;
wire x_39335;
wire x_39336;
wire x_39337;
wire x_39338;
wire x_39339;
wire x_39340;
wire x_39341;
wire x_39342;
wire x_39343;
wire x_39344;
wire x_39345;
wire x_39346;
wire x_39347;
wire x_39348;
wire x_39349;
wire x_39350;
wire x_39351;
wire x_39352;
wire x_39353;
wire x_39354;
wire x_39355;
wire x_39356;
wire x_39357;
wire x_39358;
wire x_39359;
wire x_39360;
wire x_39361;
wire x_39362;
wire x_39363;
wire x_39364;
wire x_39365;
wire x_39366;
wire x_39367;
wire x_39368;
wire x_39369;
wire x_39370;
wire x_39371;
wire x_39372;
wire x_39373;
wire x_39374;
wire x_39375;
wire x_39376;
wire x_39377;
wire x_39378;
wire x_39379;
wire x_39380;
wire x_39381;
wire x_39382;
wire x_39383;
wire x_39384;
wire x_39385;
wire x_39386;
wire x_39387;
wire x_39388;
wire x_39389;
wire x_39390;
wire x_39391;
wire x_39392;
wire x_39393;
wire x_39394;
wire x_39395;
wire x_39396;
wire x_39397;
wire x_39398;
wire x_39399;
wire x_39400;
wire x_39401;
wire x_39402;
wire x_39403;
wire x_39404;
wire x_39405;
wire x_39406;
wire x_39407;
wire x_39408;
wire x_39409;
wire x_39410;
wire x_39411;
wire x_39412;
wire x_39413;
wire x_39414;
wire x_39415;
wire x_39416;
wire x_39417;
wire x_39418;
wire x_39419;
wire x_39420;
wire x_39421;
wire x_39422;
wire x_39423;
wire x_39424;
wire x_39425;
wire x_39426;
wire x_39427;
wire x_39428;
wire x_39429;
wire x_39430;
wire x_39431;
wire x_39432;
wire x_39433;
wire x_39434;
wire x_39435;
wire x_39436;
wire x_39437;
wire x_39438;
wire x_39439;
wire x_39440;
wire x_39441;
wire x_39442;
wire x_39443;
wire x_39444;
wire x_39445;
wire x_39446;
wire x_39447;
wire x_39448;
wire x_39449;
wire x_39450;
wire x_39451;
wire x_39452;
wire x_39453;
wire x_39454;
wire x_39455;
wire x_39456;
wire x_39457;
wire x_39458;
wire x_39459;
wire x_39460;
wire x_39461;
wire x_39462;
wire x_39463;
wire x_39464;
wire x_39465;
wire x_39466;
wire x_39467;
wire x_39468;
wire x_39469;
wire x_39470;
wire x_39471;
wire x_39472;
wire x_39473;
wire x_39474;
wire x_39475;
wire x_39476;
wire x_39477;
wire x_39478;
wire x_39479;
wire x_39480;
wire x_39481;
wire x_39482;
wire x_39483;
wire x_39484;
wire x_39485;
wire x_39486;
wire x_39487;
wire x_39488;
wire x_39489;
wire x_39490;
wire x_39491;
wire x_39492;
wire x_39493;
wire x_39494;
wire x_39495;
wire x_39496;
wire x_39497;
wire x_39498;
wire x_39499;
wire x_39500;
wire x_39501;
wire x_39502;
wire x_39503;
wire x_39504;
wire x_39505;
wire x_39506;
wire x_39507;
wire x_39508;
wire x_39509;
wire x_39510;
wire x_39511;
wire x_39512;
wire x_39513;
wire x_39514;
wire x_39515;
wire x_39516;
wire x_39517;
wire x_39518;
wire x_39519;
wire x_39520;
wire x_39521;
wire x_39522;
wire x_39523;
wire x_39524;
wire x_39525;
wire x_39526;
wire x_39527;
wire x_39528;
wire x_39529;
wire x_39530;
wire x_39531;
wire x_39532;
wire x_39533;
wire x_39534;
wire x_39535;
wire x_39536;
wire x_39537;
wire x_39538;
wire x_39539;
wire x_39540;
wire x_39541;
wire x_39542;
wire x_39543;
wire x_39544;
wire x_39545;
wire x_39546;
wire x_39547;
wire x_39548;
wire x_39549;
wire x_39550;
wire x_39551;
wire x_39552;
wire x_39553;
wire x_39554;
wire x_39555;
wire x_39556;
wire x_39557;
wire x_39558;
wire x_39559;
wire x_39560;
wire x_39561;
wire x_39562;
wire x_39563;
wire x_39564;
wire x_39565;
wire x_39566;
wire x_39567;
wire x_39568;
wire x_39569;
wire x_39570;
wire x_39571;
wire x_39572;
wire x_39573;
wire x_39574;
wire x_39575;
wire x_39576;
wire x_39577;
wire x_39578;
wire x_39579;
wire x_39580;
wire x_39581;
wire x_39582;
wire x_39583;
wire x_39584;
wire x_39585;
wire x_39586;
wire x_39587;
wire x_39588;
wire x_39589;
wire x_39590;
wire x_39591;
wire x_39592;
wire x_39593;
wire x_39594;
wire x_39595;
wire x_39596;
wire x_39597;
wire x_39598;
wire x_39599;
wire x_39600;
wire x_39601;
wire x_39602;
wire x_39603;
wire x_39604;
wire x_39605;
wire x_39606;
wire x_39607;
wire x_39608;
wire x_39609;
wire x_39610;
wire x_39611;
wire x_39612;
wire x_39613;
wire x_39614;
wire x_39615;
wire x_39616;
wire x_39617;
wire x_39618;
wire x_39619;
wire x_39620;
wire x_39621;
wire x_39622;
wire x_39623;
wire x_39624;
wire x_39625;
wire x_39626;
wire x_39627;
wire x_39628;
wire x_39629;
wire x_39630;
wire x_39631;
wire x_39632;
wire x_39633;
wire x_39634;
wire x_39635;
wire x_39636;
wire x_39637;
wire x_39638;
wire x_39639;
wire x_39640;
wire x_39641;
wire x_39642;
wire x_39643;
wire x_39644;
wire x_39645;
wire x_39646;
wire x_39647;
wire x_39648;
wire x_39649;
wire x_39650;
wire x_39651;
wire x_39652;
wire x_39653;
wire x_39654;
wire x_39655;
wire x_39656;
wire x_39657;
wire x_39658;
wire x_39659;
wire x_39660;
wire x_39661;
wire x_39662;
wire x_39663;
wire x_39664;
wire x_39665;
wire x_39666;
wire x_39667;
wire x_39668;
wire x_39669;
wire x_39670;
wire x_39671;
wire x_39672;
wire x_39673;
wire x_39674;
wire x_39675;
wire x_39676;
wire x_39677;
wire x_39678;
wire x_39679;
wire x_39680;
wire x_39681;
wire x_39682;
wire x_39683;
wire x_39684;
wire x_39685;
wire x_39686;
wire x_39687;
wire x_39688;
wire x_39689;
wire x_39690;
wire x_39691;
wire x_39692;
wire x_39693;
wire x_39694;
wire x_39695;
wire x_39696;
wire x_39697;
wire x_39698;
wire x_39699;
wire x_39700;
wire x_39701;
wire x_39702;
wire x_39703;
wire x_39704;
wire x_39705;
wire x_39706;
wire x_39707;
wire x_39708;
wire x_39709;
wire x_39710;
wire x_39711;
wire x_39712;
wire x_39713;
wire x_39714;
wire x_39715;
wire x_39716;
wire x_39717;
wire x_39718;
wire x_39719;
wire x_39720;
wire x_39721;
wire x_39722;
wire x_39723;
wire x_39724;
wire x_39725;
wire x_39726;
wire x_39727;
wire x_39728;
wire x_39729;
wire x_39730;
wire x_39731;
wire x_39732;
wire x_39733;
wire x_39734;
wire x_39735;
wire x_39736;
wire x_39737;
wire x_39738;
wire x_39739;
wire x_39740;
wire x_39741;
wire x_39742;
wire x_39743;
wire x_39744;
wire x_39745;
wire x_39746;
wire x_39747;
wire x_39748;
wire x_39749;
wire x_39750;
wire x_39751;
wire x_39752;
wire x_39753;
wire x_39754;
wire x_39755;
wire x_39756;
wire x_39757;
wire x_39758;
wire x_39759;
wire x_39760;
wire x_39761;
wire x_39762;
wire x_39763;
wire x_39764;
wire x_39765;
wire x_39766;
wire x_39767;
wire x_39768;
wire x_39769;
wire x_39770;
wire x_39771;
wire x_39772;
wire x_39773;
wire x_39774;
wire x_39775;
wire x_39776;
wire x_39777;
wire x_39778;
wire x_39779;
wire x_39780;
wire x_39781;
wire x_39782;
wire x_39783;
wire x_39784;
wire x_39785;
wire x_39786;
wire x_39787;
wire x_39788;
wire x_39789;
wire x_39790;
wire x_39791;
wire x_39792;
wire x_39793;
wire x_39794;
wire x_39795;
wire x_39796;
wire x_39797;
wire x_39798;
wire x_39799;
wire x_39800;
wire x_39801;
wire x_39802;
wire x_39803;
wire x_39804;
wire x_39805;
wire x_39806;
wire x_39807;
wire x_39808;
wire x_39809;
wire x_39810;
wire x_39811;
wire x_39812;
wire x_39813;
wire x_39814;
wire x_39815;
wire x_39816;
wire x_39817;
wire x_39818;
wire x_39819;
wire x_39820;
wire x_39821;
wire x_39822;
wire x_39823;
wire x_39824;
wire x_39825;
wire x_39826;
wire x_39827;
wire x_39828;
wire x_39829;
wire x_39830;
wire x_39831;
wire x_39832;
wire x_39833;
wire x_39834;
wire x_39835;
wire x_39836;
wire x_39837;
wire x_39838;
wire x_39839;
wire x_39840;
wire x_39841;
wire x_39842;
wire x_39843;
wire x_39844;
wire x_39845;
wire x_39846;
wire x_39847;
wire x_39848;
wire x_39849;
wire x_39850;
wire x_39851;
wire x_39852;
wire x_39853;
wire x_39854;
wire x_39855;
wire x_39856;
wire x_39857;
wire x_39858;
wire x_39859;
wire x_39860;
wire x_39861;
wire x_39862;
wire x_39863;
wire x_39864;
wire x_39865;
wire x_39866;
wire x_39867;
wire x_39868;
wire x_39869;
wire x_39870;
wire x_39871;
wire x_39872;
wire x_39873;
wire x_39874;
wire x_39875;
wire x_39876;
wire x_39877;
wire x_39878;
wire x_39879;
wire x_39880;
wire x_39881;
wire x_39882;
wire x_39883;
wire x_39884;
wire x_39885;
wire x_39886;
wire x_39887;
wire x_39888;
wire x_39889;
wire x_39890;
wire x_39891;
wire x_39892;
wire x_39893;
wire x_39894;
wire x_39895;
wire x_39896;
wire x_39897;
wire x_39898;
wire x_39899;
wire x_39900;
wire x_39901;
wire x_39902;
wire x_39903;
wire x_39904;
wire x_39905;
wire x_39906;
wire x_39907;
wire x_39908;
wire x_39909;
wire x_39910;
wire x_39911;
wire x_39912;
wire x_39913;
wire x_39914;
wire x_39915;
wire x_39916;
wire x_39917;
wire x_39918;
wire x_39919;
wire x_39920;
wire x_39921;
wire x_39922;
wire x_39923;
wire x_39924;
wire x_39925;
wire x_39926;
wire x_39927;
wire x_39928;
wire x_39929;
wire x_39930;
wire x_39931;
wire x_39932;
wire x_39933;
wire x_39934;
wire x_39935;
wire x_39936;
wire x_39937;
wire x_39938;
wire x_39939;
wire x_39940;
wire x_39941;
wire x_39942;
wire x_39943;
wire x_39944;
wire x_39945;
wire x_39946;
wire x_39947;
wire x_39948;
wire x_39949;
wire x_39950;
wire x_39951;
wire x_39952;
wire x_39953;
wire x_39954;
wire x_39955;
wire x_39956;
wire x_39957;
wire x_39958;
wire x_39959;
wire x_39960;
wire x_39961;
wire x_39962;
wire x_39963;
wire x_39964;
wire x_39965;
wire x_39966;
wire x_39967;
wire x_39968;
wire x_39969;
wire x_39970;
wire x_39971;
wire x_39972;
wire x_39973;
wire x_39974;
wire x_39975;
wire x_39976;
wire x_39977;
wire x_39978;
wire x_39979;
wire x_39980;
wire x_39981;
wire x_39982;
wire x_39983;
wire x_39984;
wire x_39985;
wire x_39986;
wire x_39987;
wire x_39988;
wire x_39989;
wire x_39990;
wire x_39991;
wire x_39992;
wire x_39993;
wire x_39994;
wire x_39995;
wire x_39996;
wire x_39997;
wire x_39998;
wire x_39999;
wire x_40000;
wire x_40001;
wire x_40002;
wire x_40003;
wire x_40004;
wire x_40005;
wire x_40006;
wire x_40007;
wire x_40008;
wire x_40009;
wire x_40010;
wire x_40011;
wire x_40012;
wire x_40013;
wire x_40014;
wire x_40015;
wire x_40016;
wire x_40017;
wire x_40018;
wire x_40019;
wire x_40020;
wire x_40021;
wire x_40022;
wire x_40023;
wire x_40024;
wire x_40025;
wire x_40026;
wire x_40027;
wire x_40028;
wire x_40029;
wire x_40030;
wire x_40031;
wire x_40032;
wire x_40033;
wire x_40034;
wire x_40035;
wire x_40036;
wire x_40037;
wire x_40038;
wire x_40039;
wire x_40040;
wire x_40041;
wire x_40042;
wire x_40043;
wire x_40044;
wire x_40045;
wire x_40046;
wire x_40047;
wire x_40048;
wire x_40049;
wire x_40050;
wire x_40051;
wire x_40052;
wire x_40053;
wire x_40054;
wire x_40055;
wire x_40056;
wire x_40057;
wire x_40058;
wire x_40059;
wire x_40060;
wire x_40061;
wire x_40062;
wire x_40063;
wire x_40064;
wire x_40065;
wire x_40066;
wire x_40067;
wire x_40068;
wire x_40069;
wire x_40070;
wire x_40071;
wire x_40072;
wire x_40073;
wire x_40074;
wire x_40075;
wire x_40076;
wire x_40077;
wire x_40078;
wire x_40079;
wire x_40080;
wire x_40081;
wire x_40082;
wire x_40083;
wire x_40084;
wire x_40085;
wire x_40086;
wire x_40087;
wire x_40088;
wire x_40089;
wire x_40090;
wire x_40091;
wire x_40092;
wire x_40093;
wire x_40094;
wire x_40095;
wire x_40096;
wire x_40097;
wire x_40098;
wire x_40099;
wire x_40100;
wire x_40101;
wire x_40102;
wire x_40103;
wire x_40104;
wire x_40105;
wire x_40106;
wire x_40107;
wire x_40108;
wire x_40109;
wire x_40110;
wire x_40111;
wire x_40112;
wire x_40113;
wire x_40114;
wire x_40115;
wire x_40116;
wire x_40117;
wire x_40118;
wire x_40119;
wire x_40120;
wire x_40121;
wire x_40122;
wire x_40123;
wire x_40124;
wire x_40125;
wire x_40126;
wire x_40127;
wire x_40128;
wire x_40129;
wire x_40130;
wire x_40131;
wire x_40132;
wire x_40133;
wire x_40134;
wire x_40135;
wire x_40136;
wire x_40137;
wire x_40138;
wire x_40139;
wire x_40140;
wire x_40141;
wire x_40142;
wire x_40143;
wire x_40144;
wire x_40145;
wire x_40146;
wire x_40147;
wire x_40148;
wire x_40149;
wire x_40150;
wire x_40151;
wire x_40152;
wire x_40153;
wire x_40154;
wire x_40155;
wire x_40156;
wire x_40157;
wire x_40158;
wire x_40159;
wire x_40160;
wire x_40161;
wire x_40162;
wire x_40163;
wire x_40164;
wire x_40165;
wire x_40166;
wire x_40167;
wire x_40168;
wire x_40169;
wire x_40170;
wire x_40171;
wire x_40172;
wire x_40173;
wire x_40174;
wire x_40175;
wire x_40176;
wire x_40177;
wire x_40178;
wire x_40179;
wire x_40180;
wire x_40181;
wire x_40182;
wire x_40183;
wire x_40184;
wire x_40185;
wire x_40186;
wire x_40187;
wire x_40188;
wire x_40189;
wire x_40190;
wire x_40191;
wire x_40192;
wire x_40193;
wire x_40194;
wire x_40195;
wire x_40196;
wire x_40197;
wire x_40198;
wire x_40199;
wire x_40200;
wire x_40201;
wire x_40202;
wire x_40203;
wire x_40204;
wire x_40205;
wire x_40206;
wire x_40207;
wire x_40208;
wire x_40209;
wire x_40210;
wire x_40211;
wire x_40212;
wire x_40213;
wire x_40214;
wire x_40215;
wire x_40216;
wire x_40217;
wire x_40218;
wire x_40219;
wire x_40220;
wire x_40221;
wire x_40222;
wire x_40223;
wire x_40224;
wire x_40225;
wire x_40226;
wire x_40227;
wire x_40228;
wire x_40229;
wire x_40230;
wire x_40231;
wire x_40232;
wire x_40233;
wire x_40234;
wire x_40235;
wire x_40236;
wire x_40237;
wire x_40238;
wire x_40239;
wire x_40240;
wire x_40241;
wire x_40242;
wire x_40243;
wire x_40244;
wire x_40245;
wire x_40246;
wire x_40247;
wire x_40248;
wire x_40249;
wire x_40250;
wire x_40251;
wire x_40252;
wire x_40253;
wire x_40254;
wire x_40255;
wire x_40256;
wire x_40257;
wire x_40258;
wire x_40259;
wire x_40260;
wire x_40261;
wire x_40262;
wire x_40263;
wire x_40264;
wire x_40265;
wire x_40266;
wire x_40267;
wire x_40268;
wire x_40269;
wire x_40270;
wire x_40271;
wire x_40272;
wire x_40273;
wire x_40274;
wire x_40275;
wire x_40276;
wire x_40277;
wire x_40278;
wire x_40279;
wire x_40280;
wire x_40281;
wire x_40282;
wire x_40283;
wire x_40284;
wire x_40285;
wire x_40286;
wire x_40287;
wire x_40288;
wire x_40289;
wire x_40290;
wire x_40291;
wire x_40292;
wire x_40293;
wire x_40294;
wire x_40295;
wire x_40296;
wire x_40297;
wire x_40298;
wire x_40299;
wire x_40300;
wire x_40301;
wire x_40302;
wire x_40303;
wire x_40304;
wire x_40305;
wire x_40306;
wire x_40307;
wire x_40308;
wire x_40309;
wire x_40310;
wire x_40311;
wire x_40312;
wire x_40313;
wire x_40314;
wire x_40315;
wire x_40316;
wire x_40317;
wire x_40318;
wire x_40319;
wire x_40320;
wire x_40321;
wire x_40322;
wire x_40323;
wire x_40324;
wire x_40325;
wire x_40326;
wire x_40327;
wire x_40328;
wire x_40329;
wire x_40330;
wire x_40331;
wire x_40332;
wire x_40333;
wire x_40334;
wire x_40335;
wire x_40336;
wire x_40337;
wire x_40338;
wire x_40339;
wire x_40340;
wire x_40341;
wire x_40342;
wire x_40343;
wire x_40344;
wire x_40345;
wire x_40346;
wire x_40347;
wire x_40348;
wire x_40349;
wire x_40350;
wire x_40351;
wire x_40352;
wire x_40353;
wire x_40354;
wire x_40355;
wire x_40356;
wire x_40357;
wire x_40358;
wire x_40359;
wire x_40360;
wire x_40361;
wire x_40362;
wire x_40363;
wire x_40364;
wire x_40365;
wire x_40366;
wire x_40367;
wire x_40368;
wire x_40369;
wire x_40370;
wire x_40371;
wire x_40372;
wire x_40373;
wire x_40374;
wire x_40375;
wire x_40376;
wire x_40377;
wire x_40378;
wire x_40379;
wire x_40380;
wire x_40381;
wire x_40382;
wire x_40383;
wire x_40384;
wire x_40385;
wire x_40386;
wire x_40387;
wire x_40388;
wire x_40389;
wire x_40390;
wire x_40391;
wire x_40392;
wire x_40393;
wire x_40394;
wire x_40395;
wire x_40396;
wire x_40397;
wire x_40398;
wire x_40399;
wire x_40400;
wire x_40401;
wire x_40402;
wire x_40403;
wire x_40404;
wire x_40405;
wire x_40406;
wire x_40407;
wire x_40408;
wire x_40409;
wire x_40410;
wire x_40411;
wire x_40412;
wire x_40413;
wire x_40414;
wire x_40415;
wire x_40416;
wire x_40417;
wire x_40418;
wire x_40419;
wire x_40420;
wire x_40421;
wire x_40422;
wire x_40423;
wire x_40424;
wire x_40425;
wire x_40426;
wire x_40427;
wire x_40428;
wire x_40429;
wire x_40430;
wire x_40431;
wire x_40432;
wire x_40433;
wire x_40434;
wire x_40435;
wire x_40436;
wire x_40437;
wire x_40438;
wire x_40439;
wire x_40440;
wire x_40441;
wire x_40442;
wire x_40443;
wire x_40444;
wire x_40445;
wire x_40446;
wire x_40447;
wire x_40448;
wire x_40449;
wire x_40450;
wire x_40451;
wire x_40452;
wire x_40453;
wire x_40454;
wire x_40455;
wire x_40456;
wire x_40457;
wire x_40458;
wire x_40459;
wire x_40460;
wire x_40461;
wire x_40462;
wire x_40463;
wire x_40464;
wire x_40465;
wire x_40466;
wire x_40467;
wire x_40468;
wire x_40469;
wire x_40470;
wire x_40471;
wire x_40472;
wire x_40473;
wire x_40474;
wire x_40475;
wire x_40476;
wire x_40477;
wire x_40478;
wire x_40479;
wire x_40480;
wire x_40481;
wire x_40482;
wire x_40483;
wire x_40484;
wire x_40485;
wire x_40486;
wire x_40487;
wire x_40488;
wire x_40489;
wire x_40490;
wire x_40491;
wire x_40492;
wire x_40493;
wire x_40494;
wire x_40495;
wire x_40496;
wire x_40497;
wire x_40498;
wire x_40499;
wire x_40500;
wire x_40501;
wire x_40502;
wire x_40503;
wire x_40504;
wire x_40505;
wire x_40506;
wire x_40507;
wire x_40508;
wire x_40509;
wire x_40510;
wire x_40511;
wire x_40512;
wire x_40513;
wire x_40514;
wire x_40515;
wire x_40516;
wire x_40517;
wire x_40518;
wire x_40519;
wire x_40520;
wire x_40521;
wire x_40522;
wire x_40523;
wire x_40524;
wire x_40525;
wire x_40526;
wire x_40527;
wire x_40528;
wire x_40529;
wire x_40530;
wire x_40531;
wire x_40532;
wire x_40533;
wire x_40534;
wire x_40535;
wire x_40536;
wire x_40537;
wire x_40538;
wire x_40539;
wire x_40540;
wire x_40541;
wire x_40542;
wire x_40543;
wire x_40544;
wire x_40545;
wire x_40546;
wire x_40547;
wire x_40548;
wire x_40549;
wire x_40550;
wire x_40551;
wire x_40552;
wire x_40553;
wire x_40554;
wire x_40555;
wire x_40556;
wire x_40557;
wire x_40558;
wire x_40559;
wire x_40560;
wire x_40561;
wire x_40562;
wire x_40563;
wire x_40564;
wire x_40565;
wire x_40566;
wire x_40567;
wire x_40568;
wire x_40569;
wire x_40570;
wire x_40571;
wire x_40572;
wire x_40573;
wire x_40574;
wire x_40575;
wire x_40576;
wire x_40577;
wire x_40578;
wire x_40579;
wire x_40580;
wire x_40581;
wire x_40582;
wire x_40583;
wire x_40584;
wire x_40585;
wire x_40586;
wire x_40587;
wire x_40588;
wire x_40589;
wire x_40590;
wire x_40591;
wire x_40592;
wire x_40593;
wire x_40594;
wire x_40595;
wire x_40596;
wire x_40597;
wire x_40598;
wire x_40599;
wire x_40600;
wire x_40601;
wire x_40602;
wire x_40603;
wire x_40604;
wire x_40605;
wire x_40606;
wire x_40607;
wire x_40608;
wire x_40609;
wire x_40610;
wire x_40611;
wire x_40612;
wire x_40613;
wire x_40614;
wire x_40615;
wire x_40616;
wire x_40617;
wire x_40618;
wire x_40619;
wire x_40620;
wire x_40621;
wire x_40622;
wire x_40623;
wire x_40624;
wire x_40625;
wire x_40626;
wire x_40627;
wire x_40628;
wire x_40629;
wire x_40630;
wire x_40631;
wire x_40632;
wire x_40633;
wire x_40634;
wire x_40635;
wire x_40636;
wire x_40637;
wire x_40638;
wire x_40639;
wire x_40640;
wire x_40641;
wire x_40642;
wire x_40643;
wire x_40644;
wire x_40645;
wire x_40646;
wire x_40647;
wire x_40648;
wire x_40649;
wire x_40650;
wire x_40651;
wire x_40652;
wire x_40653;
wire x_40654;
wire x_40655;
wire x_40656;
wire x_40657;
wire x_40658;
wire x_40659;
wire x_40660;
wire x_40661;
wire x_40662;
wire x_40663;
wire x_40664;
wire x_40665;
wire x_40666;
wire x_40667;
wire x_40668;
wire x_40669;
wire x_40670;
wire x_40671;
wire x_40672;
wire x_40673;
wire x_40674;
wire x_40675;
wire x_40676;
wire x_40677;
wire x_40678;
wire x_40679;
wire x_40680;
wire x_40681;
wire x_40682;
wire x_40683;
wire x_40684;
wire x_40685;
wire x_40686;
wire x_40687;
wire x_40688;
wire x_40689;
wire x_40690;
wire x_40691;
wire x_40692;
wire x_40693;
wire x_40694;
wire x_40695;
wire x_40696;
wire x_40697;
wire x_40698;
wire x_40699;
wire x_40700;
wire x_40701;
wire x_40702;
wire x_40703;
wire x_40704;
wire x_40705;
wire x_40706;
wire x_40707;
wire x_40708;
wire x_40709;
wire x_40710;
wire x_40711;
wire x_40712;
wire x_40713;
wire x_40714;
wire x_40715;
wire x_40716;
wire x_40717;
wire x_40718;
wire x_40719;
wire x_40720;
wire x_40721;
wire x_40722;
wire x_40723;
wire x_40724;
wire x_40725;
wire x_40726;
wire x_40727;
wire x_40728;
wire x_40729;
wire x_40730;
wire x_40731;
wire x_40732;
wire x_40733;
wire x_40734;
wire x_40735;
wire x_40736;
wire x_40737;
wire x_40738;
wire x_40739;
wire x_40740;
wire x_40741;
wire x_40742;
wire x_40743;
wire x_40744;
wire x_40745;
wire x_40746;
wire x_40747;
wire x_40748;
wire x_40749;
wire x_40750;
wire x_40751;
wire x_40752;
wire x_40753;
wire x_40754;
wire x_40755;
wire x_40756;
wire x_40757;
wire x_40758;
wire x_40759;
wire x_40760;
wire x_40761;
wire x_40762;
wire x_40763;
wire x_40764;
wire x_40765;
wire x_40766;
wire x_40767;
wire x_40768;
wire x_40769;
wire x_40770;
wire x_40771;
wire x_40772;
wire x_40773;
wire x_40774;
wire x_40775;
wire x_40776;
wire x_40777;
wire x_40778;
wire x_40779;
wire x_40780;
wire x_40781;
wire x_40782;
wire x_40783;
wire x_40784;
wire x_40785;
wire x_40786;
wire x_40787;
wire x_40788;
wire x_40789;
wire x_40790;
wire x_40791;
wire x_40792;
wire x_40793;
wire x_40794;
wire x_40795;
wire x_40796;
wire x_40797;
wire x_40798;
wire x_40799;
wire x_40800;
wire x_40801;
wire x_40802;
wire x_40803;
wire x_40804;
wire x_40805;
wire x_40806;
wire x_40807;
wire x_40808;
wire x_40809;
wire x_40810;
wire x_40811;
wire x_40812;
wire x_40813;
wire x_40814;
wire x_40815;
wire x_40816;
wire x_40817;
wire x_40818;
wire x_40819;
wire x_40820;
wire x_40821;
wire x_40822;
wire x_40823;
wire x_40824;
wire x_40825;
wire x_40826;
wire x_40827;
wire x_40828;
wire x_40829;
wire x_40830;
wire x_40831;
wire x_40832;
wire x_40833;
wire x_40834;
wire x_40835;
wire x_40836;
wire x_40837;
wire x_40838;
wire x_40839;
wire x_40840;
wire x_40841;
wire x_40842;
wire x_40843;
wire x_40844;
wire x_40845;
wire x_40846;
wire x_40847;
wire x_40848;
wire x_40849;
wire x_40850;
wire x_40851;
wire x_40852;
wire x_40853;
wire x_40854;
wire x_40855;
wire x_40856;
wire x_40857;
wire x_40858;
wire x_40859;
wire x_40860;
wire x_40861;
wire x_40862;
wire x_40863;
wire x_40864;
wire x_40865;
wire x_40866;
wire x_40867;
wire x_40868;
wire x_40869;
wire x_40870;
wire x_40871;
wire x_40872;
wire x_40873;
wire x_40874;
wire x_40875;
wire x_40876;
wire x_40877;
wire x_40878;
wire x_40879;
wire x_40880;
wire x_40881;
wire x_40882;
wire x_40883;
wire x_40884;
wire x_40885;
wire x_40886;
wire x_40887;
wire x_40888;
wire x_40889;
wire x_40890;
wire x_40891;
wire x_40892;
wire x_40893;
wire x_40894;
wire x_40895;
wire x_40896;
wire x_40897;
wire x_40898;
wire x_40899;
wire x_40900;
wire x_40901;
wire x_40902;
wire x_40903;
wire x_40904;
wire x_40905;
wire x_40906;
wire x_40907;
wire x_40908;
wire x_40909;
wire x_40910;
wire x_40911;
wire x_40912;
wire x_40913;
wire x_40914;
wire x_40915;
wire x_40916;
wire x_40917;
wire x_40918;
wire x_40919;
wire x_40920;
wire x_40921;
wire x_40922;
wire x_40923;
wire x_40924;
wire x_40925;
wire x_40926;
wire x_40927;
wire x_40928;
wire x_40929;
wire x_40930;
wire x_40931;
wire x_40932;
wire x_40933;
wire x_40934;
wire x_40935;
wire x_40936;
wire x_40937;
wire x_40938;
wire x_40939;
wire x_40940;
wire x_40941;
wire x_40942;
wire x_40943;
wire x_40944;
wire x_40945;
wire x_40946;
wire x_40947;
wire x_40948;
wire x_40949;
wire x_40950;
wire x_40951;
wire x_40952;
wire x_40953;
wire x_40954;
wire x_40955;
wire x_40956;
wire x_40957;
wire x_40958;
wire x_40959;
wire x_40960;
wire x_40961;
wire x_40962;
wire x_40963;
wire x_40964;
wire x_40965;
wire x_40966;
wire x_40967;
wire x_40968;
wire x_40969;
wire x_40970;
wire x_40971;
wire x_40972;
wire x_40973;
wire x_40974;
wire x_40975;
wire x_40976;
wire x_40977;
wire x_40978;
wire x_40979;
wire x_40980;
wire x_40981;
wire x_40982;
wire x_40983;
wire x_40984;
wire x_40985;
wire x_40986;
wire x_40987;
wire x_40988;
wire x_40989;
wire x_40990;
wire x_40991;
wire x_40992;
wire x_40993;
wire x_40994;
wire x_40995;
wire x_40996;
wire x_40997;
wire x_40998;
wire x_40999;
wire x_41000;
wire x_41001;
wire x_41002;
wire x_41003;
wire x_41004;
wire x_41005;
wire x_41006;
wire x_41007;
wire x_41008;
wire x_41009;
wire x_41010;
wire x_41011;
wire x_41012;
wire x_41013;
wire x_41014;
wire x_41015;
wire x_41016;
wire x_41017;
wire x_41018;
wire x_41019;
wire x_41020;
wire x_41021;
wire x_41022;
wire x_41023;
wire x_41024;
wire x_41025;
wire x_41026;
wire x_41027;
wire x_41028;
wire x_41029;
wire x_41030;
wire x_41031;
wire x_41032;
wire x_41033;
wire x_41034;
wire x_41035;
wire x_41036;
wire x_41037;
wire x_41038;
wire x_41039;
wire x_41040;
wire x_41041;
wire x_41042;
wire x_41043;
wire x_41044;
wire x_41045;
wire x_41046;
wire x_41047;
wire x_41048;
wire x_41049;
wire x_41050;
wire x_41051;
wire x_41052;
wire x_41053;
wire x_41054;
wire x_41055;
wire x_41056;
wire x_41057;
wire x_41058;
wire x_41059;
wire x_41060;
wire x_41061;
wire x_41062;
wire x_41063;
wire x_41064;
wire x_41065;
wire x_41066;
wire x_41067;
wire x_41068;
wire x_41069;
wire x_41070;
wire x_41071;
wire x_41072;
wire x_41073;
wire x_41074;
wire x_41075;
wire x_41076;
wire x_41077;
wire x_41078;
wire x_41079;
wire x_41080;
wire x_41081;
wire x_41082;
wire x_41083;
wire x_41084;
wire x_41085;
wire x_41086;
wire x_41087;
wire x_41088;
wire x_41089;
wire x_41090;
wire x_41091;
wire x_41092;
wire x_41093;
wire x_41094;
wire x_41095;
wire x_41096;
wire x_41097;
wire x_41098;
wire x_41099;
wire x_41100;
wire x_41101;
wire x_41102;
wire x_41103;
wire x_41104;
wire x_41105;
wire x_41106;
wire x_41107;
wire x_41108;
wire x_41109;
wire x_41110;
wire x_41111;
wire x_41112;
wire x_41113;
wire x_41114;
wire x_41115;
wire x_41116;
wire x_41117;
wire x_41118;
wire x_41119;
wire x_41120;
wire x_41121;
wire x_41122;
wire x_41123;
wire x_41124;
wire x_41125;
wire x_41126;
wire x_41127;
wire x_41128;
wire x_41129;
wire x_41130;
wire x_41131;
wire x_41132;
wire x_41133;
wire x_41134;
wire x_41135;
wire x_41136;
wire x_41137;
wire x_41138;
wire x_41139;
wire x_41140;
wire x_41141;
wire x_41142;
wire x_41143;
wire x_41144;
wire x_41145;
wire x_41146;
wire x_41147;
wire x_41148;
wire x_41149;
wire x_41150;
wire x_41151;
wire x_41152;
wire x_41153;
wire x_41154;
wire x_41155;
wire x_41156;
wire x_41157;
wire x_41158;
wire x_41159;
wire x_41160;
wire x_41161;
wire x_41162;
wire x_41163;
wire x_41164;
wire x_41165;
wire x_41166;
wire x_41167;
wire x_41168;
wire x_41169;
wire x_41170;
wire x_41171;
wire x_41172;
wire x_41173;
wire x_41174;
wire x_41175;
wire x_41176;
wire x_41177;
wire x_41178;
wire x_41179;
wire x_41180;
wire x_41181;
wire x_41182;
wire x_41183;
wire x_41184;
wire x_41185;
wire x_41186;
wire x_41187;
wire x_41188;
wire x_41189;
wire x_41190;
wire x_41191;
wire x_41192;
wire x_41193;
wire x_41194;
wire x_41195;
wire x_41196;
wire x_41197;
wire x_41198;
wire x_41199;
wire x_41200;
wire x_41201;
wire x_41202;
wire x_41203;
wire x_41204;
wire x_41205;
wire x_41206;
wire x_41207;
wire x_41208;
wire x_41209;
wire x_41210;
wire x_41211;
wire x_41212;
wire x_41213;
wire x_41214;
wire x_41215;
wire x_41216;
wire x_41217;
wire x_41218;
wire x_41219;
wire x_41220;
wire x_41221;
wire x_41222;
wire x_41223;
wire x_41224;
wire x_41225;
wire x_41226;
wire x_41227;
wire x_41228;
wire x_41229;
wire x_41230;
wire x_41231;
wire x_41232;
wire x_41233;
wire x_41234;
wire x_41235;
wire x_41236;
wire x_41237;
wire x_41238;
wire x_41239;
wire x_41240;
wire x_41241;
wire x_41242;
wire x_41243;
wire x_41244;
wire x_41245;
wire x_41246;
wire x_41247;
wire x_41248;
wire x_41249;
wire x_41250;
wire x_41251;
wire x_41252;
wire x_41253;
wire x_41254;
wire x_41255;
wire x_41256;
wire x_41257;
wire x_41258;
wire x_41259;
wire x_41260;
wire x_41261;
wire x_41262;
wire x_41263;
wire x_41264;
wire x_41265;
wire x_41266;
wire x_41267;
wire x_41268;
wire x_41269;
wire x_41270;
wire x_41271;
wire x_41272;
wire x_41273;
wire x_41274;
wire x_41275;
wire x_41276;
wire x_41277;
wire x_41278;
wire x_41279;
wire x_41280;
wire x_41281;
wire x_41282;
wire x_41283;
wire x_41284;
wire x_41285;
wire x_41286;
wire x_41287;
wire x_41288;
wire x_41289;
wire x_41290;
wire x_41291;
wire x_41292;
wire x_41293;
wire x_41294;
wire x_41295;
wire x_41296;
wire x_41297;
wire x_41298;
wire x_41299;
wire x_41300;
wire x_41301;
wire x_41302;
wire x_41303;
wire x_41304;
wire x_41305;
wire x_41306;
wire x_41307;
wire x_41308;
wire x_41309;
wire x_41310;
wire x_41311;
wire x_41312;
wire x_41313;
wire x_41314;
wire x_41315;
wire x_41316;
wire x_41317;
wire x_41318;
wire x_41319;
wire x_41320;
wire x_41321;
wire x_41322;
wire x_41323;
wire x_41324;
wire x_41325;
wire x_41326;
wire x_41327;
wire x_41328;
wire x_41329;
wire x_41330;
wire x_41331;
wire x_41332;
wire x_41333;
wire x_41334;
wire x_41335;
wire x_41336;
wire x_41337;
wire x_41338;
wire x_41339;
wire x_41340;
wire x_41341;
wire x_41342;
wire x_41343;
wire x_41344;
wire x_41345;
wire x_41346;
wire x_41347;
wire x_41348;
wire x_41349;
wire x_41350;
wire x_41351;
wire x_41352;
wire x_41353;
wire x_41354;
wire x_41355;
wire x_41356;
wire x_41357;
wire x_41358;
wire x_41359;
wire x_41360;
wire x_41361;
wire x_41362;
wire x_41363;
wire x_41364;
wire x_41365;
wire x_41366;
wire x_41367;
wire x_41368;
wire x_41369;
wire x_41370;
wire x_41371;
wire x_41372;
wire x_41373;
wire x_41374;
wire x_41375;
wire x_41376;
wire x_41377;
wire x_41378;
wire x_41379;
wire x_41380;
wire x_41381;
wire x_41382;
wire x_41383;
wire x_41384;
wire x_41385;
wire x_41386;
wire x_41387;
wire x_41388;
wire x_41389;
wire x_41390;
wire x_41391;
wire x_41392;
wire x_41393;
wire x_41394;
wire x_41395;
wire x_41396;
wire x_41397;
wire x_41398;
wire x_41399;
wire x_41400;
wire x_41401;
wire x_41402;
wire x_41403;
wire x_41404;
wire x_41405;
wire x_41406;
wire x_41407;
wire x_41408;
wire x_41409;
wire x_41410;
wire x_41411;
wire x_41412;
wire x_41413;
wire x_41414;
wire x_41415;
wire x_41416;
wire x_41417;
wire x_41418;
wire x_41419;
wire x_41420;
wire x_41421;
wire x_41422;
wire x_41423;
wire x_41424;
wire x_41425;
wire x_41426;
wire x_41427;
wire x_41428;
wire x_41429;
wire x_41430;
wire x_41431;
wire x_41432;
wire x_41433;
wire x_41434;
wire x_41435;
wire x_41436;
wire x_41437;
wire x_41438;
wire x_41439;
wire x_41440;
wire x_41441;
wire x_41442;
wire x_41443;
wire x_41444;
wire x_41445;
wire x_41446;
wire x_41447;
wire x_41448;
wire x_41449;
wire x_41450;
wire x_41451;
wire x_41452;
wire x_41453;
wire x_41454;
wire x_41455;
wire x_41456;
wire x_41457;
wire x_41458;
wire x_41459;
wire x_41460;
wire x_41461;
wire x_41462;
wire x_41463;
wire x_41464;
wire x_41465;
wire x_41466;
wire x_41467;
wire x_41468;
wire x_41469;
wire x_41470;
wire x_41471;
wire x_41472;
wire x_41473;
wire x_41474;
wire x_41475;
wire x_41476;
wire x_41477;
wire x_41478;
wire x_41479;
wire x_41480;
wire x_41481;
wire x_41482;
wire x_41483;
wire x_41484;
wire x_41485;
wire x_41486;
wire x_41487;
wire x_41488;
wire x_41489;
wire x_41490;
wire x_41491;
wire x_41492;
wire x_41493;
wire x_41494;
wire x_41495;
wire x_41496;
wire x_41497;
wire x_41498;
wire x_41499;
wire x_41500;
wire x_41501;
wire x_41502;
wire x_41503;
wire x_41504;
wire x_41505;
wire x_41506;
wire x_41507;
wire x_41508;
wire x_41509;
wire x_41510;
wire x_41511;
wire x_41512;
wire x_41513;
wire x_41514;
wire x_41515;
wire x_41516;
wire x_41517;
wire x_41518;
wire x_41519;
wire x_41520;
wire x_41521;
wire x_41522;
wire x_41523;
wire x_41524;
wire x_41525;
wire x_41526;
wire x_41527;
wire x_41528;
wire x_41529;
wire x_41530;
wire x_41531;
wire x_41532;
wire x_41533;
wire x_41534;
wire x_41535;
wire x_41536;
wire x_41537;
wire x_41538;
wire x_41539;
wire x_41540;
wire x_41541;
wire x_41542;
wire x_41543;
wire x_41544;
wire x_41545;
wire x_41546;
wire x_41547;
wire x_41548;
wire x_41549;
wire x_41550;
wire x_41551;
wire x_41552;
wire x_41553;
wire x_41554;
wire x_41555;
wire x_41556;
wire x_41557;
wire x_41558;
wire x_41559;
wire x_41560;
wire x_41561;
wire x_41562;
wire x_41563;
wire x_41564;
wire x_41565;
wire x_41566;
wire x_41567;
wire x_41568;
wire x_41569;
wire x_41570;
wire x_41571;
wire x_41572;
wire x_41573;
wire x_41574;
wire x_41575;
wire x_41576;
wire x_41577;
wire x_41578;
wire x_41579;
wire x_41580;
wire x_41581;
wire x_41582;
wire x_41583;
wire x_41584;
wire x_41585;
wire x_41586;
wire x_41587;
wire x_41588;
wire x_41589;
wire x_41590;
wire x_41591;
wire x_41592;
wire x_41593;
wire x_41594;
wire x_41595;
wire x_41596;
wire x_41597;
wire x_41598;
wire x_41599;
wire x_41600;
wire x_41601;
wire x_41602;
wire x_41603;
wire x_41604;
wire x_41605;
wire x_41606;
wire x_41607;
wire x_41608;
wire x_41609;
wire x_41610;
wire x_41611;
wire x_41612;
wire x_41613;
wire x_41614;
wire x_41615;
wire x_41616;
wire x_41617;
wire x_41618;
wire x_41619;
wire x_41620;
wire x_41621;
wire x_41622;
wire x_41623;
wire x_41624;
wire x_41625;
wire x_41626;
wire x_41627;
wire x_41628;
wire x_41629;
wire x_41630;
wire x_41631;
wire x_41632;
wire x_41633;
wire x_41634;
wire x_41635;
wire x_41636;
wire x_41637;
wire x_41638;
wire x_41639;
wire x_41640;
wire x_41641;
wire x_41642;
wire x_41643;
wire x_41644;
wire x_41645;
wire x_41646;
wire x_41647;
wire x_41648;
wire x_41649;
wire x_41650;
wire x_41651;
wire x_41652;
wire x_41653;
wire x_41654;
wire x_41655;
wire x_41656;
wire x_41657;
wire x_41658;
wire x_41659;
wire x_41660;
wire x_41661;
wire x_41662;
wire x_41663;
wire x_41664;
wire x_41665;
wire x_41666;
wire x_41667;
wire x_41668;
wire x_41669;
wire x_41670;
wire x_41671;
wire x_41672;
wire x_41673;
wire x_41674;
wire x_41675;
wire x_41676;
wire x_41677;
wire x_41678;
wire x_41679;
wire x_41680;
wire x_41681;
wire x_41682;
wire x_41683;
wire x_41684;
wire x_41685;
wire x_41686;
wire x_41687;
wire x_41688;
wire x_41689;
wire x_41690;
wire x_41691;
wire x_41692;
wire x_41693;
wire x_41694;
wire x_41695;
wire x_41696;
wire x_41697;
wire x_41698;
wire x_41699;
wire x_41700;
wire x_41701;
wire x_41702;
wire x_41703;
wire x_41704;
wire x_41705;
wire x_41706;
wire x_41707;
wire x_41708;
wire x_41709;
wire x_41710;
wire x_41711;
wire x_41712;
wire x_41713;
wire x_41714;
wire x_41715;
wire x_41716;
wire x_41717;
wire x_41718;
wire x_41719;
wire x_41720;
wire x_41721;
wire x_41722;
wire x_41723;
wire x_41724;
wire x_41725;
wire x_41726;
wire x_41727;
wire x_41728;
wire x_41729;
wire x_41730;
wire x_41731;
wire x_41732;
wire x_41733;
wire x_41734;
wire x_41735;
wire x_41736;
wire x_41737;
wire x_41738;
wire x_41739;
wire x_41740;
wire x_41741;
wire x_41742;
wire x_41743;
wire x_41744;
wire x_41745;
wire x_41746;
wire x_41747;
wire x_41748;
wire x_41749;
wire x_41750;
wire x_41751;
wire x_41752;
wire x_41753;
wire x_41754;
wire x_41755;
wire x_41756;
wire x_41757;
wire x_41758;
wire x_41759;
wire x_41760;
wire x_41761;
wire x_41762;
wire x_41763;
wire x_41764;
wire x_41765;
wire x_41766;
wire x_41767;
wire x_41768;
wire x_41769;
wire x_41770;
wire x_41771;
wire x_41772;
wire x_41773;
wire x_41774;
wire x_41775;
wire x_41776;
wire x_41777;
wire x_41778;
wire x_41779;
wire x_41780;
wire x_41781;
wire x_41782;
wire x_41783;
wire x_41784;
wire x_41785;
wire x_41786;
wire x_41787;
wire x_41788;
wire x_41789;
wire x_41790;
wire x_41791;
wire x_41792;
wire x_41793;
wire x_41794;
wire x_41795;
wire x_41796;
wire x_41797;
wire x_41798;
wire x_41799;
wire x_41800;
wire x_41801;
wire x_41802;
wire x_41803;
wire x_41804;
wire x_41805;
wire x_41806;
wire x_41807;
wire x_41808;
wire x_41809;
wire x_41810;
wire x_41811;
wire x_41812;
wire x_41813;
wire x_41814;
wire x_41815;
wire x_41816;
wire x_41817;
wire x_41818;
wire x_41819;
wire x_41820;
wire x_41821;
wire x_41822;
wire x_41823;
wire x_41824;
wire x_41825;
wire x_41826;
wire x_41827;
wire x_41828;
wire x_41829;
wire x_41830;
wire x_41831;
wire x_41832;
wire x_41833;
wire x_41834;
wire x_41835;
wire x_41836;
wire x_41837;
wire x_41838;
wire x_41839;
wire x_41840;
wire x_41841;
wire x_41842;
wire x_41843;
wire x_41844;
wire x_41845;
wire x_41846;
wire x_41847;
wire x_41848;
wire x_41849;
wire x_41850;
wire x_41851;
wire x_41852;
wire x_41853;
wire x_41854;
wire x_41855;
wire x_41856;
wire x_41857;
wire x_41858;
wire x_41859;
wire x_41860;
wire x_41861;
wire x_41862;
wire x_41863;
wire x_41864;
wire x_41865;
wire x_41866;
wire x_41867;
wire x_41868;
wire x_41869;
wire x_41870;
wire x_41871;
wire x_41872;
wire x_41873;
wire x_41874;
wire x_41875;
wire x_41876;
wire x_41877;
wire x_41878;
wire x_41879;
wire x_41880;
wire x_41881;
wire x_41882;
wire x_41883;
wire x_41884;
wire x_41885;
wire x_41886;
wire x_41887;
wire x_41888;
wire x_41889;
wire x_41890;
wire x_41891;
wire x_41892;
wire x_41893;
wire x_41894;
wire x_41895;
wire x_41896;
wire x_41897;
wire x_41898;
wire x_41899;
wire x_41900;
wire x_41901;
wire x_41902;
wire x_41903;
wire x_41904;
wire x_41905;
wire x_41906;
wire x_41907;
wire x_41908;
wire x_41909;
wire x_41910;
wire x_41911;
wire x_41912;
wire x_41913;
wire x_41914;
wire x_41915;
wire x_41916;
wire x_41917;
wire x_41918;
wire x_41919;
wire x_41920;
wire x_41921;
wire x_41922;
wire x_41923;
wire x_41924;
wire x_41925;
wire x_41926;
wire x_41927;
wire x_41928;
wire x_41929;
wire x_41930;
wire x_41931;
wire x_41932;
wire x_41933;
wire x_41934;
wire x_41935;
wire x_41936;
wire x_41937;
wire x_41938;
wire x_41939;
wire x_41940;
wire x_41941;
wire x_41942;
wire x_41943;
wire x_41944;
wire x_41945;
wire x_41946;
wire x_41947;
wire x_41948;
wire x_41949;
wire x_41950;
wire x_41951;
wire x_41952;
wire x_41953;
wire x_41954;
wire x_41955;
wire x_41956;
wire x_41957;
wire x_41958;
wire x_41959;
wire x_41960;
wire x_41961;
wire x_41962;
wire x_41963;
wire x_41964;
wire x_41965;
wire x_41966;
wire x_41967;
wire x_41968;
wire x_41969;
wire x_41970;
wire x_41971;
wire x_41972;
wire x_41973;
wire x_41974;
wire x_41975;
wire x_41976;
wire x_41977;
wire x_41978;
wire x_41979;
wire x_41980;
wire x_41981;
wire x_41982;
wire x_41983;
wire x_41984;
wire x_41985;
wire x_41986;
wire x_41987;
wire x_41988;
wire x_41989;
wire x_41990;
wire x_41991;
wire x_41992;
wire x_41993;
wire x_41994;
wire x_41995;
wire x_41996;
wire x_41997;
wire x_41998;
wire x_41999;
wire x_42000;
wire x_42001;
wire x_42002;
wire x_42003;
wire x_42004;
wire x_42005;
wire x_42006;
wire x_42007;
wire x_42008;
wire x_42009;
wire x_42010;
wire x_42011;
wire x_42012;
wire x_42013;
wire x_42014;
wire x_42015;
wire x_42016;
wire x_42017;
wire x_42018;
wire x_42019;
wire x_42020;
wire x_42021;
wire x_42022;
wire x_42023;
wire x_42024;
wire x_42025;
wire x_42026;
wire x_42027;
wire x_42028;
wire x_42029;
wire x_42030;
wire x_42031;
wire x_42032;
wire x_42033;
wire x_42034;
wire x_42035;
wire x_42036;
wire x_42037;
wire x_42038;
wire x_42039;
wire x_42040;
wire x_42041;
wire x_42042;
wire x_42043;
wire x_42044;
wire x_42045;
wire x_42046;
wire x_42047;
wire x_42048;
wire x_42049;
wire x_42050;
wire x_42051;
wire x_42052;
wire x_42053;
wire x_42054;
wire x_42055;
wire x_42056;
wire x_42057;
wire x_42058;
wire x_42059;
wire x_42060;
wire x_42061;
wire x_42062;
wire x_42063;
wire x_42064;
wire x_42065;
wire x_42066;
wire x_42067;
wire x_42068;
wire x_42069;
wire x_42070;
wire x_42071;
wire x_42072;
wire x_42073;
wire x_42074;
wire x_42075;
wire x_42076;
wire x_42077;
wire x_42078;
wire x_42079;
wire x_42080;
wire x_42081;
wire x_42082;
wire x_42083;
wire x_42084;
wire x_42085;
wire x_42086;
wire x_42087;
wire x_42088;
wire x_42089;
wire x_42090;
wire x_42091;
wire x_42092;
wire x_42093;
wire x_42094;
wire x_42095;
wire x_42096;
wire x_42097;
wire x_42098;
wire x_42099;
wire x_42100;
wire x_42101;
wire x_42102;
wire x_42103;
wire x_42104;
wire x_42105;
wire x_42106;
wire x_42107;
wire x_42108;
wire x_42109;
wire x_42110;
wire x_42111;
wire x_42112;
wire x_42113;
wire x_42114;
wire x_42115;
wire x_42116;
wire x_42117;
wire x_42118;
wire x_42119;
wire x_42120;
wire x_42121;
wire x_42122;
wire x_42123;
wire x_42124;
wire x_42125;
wire x_42126;
wire x_42127;
wire x_42128;
wire x_42129;
wire x_42130;
wire x_42131;
wire x_42132;
wire x_42133;
wire x_42134;
wire x_42135;
wire x_42136;
wire x_42137;
wire x_42138;
wire x_42139;
wire x_42140;
wire x_42141;
wire x_42142;
wire x_42143;
wire x_42144;
wire x_42145;
wire x_42146;
wire x_42147;
wire x_42148;
wire x_42149;
wire x_42150;
wire x_42151;
wire x_42152;
wire x_42153;
wire x_42154;
wire x_42155;
wire x_42156;
wire x_42157;
wire x_42158;
wire x_42159;
wire x_42160;
wire x_42161;
wire x_42162;
wire x_42163;
wire x_42164;
wire x_42165;
wire x_42166;
wire x_42167;
wire x_42168;
wire x_42169;
wire x_42170;
wire x_42171;
wire x_42172;
wire x_42173;
wire x_42174;
wire x_42175;
wire x_42176;
wire x_42177;
wire x_42178;
wire x_42179;
wire x_42180;
wire x_42181;
wire x_42182;
wire x_42183;
wire x_42184;
wire x_42185;
wire x_42186;
wire x_42187;
wire x_42188;
wire x_42189;
wire x_42190;
wire x_42191;
wire x_42192;
wire x_42193;
wire x_42194;
wire x_42195;
wire x_42196;
wire x_42197;
wire x_42198;
wire x_42199;
wire x_42200;
wire x_42201;
wire x_42202;
wire x_42203;
wire x_42204;
wire x_42205;
wire x_42206;
wire x_42207;
wire x_42208;
wire x_42209;
wire x_42210;
wire x_42211;
wire x_42212;
wire x_42213;
wire x_42214;
wire x_42215;
wire x_42216;
wire x_42217;
wire x_42218;
wire x_42219;
wire x_42220;
wire x_42221;
wire x_42222;
wire x_42223;
wire x_42224;
wire x_42225;
wire x_42226;
wire x_42227;
wire x_42228;
wire x_42229;
wire x_42230;
wire x_42231;
wire x_42232;
wire x_42233;
wire x_42234;
wire x_42235;
wire x_42236;
wire x_42237;
wire x_42238;
wire x_42239;
wire x_42240;
wire x_42241;
wire x_42242;
wire x_42243;
wire x_42244;
wire x_42245;
wire x_42246;
wire x_42247;
wire x_42248;
wire x_42249;
wire x_42250;
wire x_42251;
wire x_42252;
wire x_42253;
wire x_42254;
wire x_42255;
wire x_42256;
wire x_42257;
wire x_42258;
wire x_42259;
wire x_42260;
wire x_42261;
wire x_42262;
wire x_42263;
wire x_42264;
wire x_42265;
wire x_42266;
wire x_42267;
wire x_42268;
wire x_42269;
wire x_42270;
wire x_42271;
wire x_42272;
wire x_42273;
wire x_42274;
wire x_42275;
wire x_42276;
wire x_42277;
wire x_42278;
wire x_42279;
wire x_42280;
wire x_42281;
wire x_42282;
wire x_42283;
wire x_42284;
wire x_42285;
wire x_42286;
wire x_42287;
wire x_42288;
wire x_42289;
wire x_42290;
wire x_42291;
wire x_42292;
wire x_42293;
wire x_42294;
wire x_42295;
wire x_42296;
wire x_42297;
wire x_42298;
wire x_42299;
wire x_42300;
wire x_42301;
wire x_42302;
wire x_42303;
wire x_42304;
wire x_42305;
wire x_42306;
wire x_42307;
wire x_42308;
wire x_42309;
wire x_42310;
wire x_42311;
wire x_42312;
wire x_42313;
wire x_42314;
wire x_42315;
wire x_42316;
wire x_42317;
wire x_42318;
wire x_42319;
wire x_42320;
wire x_42321;
wire x_42322;
wire x_42323;
wire x_42324;
wire x_42325;
wire x_42326;
wire x_42327;
wire x_42328;
wire x_42329;
wire x_42330;
wire x_42331;
wire x_42332;
wire x_42333;
wire x_42334;
wire x_42335;
wire x_42336;
wire x_42337;
wire x_42338;
wire x_42339;
wire x_42340;
wire x_42341;
wire x_42342;
wire x_42343;
wire x_42344;
wire x_42345;
wire x_42346;
wire x_42347;
wire x_42348;
wire x_42349;
wire x_42350;
wire x_42351;
wire x_42352;
wire x_42353;
wire x_42354;
wire x_42355;
wire x_42356;
wire x_42357;
wire x_42358;
wire x_42359;
wire x_42360;
wire x_42361;
wire x_42362;
wire x_42363;
wire x_42364;
wire x_42365;
wire x_42366;
wire x_42367;
wire x_42368;
wire x_42369;
wire x_42370;
wire x_42371;
wire x_42372;
wire x_42373;
wire x_42374;
wire x_42375;
wire x_42376;
wire x_42377;
wire x_42378;
wire x_42379;
wire x_42380;
wire x_42381;
wire x_42382;
wire x_42383;
wire x_42384;
wire x_42385;
wire x_42386;
wire x_42387;
wire x_42388;
wire x_42389;
wire x_42390;
wire x_42391;
wire x_42392;
wire x_42393;
wire x_42394;
wire x_42395;
wire x_42396;
wire x_42397;
wire x_42398;
wire x_42399;
wire x_42400;
wire x_42401;
wire x_42402;
wire x_42403;
wire x_42404;
wire x_42405;
wire x_42406;
wire x_42407;
wire x_42408;
wire x_42409;
wire x_42410;
wire x_42411;
wire x_42412;
wire x_42413;
wire x_42414;
wire x_42415;
wire x_42416;
wire x_42417;
wire x_42418;
wire x_42419;
wire x_42420;
wire x_42421;
wire x_42422;
wire x_42423;
wire x_42424;
wire x_42425;
wire x_42426;
wire x_42427;
wire x_42428;
wire x_42429;
wire x_42430;
wire x_42431;
wire x_42432;
wire x_42433;
wire x_42434;
wire x_42435;
wire x_42436;
wire x_42437;
wire x_42438;
wire x_42439;
wire x_42440;
wire x_42441;
wire x_42442;
wire x_42443;
wire x_42444;
wire x_42445;
wire x_42446;
wire x_42447;
wire x_42448;
wire x_42449;
wire x_42450;
wire x_42451;
wire x_42452;
wire x_42453;
wire x_42454;
wire x_42455;
wire x_42456;
wire x_42457;
wire x_42458;
wire x_42459;
wire x_42460;
wire x_42461;
wire x_42462;
wire x_42463;
wire x_42464;
wire x_42465;
wire x_42466;
wire x_42467;
wire x_42468;
wire x_42469;
wire x_42470;
wire x_42471;
wire x_42472;
wire x_42473;
wire x_42474;
wire x_42475;
wire x_42476;
wire x_42477;
wire x_42478;
wire x_42479;
wire x_42480;
wire x_42481;
wire x_42482;
wire x_42483;
wire x_42484;
wire x_42485;
wire x_42486;
wire x_42487;
wire x_42488;
wire x_42489;
wire x_42490;
wire x_42491;
wire x_42492;
wire x_42493;
wire x_42494;
wire x_42495;
wire x_42496;
wire x_42497;
wire x_42498;
wire x_42499;
wire x_42500;
wire x_42501;
wire x_42502;
wire x_42503;
wire x_42504;
wire x_42505;
wire x_42506;
wire x_42507;
wire x_42508;
wire x_42509;
wire x_42510;
wire x_42511;
wire x_42512;
wire x_42513;
wire x_42514;
wire x_42515;
wire x_42516;
wire x_42517;
wire x_42518;
wire x_42519;
wire x_42520;
wire x_42521;
wire x_42522;
wire x_42523;
wire x_42524;
wire x_42525;
wire x_42526;
wire x_42527;
wire x_42528;
wire x_42529;
wire x_42530;
wire x_42531;
wire x_42532;
wire x_42533;
wire x_42534;
wire x_42535;
wire x_42536;
wire x_42537;
wire x_42538;
wire x_42539;
wire x_42540;
wire x_42541;
wire x_42542;
wire x_42543;
wire x_42544;
wire x_42545;
wire x_42546;
wire x_42547;
wire x_42548;
wire x_42549;
wire x_42550;
wire x_42551;
wire x_42552;
wire x_42553;
wire x_42554;
wire x_42555;
wire x_42556;
wire x_42557;
wire x_42558;
wire x_42559;
wire x_42560;
wire x_42561;
wire x_42562;
wire x_42563;
wire x_42564;
wire x_42565;
wire x_42566;
wire x_42567;
wire x_42568;
wire x_42569;
wire x_42570;
wire x_42571;
wire x_42572;
wire x_42573;
wire x_42574;
wire x_42575;
wire x_42576;
wire x_42577;
wire x_42578;
wire x_42579;
wire x_42580;
wire x_42581;
wire x_42582;
wire x_42583;
wire x_42584;
wire x_42585;
wire x_42586;
wire x_42587;
wire x_42588;
wire x_42589;
wire x_42590;
wire x_42591;
wire x_42592;
wire x_42593;
wire x_42594;
wire x_42595;
wire x_42596;
wire x_42597;
wire x_42598;
wire x_42599;
wire x_42600;
wire x_42601;
wire x_42602;
wire x_42603;
wire x_42604;
wire x_42605;
wire x_42606;
wire x_42607;
wire x_42608;
wire x_42609;
wire x_42610;
wire x_42611;
wire x_42612;
wire x_42613;
wire x_42614;
wire x_42615;
wire x_42616;
wire x_42617;
wire x_42618;
wire x_42619;
wire x_42620;
wire x_42621;
wire x_42622;
wire x_42623;
wire x_42624;
wire x_42625;
wire x_42626;
wire x_42627;
wire x_42628;
wire x_42629;
wire x_42630;
wire x_42631;
wire x_42632;
wire x_42633;
wire x_42634;
wire x_42635;
wire x_42636;
wire x_42637;
wire x_42638;
wire x_42639;
wire x_42640;
wire x_42641;
wire x_42642;
wire x_42643;
wire x_42644;
wire x_42645;
wire x_42646;
wire x_42647;
wire x_42648;
wire x_42649;
wire x_42650;
wire x_42651;
wire x_42652;
wire x_42653;
wire x_42654;
wire x_42655;
wire x_42656;
wire x_42657;
wire x_42658;
wire x_42659;
wire x_42660;
wire x_42661;
wire x_42662;
wire x_42663;
wire x_42664;
wire x_42665;
wire x_42666;
wire x_42667;
wire x_42668;
wire x_42669;
wire x_42670;
wire x_42671;
wire x_42672;
wire x_42673;
wire x_42674;
wire x_42675;
wire x_42676;
wire x_42677;
wire x_42678;
wire x_42679;
wire x_42680;
wire x_42681;
wire x_42682;
wire x_42683;
wire x_42684;
wire x_42685;
wire x_42686;
wire x_42687;
wire x_42688;
wire x_42689;
wire x_42690;
wire x_42691;
wire x_42692;
wire x_42693;
wire x_42694;
wire x_42695;
wire x_42696;
wire x_42697;
wire x_42698;
wire x_42699;
wire x_42700;
wire x_42701;
wire x_42702;
wire x_42703;
wire x_42704;
wire x_42705;
wire x_42706;
wire x_42707;
wire x_42708;
wire x_42709;
wire x_42710;
wire x_42711;
wire x_42712;
wire x_42713;
wire x_42714;
wire x_42715;
wire x_42716;
wire x_42717;
wire x_42718;
wire x_42719;
wire x_42720;
wire x_42721;
wire x_42722;
wire x_42723;
wire x_42724;
wire x_42725;
wire x_42726;
wire x_42727;
wire x_42728;
wire x_42729;
wire x_42730;
wire x_42731;
wire x_42732;
wire x_42733;
wire x_42734;
wire x_42735;
wire x_42736;
wire x_42737;
wire x_42738;
wire x_42739;
wire x_42740;
wire x_42741;
wire x_42742;
wire x_42743;
wire x_42744;
wire x_42745;
wire x_42746;
wire x_42747;
wire x_42748;
wire x_42749;
wire x_42750;
wire x_42751;
wire x_42752;
wire x_42753;
wire x_42754;
wire x_42755;
wire x_42756;
wire x_42757;
wire x_42758;
wire x_42759;
wire x_42760;
wire x_42761;
wire x_42762;
wire x_42763;
wire x_42764;
wire x_42765;
wire x_42766;
wire x_42767;
wire x_42768;
wire x_42769;
wire x_42770;
wire x_42771;
wire x_42772;
wire x_42773;
wire x_42774;
wire x_42775;
wire x_42776;
wire x_42777;
wire x_42778;
wire x_42779;
wire x_42780;
wire x_42781;
wire x_42782;
wire x_42783;
wire x_42784;
wire x_42785;
wire x_42786;
wire x_42787;
wire x_42788;
wire x_42789;
wire x_42790;
wire x_42791;
wire x_42792;
wire x_42793;
wire x_42794;
wire x_42795;
wire x_42796;
wire x_42797;
wire x_42798;
wire x_42799;
wire x_42800;
wire x_42801;
wire x_42802;
wire x_42803;
wire x_42804;
wire x_42805;
wire x_42806;
wire x_42807;
wire x_42808;
wire x_42809;
wire x_42810;
wire x_42811;
wire x_42812;
wire x_42813;
wire x_42814;
wire x_42815;
wire x_42816;
wire x_42817;
wire x_42818;
wire x_42819;
wire x_42820;
wire x_42821;
wire x_42822;
wire x_42823;
wire x_42824;
wire x_42825;
wire x_42826;
wire x_42827;
wire x_42828;
wire x_42829;
wire x_42830;
wire x_42831;
wire x_42832;
wire x_42833;
wire x_42834;
wire x_42835;
wire x_42836;
wire x_42837;
wire x_42838;
wire x_42839;
wire x_42840;
wire x_42841;
wire x_42842;
wire x_42843;
wire x_42844;
wire x_42845;
wire x_42846;
wire x_42847;
wire x_42848;
wire x_42849;
wire x_42850;
wire x_42851;
wire x_42852;
wire x_42853;
wire x_42854;
wire x_42855;
wire x_42856;
wire x_42857;
wire x_42858;
wire x_42859;
wire x_42860;
wire x_42861;
wire x_42862;
wire x_42863;
wire x_42864;
wire x_42865;
wire x_42866;
wire x_42867;
wire x_42868;
wire x_42869;
wire x_42870;
wire x_42871;
wire x_42872;
wire x_42873;
wire x_42874;
wire x_42875;
wire x_42876;
wire x_42877;
wire x_42878;
wire x_42879;
wire x_42880;
wire x_42881;
wire x_42882;
wire x_42883;
wire x_42884;
wire x_42885;
wire x_42886;
wire x_42887;
wire x_42888;
wire x_42889;
wire x_42890;
wire x_42891;
wire x_42892;
wire x_42893;
wire x_42894;
wire x_42895;
wire x_42896;
wire x_42897;
wire x_42898;
wire x_42899;
wire x_42900;
wire x_42901;
wire x_42902;
wire x_42903;
wire x_42904;
wire x_42905;
wire x_42906;
wire x_42907;
wire x_42908;
wire x_42909;
wire x_42910;
wire x_42911;
wire x_42912;
wire x_42913;
wire x_42914;
wire x_42915;
wire x_42916;
wire x_42917;
wire x_42918;
wire x_42919;
wire x_42920;
wire x_42921;
wire x_42922;
wire x_42923;
wire x_42924;
wire x_42925;
wire x_42926;
wire x_42927;
wire x_42928;
wire x_42929;
wire x_42930;
wire x_42931;
wire x_42932;
wire x_42933;
wire x_42934;
wire x_42935;
wire x_42936;
wire x_42937;
wire x_42938;
wire x_42939;
wire x_42940;
wire x_42941;
wire x_42942;
wire x_42943;
wire x_42944;
wire x_42945;
wire x_42946;
wire x_42947;
wire x_42948;
wire x_42949;
wire x_42950;
wire x_42951;
wire x_42952;
wire x_42953;
wire x_42954;
wire x_42955;
wire x_42956;
wire x_42957;
wire x_42958;
wire x_42959;
wire x_42960;
wire x_42961;
wire x_42962;
wire x_42963;
wire x_42964;
wire x_42965;
wire x_42966;
wire x_42967;
wire x_42968;
wire x_42969;
wire x_42970;
wire x_42971;
wire x_42972;
wire x_42973;
wire x_42974;
wire x_42975;
wire x_42976;
wire x_42977;
wire x_42978;
wire x_42979;
wire x_42980;
wire x_42981;
wire x_42982;
wire x_42983;
wire x_42984;
wire x_42985;
wire x_42986;
wire x_42987;
wire x_42988;
wire x_42989;
wire x_42990;
wire x_42991;
wire x_42992;
wire x_42993;
wire x_42994;
wire x_42995;
wire x_42996;
wire x_42997;
wire x_42998;
wire x_42999;
wire x_43000;
wire x_43001;
wire x_43002;
wire x_43003;
wire x_43004;
wire x_43005;
wire x_43006;
wire x_43007;
wire x_43008;
wire x_43009;
wire x_43010;
wire x_43011;
wire x_43012;
wire x_43013;
wire x_43014;
wire x_43015;
wire x_43016;
wire x_43017;
wire x_43018;
wire x_43019;
wire x_43020;
wire x_43021;
wire x_43022;
wire x_43023;
wire x_43024;
wire x_43025;
wire x_43026;
wire x_43027;
wire x_43028;
wire x_43029;
wire x_43030;
wire x_43031;
wire x_43032;
wire x_43033;
wire x_43034;
wire x_43035;
wire x_43036;
wire x_43037;
wire x_43038;
wire x_43039;
wire x_43040;
wire x_43041;
wire x_43042;
wire x_43043;
wire x_43044;
wire x_43045;
wire x_43046;
wire x_43047;
wire x_43048;
wire x_43049;
wire x_43050;
wire x_43051;
wire x_43052;
wire x_43053;
wire x_43054;
wire x_43055;
wire x_43056;
wire x_43057;
wire x_43058;
wire x_43059;
wire x_43060;
wire x_43061;
wire x_43062;
wire x_43063;
wire x_43064;
wire x_43065;
wire x_43066;
wire x_43067;
wire x_43068;
wire x_43069;
wire x_43070;
wire x_43071;
wire x_43072;
wire x_43073;
wire x_43074;
wire x_43075;
wire x_43076;
wire x_43077;
wire x_43078;
wire x_43079;
wire x_43080;
wire x_43081;
wire x_43082;
wire x_43083;
wire x_43084;
wire x_43085;
wire x_43086;
wire x_43087;
wire x_43088;
wire x_43089;
wire x_43090;
wire x_43091;
wire x_43092;
wire x_43093;
wire x_43094;
wire x_43095;
wire x_43096;
wire x_43097;
wire x_43098;
wire x_43099;
wire x_43100;
wire x_43101;
wire x_43102;
wire x_43103;
wire x_43104;
wire x_43105;
wire x_43106;
wire x_43107;
wire x_43108;
wire x_43109;
wire x_43110;
wire x_43111;
wire x_43112;
wire x_43113;
wire x_43114;
wire x_43115;
wire x_43116;
wire x_43117;
wire x_43118;
wire x_43119;
wire x_43120;
wire x_43121;
wire x_43122;
wire x_43123;
wire x_43124;
wire x_43125;
wire x_43126;
wire x_43127;
wire x_43128;
wire x_43129;
wire x_43130;
wire x_43131;
wire x_43132;
wire x_43133;
wire x_43134;
wire x_43135;
wire x_43136;
wire x_43137;
wire x_43138;
wire x_43139;
wire x_43140;
wire x_43141;
wire x_43142;
wire x_43143;
wire x_43144;
wire x_43145;
wire x_43146;
wire x_43147;
wire x_43148;
wire x_43149;
wire x_43150;
wire x_43151;
wire x_43152;
wire x_43153;
wire x_43154;
wire x_43155;
wire x_43156;
wire x_43157;
wire x_43158;
wire x_43159;
wire x_43160;
wire x_43161;
wire x_43162;
wire x_43163;
wire x_43164;
wire x_43165;
wire x_43166;
wire x_43167;
wire x_43168;
wire x_43169;
wire x_43170;
wire x_43171;
wire x_43172;
wire x_43173;
wire x_43174;
wire x_43175;
wire x_43176;
wire x_43177;
wire x_43178;
wire x_43179;
wire x_43180;
wire x_43181;
wire x_43182;
wire x_43183;
wire x_43184;
wire x_43185;
wire x_43186;
wire x_43187;
wire x_43188;
wire x_43189;
wire x_43190;
wire x_43191;
wire x_43192;
wire x_43193;
wire x_43194;
wire x_43195;
wire x_43196;
wire x_43197;
wire x_43198;
wire x_43199;
wire x_43200;
wire x_43201;
wire x_43202;
wire x_43203;
wire x_43204;
wire x_43205;
wire x_43206;
wire x_43207;
wire x_43208;
wire x_43209;
wire x_43210;
wire x_43211;
wire x_43212;
wire x_43213;
wire x_43214;
wire x_43215;
wire x_43216;
wire x_43217;
wire x_43218;
wire x_43219;
wire x_43220;
wire x_43221;
wire x_43222;
wire x_43223;
wire x_43224;
wire x_43225;
wire x_43226;
wire x_43227;
wire x_43228;
wire x_43229;
wire x_43230;
wire x_43231;
wire x_43232;
wire x_43233;
wire x_43234;
wire x_43235;
wire x_43236;
wire x_43237;
wire x_43238;
wire x_43239;
wire x_43240;
wire x_43241;
wire x_43242;
wire x_43243;
wire x_43244;
wire x_43245;
wire x_43246;
wire x_43247;
wire x_43248;
wire x_43249;
wire x_43250;
wire x_43251;
wire x_43252;
wire x_43253;
wire x_43254;
wire x_43255;
wire x_43256;
wire x_43257;
wire x_43258;
wire x_43259;
wire x_43260;
wire x_43261;
wire x_43262;
wire x_43263;
wire x_43264;
wire x_43265;
wire x_43266;
wire x_43267;
wire x_43268;
wire x_43269;
wire x_43270;
wire x_43271;
wire x_43272;
wire x_43273;
wire x_43274;
wire x_43275;
wire x_43276;
wire x_43277;
wire x_43278;
wire x_43279;
wire x_43280;
wire x_43281;
wire x_43282;
wire x_43283;
wire x_43284;
wire x_43285;
wire x_43286;
wire x_43287;
wire x_43288;
wire x_43289;
wire x_43290;
wire x_43291;
wire x_43292;
wire x_43293;
wire x_43294;
wire x_43295;
wire x_43296;
wire x_43297;
wire x_43298;
wire x_43299;
wire x_43300;
wire x_43301;
wire x_43302;
wire x_43303;
wire x_43304;
wire x_43305;
wire x_43306;
wire x_43307;
wire x_43308;
wire x_43309;
wire x_43310;
wire x_43311;
wire x_43312;
wire x_43313;
wire x_43314;
wire x_43315;
wire x_43316;
wire x_43317;
wire x_43318;
wire x_43319;
wire x_43320;
wire x_43321;
wire x_43322;
wire x_43323;
wire x_43324;
wire x_43325;
wire x_43326;
wire x_43327;
wire x_43328;
wire x_43329;
wire x_43330;
wire x_43331;
wire x_43332;
wire x_43333;
wire x_43334;
wire x_43335;
wire x_43336;
wire x_43337;
wire x_43338;
wire x_43339;
wire x_43340;
wire x_43341;
wire x_43342;
wire x_43343;
wire x_43344;
wire x_43345;
wire x_43346;
wire x_43347;
wire x_43348;
wire x_43349;
wire x_43350;
wire x_43351;
wire x_43352;
wire x_43353;
wire x_43354;
wire x_43355;
wire x_43356;
wire x_43357;
wire x_43358;
wire x_43359;
wire x_43360;
wire x_43361;
wire x_43362;
wire x_43363;
wire x_43364;
wire x_43365;
wire x_43366;
wire x_43367;
wire x_43368;
wire x_43369;
wire x_43370;
wire x_43371;
wire x_43372;
wire x_43373;
wire x_43374;
wire x_43375;
wire x_43376;
wire x_43377;
wire x_43378;
wire x_43379;
wire x_43380;
wire x_43381;
wire x_43382;
wire x_43383;
wire x_43384;
wire x_43385;
wire x_43386;
wire x_43387;
wire x_43388;
wire x_43389;
wire x_43390;
wire x_43391;
wire x_43392;
wire x_43393;
wire x_43394;
wire x_43395;
wire x_43396;
wire x_43397;
wire x_43398;
wire x_43399;
wire x_43400;
wire x_43401;
wire x_43402;
wire x_43403;
wire x_43404;
wire x_43405;
wire x_43406;
wire x_43407;
wire x_43408;
wire x_43409;
wire x_43410;
wire x_43411;
wire x_43412;
wire x_43413;
wire x_43414;
wire x_43415;
wire x_43416;
wire x_43417;
wire x_43418;
wire x_43419;
wire x_43420;
wire x_43421;
wire x_43422;
wire x_43423;
wire x_43424;
wire x_43425;
wire x_43426;
wire x_43427;
wire x_43428;
wire x_43429;
wire x_43430;
wire x_43431;
wire x_43432;
wire x_43433;
wire x_43434;
wire x_43435;
wire x_43436;
wire x_43437;
wire x_43438;
wire x_43439;
wire x_43440;
wire x_43441;
wire x_43442;
wire x_43443;
wire x_43444;
wire x_43445;
wire x_43446;
wire x_43447;
wire x_43448;
wire x_43449;
wire x_43450;
wire x_43451;
wire x_43452;
wire x_43453;
wire x_43454;
wire x_43455;
wire x_43456;
wire x_43457;
wire x_43458;
wire x_43459;
wire x_43460;
wire x_43461;
wire x_43462;
wire x_43463;
wire x_43464;
wire x_43465;
wire x_43466;
wire x_43467;
wire x_43468;
wire x_43469;
wire x_43470;
wire x_43471;
wire x_43472;
wire x_43473;
wire x_43474;
wire x_43475;
wire x_43476;
wire x_43477;
wire x_43478;
wire x_43479;
wire x_43480;
wire x_43481;
wire x_43482;
wire x_43483;
wire x_43484;
wire x_43485;
wire x_43486;
wire x_43487;
wire x_43488;
wire x_43489;
wire x_43490;
wire x_43491;
wire x_43492;
wire x_43493;
wire x_43494;
wire x_43495;
wire x_43496;
wire x_43497;
wire x_43498;
wire x_43499;
wire x_43500;
wire x_43501;
wire x_43502;
wire x_43503;
wire x_43504;
wire x_43505;
wire x_43506;
wire x_43507;
wire x_43508;
wire x_43509;
wire x_43510;
wire x_43511;
wire x_43512;
wire x_43513;
wire x_43514;
wire x_43515;
wire x_43516;
wire x_43517;
wire x_43518;
wire x_43519;
wire x_43520;
wire x_43521;
wire x_43522;
wire x_43523;
wire x_43524;
wire x_43525;
wire x_43526;
wire x_43527;
wire x_43528;
wire x_43529;
wire x_43530;
wire x_43531;
wire x_43532;
wire x_43533;
wire x_43534;
wire x_43535;
wire x_43536;
wire x_43537;
wire x_43538;
wire x_43539;
wire x_43540;
wire x_43541;
wire x_43542;
wire x_43543;
wire x_43544;
wire x_43545;
wire x_43546;
wire x_43547;
wire x_43548;
wire x_43549;
wire x_43550;
wire x_43551;
wire x_43552;
wire x_43553;
wire x_43554;
wire x_43555;
wire x_43556;
wire x_43557;
wire x_43558;
wire x_43559;
wire x_43560;
wire x_43561;
wire x_43562;
wire x_43563;
wire x_43564;
wire x_43565;
wire x_43566;
wire x_43567;
wire x_43568;
wire x_43569;
wire x_43570;
wire x_43571;
wire x_43572;
wire x_43573;
wire x_43574;
wire x_43575;
wire x_43576;
wire x_43577;
wire x_43578;
wire x_43579;
wire x_43580;
wire x_43581;
wire x_43582;
wire x_43583;
wire x_43584;
wire x_43585;
wire x_43586;
wire x_43587;
wire x_43588;
wire x_43589;
wire x_43590;
wire x_43591;
wire x_43592;
wire x_43593;
wire x_43594;
wire x_43595;
wire x_43596;
wire x_43597;
wire x_43598;
wire x_43599;
wire x_43600;
wire x_43601;
wire x_43602;
wire x_43603;
wire x_43604;
wire x_43605;
wire x_43606;
wire x_43607;
wire x_43608;
wire x_43609;
wire x_43610;
wire x_43611;
wire x_43612;
wire x_43613;
wire x_43614;
wire x_43615;
wire x_43616;
wire x_43617;
wire x_43618;
wire x_43619;
wire x_43620;
wire x_43621;
wire x_43622;
wire x_43623;
wire x_43624;
wire x_43625;
wire x_43626;
wire x_43627;
wire x_43628;
wire x_43629;
wire x_43630;
wire x_43631;
wire x_43632;
wire x_43633;
wire x_43634;
wire x_43635;
wire x_43636;
wire x_43637;
wire x_43638;
wire x_43639;
wire x_43640;
wire x_43641;
wire x_43642;
wire x_43643;
wire x_43644;
wire x_43645;
wire x_43646;
wire x_43647;
wire x_43648;
wire x_43649;
wire x_43650;
wire x_43651;
wire x_43652;
wire x_43653;
wire x_43654;
wire x_43655;
wire x_43656;
wire x_43657;
wire x_43658;
wire x_43659;
wire x_43660;
wire x_43661;
wire x_43662;
wire x_43663;
wire x_43664;
wire x_43665;
wire x_43666;
wire x_43667;
wire x_43668;
wire x_43669;
wire x_43670;
wire x_43671;
wire x_43672;
wire x_43673;
wire x_43674;
wire x_43675;
wire x_43676;
wire x_43677;
wire x_43678;
wire x_43679;
wire x_43680;
wire x_43681;
wire x_43682;
wire x_43683;
wire x_43684;
wire x_43685;
wire x_43686;
wire x_43687;
wire x_43688;
wire x_43689;
wire x_43690;
wire x_43691;
wire x_43692;
wire x_43693;
wire x_43694;
wire x_43695;
wire x_43696;
wire x_43697;
wire x_43698;
wire x_43699;
wire x_43700;
wire x_43701;
wire x_43702;
wire x_43703;
wire x_43704;
wire x_43705;
wire x_43706;
wire x_43707;
wire x_43708;
wire x_43709;
wire x_43710;
wire x_43711;
wire x_43712;
wire x_43713;
wire x_43714;
wire x_43715;
wire x_43716;
wire x_43717;
wire x_43718;
wire x_43719;
wire x_43720;
wire x_43721;
wire x_43722;
wire x_43723;
wire x_43724;
wire x_43725;
wire x_43726;
wire x_43727;
wire x_43728;
wire x_43729;
wire x_43730;
wire x_43731;
wire x_43732;
wire x_43733;
wire x_43734;
wire x_43735;
wire x_43736;
wire x_43737;
wire x_43738;
wire x_43739;
wire x_43740;
wire x_43741;
wire x_43742;
wire x_43743;
wire x_43744;
wire x_43745;
wire x_43746;
wire x_43747;
wire x_43748;
wire x_43749;
wire x_43750;
wire x_43751;
wire x_43752;
wire x_43753;
wire x_43754;
wire x_43755;
wire x_43756;
wire x_43757;
wire x_43758;
wire x_43759;
wire x_43760;
wire x_43761;
wire x_43762;
wire x_43763;
wire x_43764;
wire x_43765;
wire x_43766;
wire x_43767;
wire x_43768;
wire x_43769;
wire x_43770;
wire x_43771;
wire x_43772;
wire x_43773;
wire x_43774;
wire x_43775;
wire x_43776;
wire x_43777;
wire x_43778;
wire x_43779;
wire x_43780;
wire x_43781;
wire x_43782;
wire x_43783;
wire x_43784;
wire x_43785;
wire x_43786;
wire x_43787;
wire x_43788;
wire x_43789;
wire x_43790;
wire x_43791;
wire x_43792;
wire x_43793;
wire x_43794;
wire x_43795;
wire x_43796;
wire x_43797;
wire x_43798;
wire x_43799;
wire x_43800;
wire x_43801;
wire x_43802;
wire x_43803;
wire x_43804;
wire x_43805;
wire x_43806;
wire x_43807;
wire x_43808;
wire x_43809;
wire x_43810;
wire x_43811;
wire x_43812;
wire x_43813;
wire x_43814;
wire x_43815;
wire x_43816;
wire x_43817;
wire x_43818;
wire x_43819;
wire x_43820;
wire x_43821;
wire x_43822;
wire x_43823;
wire x_43824;
wire x_43825;
wire x_43826;
wire x_43827;
wire x_43828;
wire x_43829;
wire x_43830;
wire x_43831;
wire x_43832;
wire x_43833;
wire x_43834;
wire x_43835;
wire x_43836;
wire x_43837;
wire x_43838;
wire x_43839;
wire x_43840;
wire x_43841;
wire x_43842;
wire x_43843;
wire x_43844;
wire x_43845;
wire x_43846;
wire x_43847;
wire x_43848;
wire x_43849;
wire x_43850;
wire x_43851;
wire x_43852;
wire x_43853;
wire x_43854;
wire x_43855;
wire x_43856;
wire x_43857;
wire x_43858;
wire x_43859;
wire x_43860;
wire x_43861;
wire x_43862;
wire x_43863;
wire x_43864;
wire x_43865;
wire x_43866;
wire x_43867;
wire x_43868;
wire x_43869;
wire x_43870;
wire x_43871;
wire x_43872;
wire x_43873;
wire x_43874;
wire x_43875;
wire x_43876;
wire x_43877;
wire x_43878;
wire x_43879;
wire x_43880;
wire x_43881;
wire x_43882;
wire x_43883;
wire x_43884;
wire x_43885;
wire x_43886;
wire x_43887;
wire x_43888;
wire x_43889;
wire x_43890;
wire x_43891;
wire x_43892;
wire x_43893;
wire x_43894;
wire x_43895;
wire x_43896;
wire x_43897;
wire x_43898;
wire x_43899;
wire x_43900;
wire x_43901;
wire x_43902;
wire x_43903;
wire x_43904;
wire x_43905;
wire x_43906;
wire x_43907;
wire x_43908;
wire x_43909;
wire x_43910;
wire x_43911;
wire x_43912;
wire x_43913;
wire x_43914;
wire x_43915;
wire x_43916;
wire x_43917;
wire x_43918;
wire x_43919;
wire x_43920;
wire x_43921;
wire x_43922;
wire x_43923;
wire x_43924;
wire x_43925;
wire x_43926;
wire x_43927;
wire x_43928;
wire x_43929;
wire x_43930;
wire x_43931;
wire x_43932;
wire x_43933;
wire x_43934;
wire x_43935;
wire x_43936;
wire x_43937;
wire x_43938;
wire x_43939;
wire x_43940;
wire x_43941;
wire x_43942;
wire x_43943;
wire x_43944;
wire x_43945;
wire x_43946;
wire x_43947;
wire x_43948;
wire x_43949;
wire x_43950;
wire x_43951;
wire x_43952;
wire x_43953;
wire x_43954;
wire x_43955;
wire x_43956;
wire x_43957;
wire x_43958;
wire x_43959;
wire x_43960;
wire x_43961;
wire x_43962;
wire x_43963;
wire x_43964;
wire x_43965;
wire x_43966;
wire x_43967;
wire x_43968;
wire x_43969;
wire x_43970;
wire x_43971;
wire x_43972;
wire x_43973;
wire x_43974;
wire x_43975;
wire x_43976;
wire x_43977;
wire x_43978;
wire x_43979;
wire x_43980;
wire x_43981;
wire x_43982;
wire x_43983;
wire x_43984;
wire x_43985;
wire x_43986;
wire x_43987;
wire x_43988;
wire x_43989;
wire x_43990;
wire x_43991;
wire x_43992;
wire x_43993;
wire x_43994;
wire x_43995;
wire x_43996;
wire x_43997;
wire x_43998;
wire x_43999;
wire x_44000;
wire x_44001;
wire x_44002;
wire x_44003;
wire x_44004;
wire x_44005;
wire x_44006;
wire x_44007;
wire x_44008;
wire x_44009;
wire x_44010;
wire x_44011;
wire x_44012;
wire x_44013;
wire x_44014;
wire x_44015;
wire x_44016;
wire x_44017;
wire x_44018;
wire x_44019;
wire x_44020;
wire x_44021;
wire x_44022;
wire x_44023;
wire x_44024;
wire x_44025;
wire x_44026;
wire x_44027;
wire x_44028;
wire x_44029;
wire x_44030;
wire x_44031;
wire x_44032;
wire x_44033;
wire x_44034;
wire x_44035;
wire x_44036;
wire x_44037;
wire x_44038;
wire x_44039;
wire x_44040;
wire x_44041;
wire x_44042;
wire x_44043;
wire x_44044;
wire x_44045;
wire x_44046;
wire x_44047;
wire x_44048;
wire x_44049;
wire x_44050;
wire x_44051;
wire x_44052;
wire x_44053;
wire x_44054;
wire x_44055;
wire x_44056;
wire x_44057;
wire x_44058;
wire x_44059;
wire x_44060;
wire x_44061;
wire x_44062;
wire x_44063;
wire x_44064;
wire x_44065;
wire x_44066;
wire x_44067;
wire x_44068;
wire x_44069;
wire x_44070;
wire x_44071;
wire x_44072;
wire x_44073;
wire x_44074;
wire x_44075;
wire x_44076;
wire x_44077;
wire x_44078;
wire x_44079;
wire x_44080;
wire x_44081;
wire x_44082;
wire x_44083;
wire x_44084;
wire x_44085;
wire x_44086;
wire x_44087;
wire x_44088;
wire x_44089;
wire x_44090;
wire x_44091;
wire x_44092;
wire x_44093;
wire x_44094;
wire x_44095;
wire x_44096;
wire x_44097;
wire x_44098;
wire x_44099;
wire x_44100;
wire x_44101;
wire x_44102;
wire x_44103;
wire x_44104;
wire x_44105;
wire x_44106;
wire x_44107;
wire x_44108;
wire x_44109;
wire x_44110;
wire x_44111;
wire x_44112;
wire x_44113;
wire x_44114;
wire x_44115;
wire x_44116;
wire x_44117;
wire x_44118;
wire x_44119;
wire x_44120;
wire x_44121;
wire x_44122;
wire x_44123;
wire x_44124;
wire x_44125;
wire x_44126;
wire x_44127;
wire x_44128;
wire x_44129;
wire x_44130;
wire x_44131;
wire x_44132;
wire x_44133;
wire x_44134;
wire x_44135;
wire x_44136;
wire x_44137;
wire x_44138;
wire x_44139;
wire x_44140;
wire x_44141;
wire x_44142;
wire x_44143;
wire x_44144;
wire x_44145;
wire x_44146;
wire x_44147;
wire x_44148;
wire x_44149;
wire x_44150;
wire x_44151;
wire x_44152;
wire x_44153;
wire x_44154;
wire x_44155;
wire x_44156;
wire x_44157;
wire x_44158;
wire x_44159;
wire x_44160;
wire x_44161;
wire x_44162;
wire x_44163;
wire x_44164;
wire x_44165;
wire x_44166;
wire x_44167;
wire x_44168;
wire x_44169;
wire x_44170;
wire x_44171;
wire x_44172;
wire x_44173;
wire x_44174;
wire x_44175;
wire x_44176;
wire x_44177;
wire x_44178;
wire x_44179;
wire x_44180;
wire x_44181;
wire x_44182;
wire x_44183;
wire x_44184;
wire x_44185;
wire x_44186;
wire x_44187;
wire x_44188;
wire x_44189;
wire x_44190;
wire x_44191;
wire x_44192;
wire x_44193;
wire x_44194;
wire x_44195;
wire x_44196;
wire x_44197;
wire x_44198;
wire x_44199;
wire x_44200;
wire x_44201;
wire x_44202;
wire x_44203;
wire x_44204;
wire x_44205;
wire x_44206;
wire x_44207;
wire x_44208;
wire x_44209;
wire x_44210;
wire x_44211;
wire x_44212;
wire x_44213;
wire x_44214;
wire x_44215;
wire x_44216;
wire x_44217;
wire x_44218;
wire x_44219;
wire x_44220;
wire x_44221;
wire x_44222;
wire x_44223;
wire x_44224;
wire x_44225;
wire x_44226;
wire x_44227;
wire x_44228;
wire x_44229;
wire x_44230;
wire x_44231;
wire x_44232;
wire x_44233;
wire x_44234;
wire x_44235;
wire x_44236;
wire x_44237;
wire x_44238;
wire x_44239;
wire x_44240;
wire x_44241;
wire x_44242;
wire x_44243;
wire x_44244;
wire x_44245;
wire x_44246;
wire x_44247;
wire x_44248;
wire x_44249;
wire x_44250;
wire x_44251;
wire x_44252;
wire x_44253;
wire x_44254;
wire x_44255;
wire x_44256;
wire x_44257;
wire x_44258;
wire x_44259;
wire x_44260;
wire x_44261;
wire x_44262;
wire x_44263;
wire x_44264;
wire x_44265;
wire x_44266;
wire x_44267;
wire x_44268;
wire x_44269;
wire x_44270;
wire x_44271;
wire x_44272;
wire x_44273;
wire x_44274;
wire x_44275;
wire x_44276;
wire x_44277;
wire x_44278;
wire x_44279;
wire x_44280;
wire x_44281;
wire x_44282;
wire x_44283;
wire x_44284;
wire x_44285;
wire x_44286;
wire x_44287;
wire x_44288;
wire x_44289;
wire x_44290;
wire x_44291;
wire x_44292;
wire x_44293;
wire x_44294;
wire x_44295;
wire x_44296;
wire x_44297;
wire x_44298;
wire x_44299;
wire x_44300;
wire x_44301;
wire x_44302;
wire x_44303;
wire x_44304;
wire x_44305;
wire x_44306;
wire x_44307;
wire x_44308;
wire x_44309;
wire x_44310;
wire x_44311;
wire x_44312;
wire x_44313;
wire x_44314;
wire x_44315;
wire x_44316;
wire x_44317;
wire x_44318;
wire x_44319;
wire x_44320;
wire x_44321;
wire x_44322;
wire x_44323;
wire x_44324;
wire x_44325;
wire x_44326;
wire x_44327;
wire x_44328;
wire x_44329;
wire x_44330;
wire x_44331;
wire x_44332;
wire x_44333;
wire x_44334;
wire x_44335;
wire x_44336;
wire x_44337;
wire x_44338;
wire x_44339;
wire x_44340;
wire x_44341;
wire x_44342;
wire x_44343;
wire x_44344;
wire x_44345;
wire x_44346;
wire x_44347;
wire x_44348;
wire x_44349;
wire x_44350;
wire x_44351;
wire x_44352;
wire x_44353;
wire x_44354;
wire x_44355;
wire x_44356;
wire x_44357;
wire x_44358;
wire x_44359;
wire x_44360;
wire x_44361;
wire x_44362;
wire x_44363;
wire x_44364;
wire x_44365;
wire x_44366;
wire x_44367;
wire x_44368;
wire x_44369;
wire x_44370;
wire x_44371;
wire x_44372;
wire x_44373;
wire x_44374;
wire x_44375;
wire x_44376;
wire x_44377;
wire x_44378;
wire x_44379;
wire x_44380;
wire x_44381;
wire x_44382;
wire x_44383;
wire x_44384;
wire x_44385;
wire x_44386;
wire x_44387;
wire x_44388;
wire x_44389;
wire x_44390;
wire x_44391;
wire x_44392;
wire x_44393;
wire x_44394;
wire x_44395;
wire x_44396;
wire x_44397;
wire x_44398;
wire x_44399;
wire x_44400;
wire x_44401;
wire x_44402;
wire x_44403;
wire x_44404;
wire x_44405;
wire x_44406;
wire x_44407;
wire x_44408;
wire x_44409;
wire x_44410;
wire x_44411;
wire x_44412;
wire x_44413;
wire x_44414;
wire x_44415;
wire x_44416;
wire x_44417;
wire x_44418;
wire x_44419;
wire x_44420;
wire x_44421;
wire x_44422;
wire x_44423;
wire x_44424;
wire x_44425;
wire x_44426;
wire x_44427;
wire x_44428;
wire x_44429;
wire x_44430;
wire x_44431;
wire x_44432;
wire x_44433;
wire x_44434;
wire x_44435;
wire x_44436;
wire x_44437;
wire x_44438;
wire x_44439;
wire x_44440;
wire x_44441;
wire x_44442;
wire x_44443;
wire x_44444;
wire x_44445;
wire x_44446;
wire x_44447;
wire x_44448;
wire x_44449;
wire x_44450;
wire x_44451;
wire x_44452;
wire x_44453;
wire x_44454;
wire x_44455;
wire x_44456;
wire x_44457;
wire x_44458;
wire x_44459;
wire x_44460;
wire x_44461;
wire x_44462;
wire x_44463;
wire x_44464;
wire x_44465;
wire x_44466;
wire x_44467;
wire x_44468;
wire x_44469;
wire x_44470;
wire x_44471;
wire x_44472;
wire x_44473;
wire x_44474;
wire x_44475;
wire x_44476;
wire x_44477;
wire x_44478;
wire x_44479;
wire x_44480;
wire x_44481;
wire x_44482;
wire x_44483;
wire x_44484;
wire x_44485;
wire x_44486;
wire x_44487;
wire x_44488;
wire x_44489;
wire x_44490;
wire x_44491;
wire x_44492;
wire x_44493;
wire x_44494;
wire x_44495;
wire x_44496;
wire x_44497;
wire x_44498;
wire x_44499;
wire x_44500;
wire x_44501;
wire x_44502;
wire x_44503;
wire x_44504;
wire x_44505;
wire x_44506;
wire x_44507;
wire x_44508;
wire x_44509;
wire x_44510;
wire x_44511;
wire x_44512;
wire x_44513;
wire x_44514;
wire x_44515;
wire x_44516;
wire x_44517;
wire x_44518;
wire x_44519;
wire x_44520;
wire x_44521;
wire x_44522;
wire x_44523;
wire x_44524;
wire x_44525;
wire x_44526;
wire x_44527;
wire x_44528;
wire x_44529;
wire x_44530;
wire x_44531;
wire x_44532;
wire x_44533;
wire x_44534;
wire x_44535;
wire x_44536;
wire x_44537;
wire x_44538;
wire x_44539;
wire x_44540;
wire x_44541;
wire x_44542;
wire x_44543;
wire x_44544;
wire x_44545;
wire x_44546;
wire x_44547;
wire x_44548;
wire x_44549;
wire x_44550;
wire x_44551;
wire x_44552;
wire x_44553;
wire x_44554;
wire x_44555;
wire x_44556;
wire x_44557;
wire x_44558;
wire x_44559;
wire x_44560;
wire x_44561;
wire x_44562;
wire x_44563;
wire x_44564;
wire x_44565;
wire x_44566;
wire x_44567;
wire x_44568;
wire x_44569;
wire x_44570;
wire x_44571;
wire x_44572;
wire x_44573;
wire x_44574;
wire x_44575;
wire x_44576;
wire x_44577;
wire x_44578;
wire x_44579;
wire x_44580;
wire x_44581;
wire x_44582;
wire x_44583;
wire x_44584;
wire x_44585;
wire x_44586;
wire x_44587;
wire x_44588;
wire x_44589;
wire x_44590;
wire x_44591;
wire x_44592;
wire x_44593;
wire x_44594;
wire x_44595;
wire x_44596;
wire x_44597;
wire x_44598;
wire x_44599;
wire x_44600;
wire x_44601;
wire x_44602;
wire x_44603;
wire x_44604;
wire x_44605;
wire x_44606;
wire x_44607;
wire x_44608;
wire x_44609;
wire x_44610;
wire x_44611;
wire x_44612;
wire x_44613;
wire x_44614;
wire x_44615;
wire x_44616;
wire x_44617;
wire x_44618;
wire x_44619;
wire x_44620;
wire x_44621;
wire x_44622;
wire x_44623;
wire x_44624;
wire x_44625;
wire x_44626;
wire x_44627;
wire x_44628;
wire x_44629;
wire x_44630;
wire x_44631;
wire x_44632;
wire x_44633;
wire x_44634;
wire x_44635;
wire x_44636;
wire x_44637;
wire x_44638;
wire x_44639;
wire x_44640;
wire x_44641;
wire x_44642;
wire x_44643;
wire x_44644;
wire x_44645;
wire x_44646;
wire x_44647;
wire x_44648;
wire x_44649;
wire x_44650;
wire x_44651;
wire x_44652;
wire x_44653;
wire x_44654;
wire x_44655;
wire x_44656;
wire x_44657;
wire x_44658;
wire x_44659;
wire x_44660;
wire x_44661;
wire x_44662;
wire x_44663;
wire x_44664;
wire x_44665;
wire x_44666;
wire x_44667;
wire x_44668;
wire x_44669;
wire x_44670;
wire x_44671;
wire x_44672;
wire x_44673;
wire x_44674;
wire x_44675;
wire x_44676;
wire x_44677;
wire x_44678;
wire x_44679;
wire x_44680;
wire x_44681;
wire x_44682;
wire x_44683;
wire x_44684;
wire x_44685;
wire x_44686;
wire x_44687;
wire x_44688;
wire x_44689;
wire x_44690;
wire x_44691;
wire x_44692;
wire x_44693;
wire x_44694;
wire x_44695;
wire x_44696;
wire x_44697;
wire x_44698;
wire x_44699;
wire x_44700;
wire x_44701;
wire x_44702;
wire x_44703;
wire x_44704;
wire x_44705;
wire x_44706;
wire x_44707;
wire x_44708;
wire x_44709;
wire x_44710;
wire x_44711;
wire x_44712;
wire x_44713;
wire x_44714;
wire x_44715;
wire x_44716;
wire x_44717;
wire x_44718;
wire x_44719;
wire x_44720;
wire x_44721;
wire x_44722;
wire x_44723;
wire x_44724;
wire x_44725;
wire x_44726;
wire x_44727;
wire x_44728;
wire x_44729;
wire x_44730;
wire x_44731;
wire x_44732;
wire x_44733;
wire x_44734;
wire x_44735;
wire x_44736;
wire x_44737;
wire x_44738;
wire x_44739;
wire x_44740;
wire x_44741;
wire x_44742;
wire x_44743;
wire x_44744;
wire x_44745;
wire x_44746;
wire x_44747;
wire x_44748;
wire x_44749;
wire x_44750;
wire x_44751;
wire x_44752;
wire x_44753;
wire x_44754;
wire x_44755;
wire x_44756;
wire x_44757;
wire x_44758;
wire x_44759;
wire x_44760;
wire x_44761;
wire x_44762;
wire x_44763;
wire x_44764;
wire x_44765;
wire x_44766;
wire x_44767;
wire x_44768;
wire x_44769;
wire x_44770;
wire x_44771;
wire x_44772;
wire x_44773;
wire x_44774;
wire x_44775;
wire x_44776;
wire x_44777;
wire x_44778;
wire x_44779;
wire x_44780;
wire x_44781;
wire x_44782;
wire x_44783;
wire x_44784;
wire x_44785;
wire x_44786;
wire x_44787;
wire x_44788;
wire x_44789;
wire x_44790;
wire x_44791;
wire x_44792;
wire x_44793;
wire x_44794;
wire x_44795;
wire x_44796;
wire x_44797;
wire x_44798;
wire x_44799;
wire x_44800;
wire x_44801;
wire x_44802;
wire x_44803;
wire x_44804;
wire x_44805;
wire x_44806;
wire x_44807;
wire x_44808;
wire x_44809;
wire x_44810;
wire x_44811;
wire x_44812;
wire x_44813;
wire x_44814;
wire x_44815;
wire x_44816;
wire x_44817;
wire x_44818;
wire x_44819;
wire x_44820;
wire x_44821;
wire x_44822;
wire x_44823;
wire x_44824;
wire x_44825;
wire x_44826;
wire x_44827;
wire x_44828;
wire x_44829;
wire x_44830;
wire x_44831;
wire x_44832;
wire x_44833;
wire x_44834;
wire x_44835;
wire x_44836;
wire x_44837;
wire x_44838;
wire x_44839;
wire x_44840;
wire x_44841;
wire x_44842;
wire x_44843;
wire x_44844;
wire x_44845;
wire x_44846;
wire x_44847;
wire x_44848;
wire x_44849;
wire x_44850;
wire x_44851;
wire x_44852;
wire x_44853;
wire x_44854;
wire x_44855;
wire x_44856;
wire x_44857;
wire x_44858;
wire x_44859;
wire x_44860;
wire x_44861;
wire x_44862;
wire x_44863;
wire x_44864;
wire x_44865;
wire x_44866;
wire x_44867;
wire x_44868;
wire x_44869;
wire x_44870;
wire x_44871;
wire x_44872;
wire x_44873;
wire x_44874;
wire x_44875;
wire x_44876;
wire x_44877;
wire x_44878;
wire x_44879;
wire x_44880;
wire x_44881;
wire x_44882;
wire x_44883;
wire x_44884;
wire x_44885;
wire x_44886;
wire x_44887;
wire x_44888;
wire x_44889;
wire x_44890;
wire x_44891;
wire x_44892;
wire x_44893;
wire x_44894;
wire x_44895;
wire x_44896;
wire x_44897;
wire x_44898;
wire x_44899;
wire x_44900;
wire x_44901;
wire x_44902;
wire x_44903;
wire x_44904;
wire x_44905;
wire x_44906;
wire x_44907;
wire x_44908;
wire x_44909;
wire x_44910;
wire x_44911;
wire x_44912;
wire x_44913;
wire x_44914;
wire x_44915;
wire x_44916;
wire x_44917;
wire x_44918;
wire x_44919;
wire x_44920;
wire x_44921;
wire x_44922;
wire x_44923;
wire x_44924;
wire x_44925;
wire x_44926;
wire x_44927;
wire x_44928;
wire x_44929;
wire x_44930;
wire x_44931;
wire x_44932;
wire x_44933;
wire x_44934;
wire x_44935;
wire x_44936;
wire x_44937;
wire x_44938;
wire x_44939;
wire x_44940;
wire x_44941;
wire x_44942;
wire x_44943;
wire x_44944;
wire x_44945;
wire x_44946;
wire x_44947;
wire x_44948;
wire x_44949;
wire x_44950;
wire x_44951;
wire x_44952;
wire x_44953;
wire x_44954;
wire x_44955;
wire x_44956;
wire x_44957;
wire x_44958;
wire x_44959;
wire x_44960;
wire x_44961;
wire x_44962;
wire x_44963;
wire x_44964;
wire x_44965;
wire x_44966;
wire x_44967;
wire x_44968;
wire x_44969;
wire x_44970;
wire x_44971;
wire x_44972;
wire x_44973;
wire x_44974;
wire x_44975;
wire x_44976;
wire x_44977;
wire x_44978;
wire x_44979;
wire x_44980;
wire x_44981;
wire x_44982;
wire x_44983;
wire x_44984;
wire x_44985;
wire x_44986;
wire x_44987;
wire x_44988;
wire x_44989;
wire x_44990;
wire x_44991;
wire x_44992;
wire x_44993;
wire x_44994;
wire x_44995;
wire x_44996;
wire x_44997;
wire x_44998;
wire x_44999;
wire x_45000;
wire x_45001;
wire x_45002;
wire x_45003;
wire x_45004;
wire x_45005;
wire x_45006;
wire x_45007;
wire x_45008;
wire x_45009;
wire x_45010;
wire x_45011;
wire x_45012;
wire x_45013;
wire x_45014;
wire x_45015;
wire x_45016;
wire x_45017;
wire x_45018;
wire x_45019;
wire x_45020;
wire x_45021;
wire x_45022;
wire x_45023;
wire x_45024;
wire x_45025;
wire x_45026;
wire x_45027;
wire x_45028;
wire x_45029;
wire x_45030;
wire x_45031;
wire x_45032;
wire x_45033;
wire x_45034;
wire x_45035;
wire x_45036;
wire x_45037;
wire x_45038;
wire x_45039;
wire x_45040;
wire x_45041;
wire x_45042;
wire x_45043;
wire x_45044;
wire x_45045;
wire x_45046;
wire x_45047;
wire x_45048;
wire x_45049;
wire x_45050;
wire x_45051;
wire x_45052;
wire x_45053;
wire x_45054;
wire x_45055;
wire x_45056;
wire x_45057;
wire x_45058;
wire x_45059;
wire x_45060;
wire x_45061;
wire x_45062;
wire x_45063;
wire x_45064;
wire x_45065;
wire x_45066;
wire x_45067;
wire x_45068;
wire x_45069;
wire x_45070;
wire x_45071;
wire x_45072;
wire x_45073;
wire x_45074;
wire x_45075;
wire x_45076;
wire x_45077;
wire x_45078;
wire x_45079;
wire x_45080;
wire x_45081;
wire x_45082;
wire x_45083;
wire x_45084;
wire x_45085;
wire x_45086;
wire x_45087;
wire x_45088;
wire x_45089;
wire x_45090;
wire x_45091;
wire x_45092;
wire x_45093;
wire x_45094;
wire x_45095;
wire x_45096;
wire x_45097;
wire x_45098;
wire x_45099;
wire x_45100;
wire x_45101;
wire x_45102;
wire x_45103;
wire x_45104;
wire x_45105;
wire x_45106;
wire x_45107;
wire x_45108;
wire x_45109;
wire x_45110;
wire x_45111;
wire x_45112;
wire x_45113;
wire x_45114;
wire x_45115;
wire x_45116;
wire x_45117;
wire x_45118;
wire x_45119;
wire x_45120;
wire x_45121;
wire x_45122;
wire x_45123;
wire x_45124;
wire x_45125;
wire x_45126;
wire x_45127;
wire x_45128;
wire x_45129;
wire x_45130;
wire x_45131;
wire x_45132;
wire x_45133;
wire x_45134;
wire x_45135;
wire x_45136;
wire x_45137;
wire x_45138;
wire x_45139;
wire x_45140;
wire x_45141;
wire x_45142;
wire x_45143;
wire x_45144;
wire x_45145;
wire x_45146;
wire x_45147;
wire x_45148;
wire x_45149;
wire x_45150;
wire x_45151;
wire x_45152;
wire x_45153;
wire x_45154;
wire x_45155;
wire x_45156;
wire x_45157;
wire x_45158;
wire x_45159;
wire x_45160;
wire x_45161;
wire x_45162;
wire x_45163;
wire x_45164;
wire x_45165;
wire x_45166;
wire x_45167;
wire x_45168;
wire x_45169;
wire x_45170;
wire x_45171;
wire x_45172;
wire x_45173;
wire x_45174;
wire x_45175;
wire x_45176;
wire x_45177;
wire x_45178;
wire x_45179;
wire x_45180;
wire x_45181;
wire x_45182;
wire x_45183;
wire x_45184;
wire x_45185;
wire x_45186;
wire x_45187;
wire x_45188;
wire x_45189;
wire x_45190;
wire x_45191;
wire x_45192;
wire x_45193;
wire x_45194;
wire x_45195;
wire x_45196;
wire x_45197;
wire x_45198;
wire x_45199;
wire x_45200;
wire x_45201;
wire x_45202;
wire x_45203;
wire x_45204;
wire x_45205;
wire x_45206;
wire x_45207;
wire x_45208;
wire x_45209;
wire x_45210;
wire x_45211;
wire x_45212;
wire x_45213;
wire x_45214;
wire x_45215;
wire x_45216;
wire x_45217;
wire x_45218;
wire x_45219;
wire x_45220;
wire x_45221;
wire x_45222;
wire x_45223;
wire x_45224;
wire x_45225;
wire x_45226;
wire x_45227;
wire x_45228;
wire x_45229;
wire x_45230;
wire x_45231;
wire x_45232;
wire x_45233;
wire x_45234;
wire x_45235;
wire x_45236;
wire x_45237;
wire x_45238;
wire x_45239;
wire x_45240;
wire x_45241;
wire x_45242;
wire x_45243;
wire x_45244;
wire x_45245;
wire x_45246;
wire x_45247;
wire x_45248;
wire x_45249;
wire x_45250;
wire x_45251;
wire x_45252;
wire x_45253;
wire x_45254;
wire x_45255;
wire x_45256;
wire x_45257;
wire x_45258;
wire x_45259;
wire x_45260;
wire x_45261;
wire x_45262;
wire x_45263;
wire x_45264;
wire x_45265;
wire x_45266;
wire x_45267;
wire x_45268;
wire x_45269;
wire x_45270;
wire x_45271;
wire x_45272;
wire x_45273;
wire x_45274;
wire x_45275;
wire x_45276;
wire x_45277;
wire x_45278;
wire x_45279;
wire x_45280;
wire x_45281;
wire x_45282;
wire x_45283;
wire x_45284;
wire x_45285;
wire x_45286;
wire x_45287;
wire x_45288;
wire x_45289;
wire x_45290;
wire x_45291;
wire x_45292;
wire x_45293;
wire x_45294;
wire x_45295;
wire x_45296;
wire x_45297;
wire x_45298;
wire x_45299;
wire x_45300;
wire x_45301;
wire x_45302;
wire x_45303;
wire x_45304;
wire x_45305;
wire x_45306;
wire x_45307;
wire x_45308;
wire x_45309;
wire x_45310;
wire x_45311;
wire x_45312;
wire x_45313;
wire x_45314;
wire x_45315;
wire x_45316;
wire x_45317;
wire x_45318;
wire x_45319;
wire x_45320;
wire x_45321;
wire x_45322;
wire x_45323;
wire x_45324;
wire x_45325;
wire x_45326;
wire x_45327;
wire x_45328;
wire x_45329;
wire x_45330;
wire x_45331;
wire x_45332;
wire x_45333;
wire x_45334;
wire x_45335;
wire x_45336;
wire x_45337;
wire x_45338;
wire x_45339;
wire x_45340;
wire x_45341;
wire x_45342;
wire x_45343;
wire x_45344;
wire x_45345;
wire x_45346;
wire x_45347;
wire x_45348;
wire x_45349;
wire x_45350;
wire x_45351;
wire x_45352;
wire x_45353;
wire x_45354;
wire x_45355;
wire x_45356;
wire x_45357;
wire x_45358;
wire x_45359;
wire x_45360;
wire x_45361;
wire x_45362;
wire x_45363;
wire x_45364;
wire x_45365;
wire x_45366;
wire x_45367;
wire x_45368;
wire x_45369;
wire x_45370;
wire x_45371;
wire x_45372;
wire x_45373;
wire x_45374;
wire x_45375;
wire x_45376;
wire x_45377;
wire x_45378;
wire x_45379;
wire x_45380;
wire x_45381;
wire x_45382;
wire x_45383;
wire x_45384;
wire x_45385;
wire x_45386;
wire x_45387;
wire x_45388;
wire x_45389;
wire x_45390;
wire x_45391;
wire x_45392;
wire x_45393;
wire x_45394;
wire x_45395;
wire x_45396;
wire x_45397;
wire x_45398;
wire x_45399;
wire x_45400;
wire x_45401;
wire x_45402;
wire x_45403;
wire x_45404;
wire x_45405;
wire x_45406;
wire x_45407;
wire x_45408;
wire x_45409;
wire x_45410;
wire x_45411;
wire x_45412;
wire x_45413;
wire x_45414;
wire x_45415;
wire x_45416;
wire x_45417;
wire x_45418;
wire x_45419;
wire x_45420;
wire x_45421;
wire x_45422;
wire x_45423;
wire x_45424;
wire x_45425;
wire x_45426;
wire x_45427;
wire x_45428;
wire x_45429;
wire x_45430;
wire x_45431;
wire x_45432;
wire x_45433;
wire x_45434;
wire x_45435;
wire x_45436;
wire x_45437;
wire x_45438;
wire x_45439;
wire x_45440;
wire x_45441;
wire x_45442;
wire x_45443;
wire x_45444;
wire x_45445;
wire x_45446;
wire x_45447;
wire x_45448;
wire x_45449;
wire x_45450;
wire x_45451;
wire x_45452;
wire x_45453;
wire x_45454;
wire x_45455;
wire x_45456;
wire x_45457;
wire x_45458;
wire x_45459;
wire x_45460;
wire x_45461;
wire x_45462;
wire x_45463;
wire x_45464;
wire x_45465;
wire x_45466;
wire x_45467;
wire x_45468;
wire x_45469;
wire x_45470;
wire x_45471;
wire x_45472;
wire x_45473;
wire x_45474;
wire x_45475;
wire x_45476;
wire x_45477;
wire x_45478;
wire x_45479;
wire x_45480;
wire x_45481;
wire x_45482;
wire x_45483;
wire x_45484;
wire x_45485;
wire x_45486;
wire x_45487;
wire x_45488;
wire x_45489;
wire x_45490;
wire x_45491;
wire x_45492;
wire x_45493;
wire x_45494;
wire x_45495;
wire x_45496;
wire x_45497;
wire x_45498;
wire x_45499;
wire x_45500;
wire x_45501;
wire x_45502;
wire x_45503;
wire x_45504;
wire x_45505;
wire x_45506;
wire x_45507;
wire x_45508;
wire x_45509;
wire x_45510;
wire x_45511;
wire x_45512;
wire x_45513;
wire x_45514;
wire x_45515;
wire x_45516;
wire x_45517;
wire x_45518;
wire x_45519;
wire x_45520;
wire x_45521;
wire x_45522;
wire x_45523;
wire x_45524;
wire x_45525;
wire x_45526;
wire x_45527;
wire x_45528;
wire x_45529;
wire x_45530;
wire x_45531;
wire x_45532;
wire x_45533;
wire x_45534;
wire x_45535;
wire x_45536;
wire x_45537;
wire x_45538;
wire x_45539;
wire x_45540;
wire x_45541;
wire x_45542;
wire x_45543;
wire x_45544;
wire x_45545;
wire x_45546;
wire x_45547;
wire x_45548;
wire x_45549;
wire x_45550;
wire x_45551;
wire x_45552;
wire x_45553;
wire x_45554;
wire x_45555;
wire x_45556;
wire x_45557;
wire x_45558;
wire x_45559;
wire x_45560;
wire x_45561;
wire x_45562;
wire x_45563;
wire x_45564;
wire x_45565;
wire x_45566;
wire x_45567;
wire x_45568;
wire x_45569;
wire x_45570;
wire x_45571;
wire x_45572;
wire x_45573;
wire x_45574;
wire x_45575;
wire x_45576;
wire x_45577;
wire x_45578;
wire x_45579;
wire x_45580;
wire x_45581;
wire x_45582;
wire x_45583;
wire x_45584;
wire x_45585;
wire x_45586;
wire x_45587;
wire x_45588;
wire x_45589;
wire x_45590;
wire x_45591;
wire x_45592;
wire x_45593;
wire x_45594;
wire x_45595;
wire x_45596;
wire x_45597;
wire x_45598;
wire x_45599;
wire x_45600;
wire x_45601;
wire x_45602;
wire x_45603;
wire x_45604;
wire x_45605;
wire x_45606;
wire x_45607;
wire x_45608;
wire x_45609;
wire x_45610;
wire x_45611;
wire x_45612;
wire x_45613;
wire x_45614;
wire x_45615;
wire x_45616;
wire x_45617;
wire x_45618;
wire x_45619;
wire x_45620;
wire x_45621;
wire x_45622;
wire x_45623;
wire x_45624;
wire x_45625;
wire x_45626;
wire x_45627;
wire x_45628;
wire x_45629;
wire x_45630;
wire x_45631;
wire x_45632;
wire x_45633;
wire x_45634;
wire x_45635;
wire x_45636;
wire x_45637;
wire x_45638;
wire x_45639;
wire x_45640;
wire x_45641;
wire x_45642;
wire x_45643;
wire x_45644;
wire x_45645;
wire x_45646;
wire x_45647;
wire x_45648;
wire x_45649;
wire x_45650;
wire x_45651;
wire x_45652;
wire x_45653;
wire x_45654;
wire x_45655;
wire x_45656;
wire x_45657;
wire x_45658;
wire x_45659;
wire x_45660;
wire x_45661;
wire x_45662;
wire x_45663;
wire x_45664;
wire x_45665;
wire x_45666;
wire x_45667;
wire x_45668;
wire x_45669;
wire x_45670;
wire x_45671;
wire x_45672;
wire x_45673;
wire x_45674;
wire x_45675;
wire x_45676;
wire x_45677;
wire x_45678;
wire x_45679;
wire x_45680;
wire x_45681;
wire x_45682;
wire x_45683;
wire x_45684;
wire x_45685;
wire x_45686;
wire x_45687;
wire x_45688;
wire x_45689;
wire x_45690;
wire x_45691;
wire x_45692;
wire x_45693;
wire x_45694;
wire x_45695;
wire x_45696;
wire x_45697;
wire x_45698;
wire x_45699;
wire x_45700;
wire x_45701;
wire x_45702;
wire x_45703;
wire x_45704;
wire x_45705;
wire x_45706;
wire x_45707;
wire x_45708;
wire x_45709;
wire x_45710;
wire x_45711;
wire x_45712;
wire x_45713;
wire x_45714;
wire x_45715;
wire x_45716;
wire x_45717;
wire x_45718;
wire x_45719;
wire x_45720;
wire x_45721;
wire x_45722;
wire x_45723;
wire x_45724;
wire x_45725;
wire x_45726;
wire x_45727;
wire x_45728;
wire x_45729;
wire x_45730;
wire x_45731;
wire x_45732;
wire x_45733;
wire x_45734;
wire x_45735;
wire x_45736;
wire x_45737;
wire x_45738;
wire x_45739;
wire x_45740;
wire x_45741;
wire x_45742;
wire x_45743;
wire x_45744;
wire x_45745;
wire x_45746;
wire x_45747;
wire x_45748;
wire x_45749;
wire x_45750;
wire x_45751;
wire x_45752;
wire x_45753;
wire x_45754;
wire x_45755;
wire x_45756;
wire x_45757;
wire x_45758;
wire x_45759;
wire x_45760;
wire x_45761;
wire x_45762;
wire x_45763;
wire x_45764;
wire x_45765;
wire x_45766;
wire x_45767;
wire x_45768;
wire x_45769;
wire x_45770;
wire x_45771;
wire x_45772;
wire x_45773;
wire x_45774;
wire x_45775;
wire x_45776;
wire x_45777;
wire x_45778;
wire x_45779;
wire x_45780;
wire x_45781;
wire x_45782;
wire x_45783;
wire x_45784;
wire x_45785;
wire x_45786;
wire x_45787;
wire x_45788;
wire x_45789;
wire x_45790;
wire x_45791;
wire x_45792;
wire x_45793;
wire x_45794;
wire x_45795;
wire x_45796;
wire x_45797;
wire x_45798;
wire x_45799;
wire x_45800;
wire x_45801;
wire x_45802;
wire x_45803;
wire x_45804;
wire x_45805;
wire x_45806;
wire x_45807;
wire x_45808;
wire x_45809;
wire x_45810;
wire x_45811;
wire x_45812;
wire x_45813;
wire x_45814;
wire x_45815;
wire x_45816;
wire x_45817;
wire x_45818;
wire x_45819;
wire x_45820;
wire x_45821;
wire x_45822;
wire x_45823;
wire x_45824;
wire x_45825;
wire x_45826;
wire x_45827;
wire x_45828;
wire x_45829;
wire x_45830;
wire x_45831;
wire x_45832;
wire x_45833;
wire x_45834;
wire x_45835;
wire x_45836;
wire x_45837;
wire x_45838;
wire x_45839;
wire x_45840;
wire x_45841;
wire x_45842;
wire x_45843;
wire x_45844;
wire x_45845;
wire x_45846;
wire x_45847;
wire x_45848;
wire x_45849;
wire x_45850;
wire x_45851;
wire x_45852;
wire x_45853;
wire x_45854;
wire x_45855;
wire x_45856;
wire x_45857;
wire x_45858;
wire x_45859;
wire x_45860;
wire x_45861;
wire x_45862;
wire x_45863;
wire x_45864;
wire x_45865;
wire x_45866;
wire x_45867;
wire x_45868;
wire x_45869;
wire x_45870;
wire x_45871;
wire x_45872;
wire x_45873;
wire x_45874;
wire x_45875;
wire x_45876;
wire x_45877;
wire x_45878;
wire x_45879;
wire x_45880;
wire x_45881;
wire x_45882;
wire x_45883;
wire x_45884;
wire x_45885;
wire x_45886;
wire x_45887;
wire x_45888;
wire x_45889;
wire x_45890;
wire x_45891;
wire x_45892;
wire x_45893;
wire x_45894;
wire x_45895;
wire x_45896;
wire x_45897;
wire x_45898;
wire x_45899;
wire x_45900;
wire x_45901;
wire x_45902;
wire x_45903;
wire x_45904;
wire x_45905;
wire x_45906;
wire x_45907;
wire x_45908;
wire x_45909;
wire x_45910;
wire x_45911;
wire x_45912;
wire x_45913;
wire x_45914;
wire x_45915;
wire x_45916;
wire x_45917;
wire x_45918;
wire x_45919;
wire x_45920;
wire x_45921;
wire x_45922;
wire x_45923;
wire x_45924;
wire x_45925;
wire x_45926;
wire x_45927;
wire x_45928;
wire x_45929;
wire x_45930;
wire x_45931;
wire x_45932;
wire x_45933;
wire x_45934;
wire x_45935;
wire x_45936;
wire x_45937;
wire x_45938;
wire x_45939;
wire x_45940;
wire x_45941;
wire x_45942;
wire x_45943;
wire x_45944;
wire x_45945;
wire x_45946;
wire x_45947;
wire x_45948;
wire x_45949;
wire x_45950;
wire x_45951;
wire x_45952;
wire x_45953;
wire x_45954;
wire x_45955;
wire x_45956;
wire x_45957;
wire x_45958;
wire x_45959;
wire x_45960;
wire x_45961;
wire x_45962;
wire x_45963;
wire x_45964;
wire x_45965;
wire x_45966;
wire x_45967;
wire x_45968;
wire x_45969;
wire x_45970;
wire x_45971;
wire x_45972;
wire x_45973;
wire x_45974;
wire x_45975;
wire x_45976;
wire x_45977;
wire x_45978;
wire x_45979;
wire x_45980;
wire x_45981;
wire x_45982;
wire x_45983;
wire x_45984;
wire x_45985;
wire x_45986;
wire x_45987;
wire x_45988;
wire x_45989;
wire x_45990;
wire x_45991;
wire x_45992;
wire x_45993;
wire x_45994;
wire x_45995;
wire x_45996;
wire x_45997;
wire x_45998;
wire x_45999;
wire x_46000;
wire x_46001;
wire x_46002;
wire x_46003;
wire x_46004;
wire x_46005;
wire x_46006;
wire x_46007;
wire x_46008;
wire x_46009;
wire x_46010;
wire x_46011;
wire x_46012;
wire x_46013;
wire x_46014;
wire x_46015;
wire x_46016;
wire x_46017;
wire x_46018;
wire x_46019;
wire x_46020;
wire x_46021;
wire x_46022;
wire x_46023;
wire x_46024;
wire x_46025;
wire x_46026;
wire x_46027;
wire x_46028;
wire x_46029;
wire x_46030;
wire x_46031;
wire x_46032;
wire x_46033;
wire x_46034;
wire x_46035;
wire x_46036;
wire x_46037;
wire x_46038;
wire x_46039;
wire x_46040;
wire x_46041;
wire x_46042;
wire x_46043;
wire x_46044;
wire x_46045;
wire x_46046;
wire x_46047;
wire x_46048;
wire x_46049;
wire x_46050;
wire x_46051;
wire x_46052;
wire x_46053;
wire x_46054;
wire x_46055;
wire x_46056;
wire x_46057;
wire x_46058;
wire x_46059;
wire x_46060;
wire x_46061;
wire x_46062;
wire x_46063;
wire x_46064;
wire x_46065;
wire x_46066;
wire x_46067;
wire x_46068;
wire x_46069;
wire x_46070;
wire x_46071;
wire x_46072;
wire x_46073;
wire x_46074;
wire x_46075;
wire x_46076;
wire x_46077;
wire x_46078;
wire x_46079;
wire x_46080;
wire x_46081;
wire x_46082;
wire x_46083;
wire x_46084;
wire x_46085;
wire x_46086;
wire x_46087;
wire x_46088;
wire x_46089;
wire x_46090;
wire x_46091;
wire x_46092;
wire x_46093;
wire x_46094;
wire x_46095;
wire x_46096;
wire x_46097;
wire x_46098;
wire x_46099;
wire x_46100;
wire x_46101;
wire x_46102;
wire x_46103;
wire x_46104;
wire x_46105;
wire x_46106;
wire x_46107;
wire x_46108;
wire x_46109;
wire x_46110;
wire x_46111;
wire x_46112;
wire x_46113;
wire x_46114;
wire x_46115;
wire x_46116;
wire x_46117;
wire x_46118;
wire x_46119;
wire x_46120;
wire x_46121;
wire x_46122;
wire x_46123;
wire x_46124;
wire x_46125;
wire x_46126;
wire x_46127;
wire x_46128;
wire x_46129;
wire x_46130;
wire x_46131;
wire x_46132;
wire x_46133;
wire x_46134;
wire x_46135;
wire x_46136;
wire x_46137;
wire x_46138;
wire x_46139;
wire x_46140;
wire x_46141;
wire x_46142;
wire x_46143;
wire x_46144;
wire x_46145;
wire x_46146;
wire x_46147;
wire x_46148;
wire x_46149;
wire x_46150;
wire x_46151;
wire x_46152;
wire x_46153;
wire x_46154;
wire x_46155;
wire x_46156;
wire x_46157;
wire x_46158;
wire x_46159;
wire x_46160;
wire x_46161;
wire x_46162;
wire x_46163;
wire x_46164;
wire x_46165;
wire x_46166;
wire x_46167;
wire x_46168;
wire x_46169;
wire x_46170;
wire x_46171;
wire x_46172;
wire x_46173;
wire x_46174;
wire x_46175;
wire x_46176;
wire x_46177;
wire x_46178;
wire x_46179;
wire x_46180;
wire x_46181;
wire x_46182;
wire x_46183;
wire x_46184;
wire x_46185;
wire x_46186;
wire x_46187;
wire x_46188;
wire x_46189;
wire x_46190;
wire x_46191;
wire x_46192;
wire x_46193;
wire x_46194;
wire x_46195;
wire x_46196;
wire x_46197;
wire x_46198;
wire x_46199;
wire x_46200;
wire x_46201;
wire x_46202;
wire x_46203;
wire x_46204;
wire x_46205;
wire x_46206;
wire x_46207;
wire x_46208;
wire x_46209;
wire x_46210;
wire x_46211;
wire x_46212;
wire x_46213;
wire x_46214;
wire x_46215;
wire x_46216;
wire x_46217;
wire x_46218;
wire x_46219;
wire x_46220;
wire x_46221;
wire x_46222;
wire x_46223;
wire x_46224;
wire x_46225;
wire x_46226;
wire x_46227;
wire x_46228;
wire x_46229;
wire x_46230;
wire x_46231;
wire x_46232;
wire x_46233;
wire x_46234;
wire x_46235;
wire x_46236;
wire x_46237;
wire x_46238;
wire x_46239;
wire x_46240;
wire x_46241;
wire x_46242;
wire x_46243;
wire x_46244;
wire x_46245;
wire x_46246;
wire x_46247;
wire x_46248;
wire x_46249;
wire x_46250;
wire x_46251;
wire x_46252;
wire x_46253;
wire x_46254;
wire x_46255;
wire x_46256;
wire x_46257;
wire x_46258;
wire x_46259;
wire x_46260;
wire x_46261;
wire x_46262;
wire x_46263;
wire x_46264;
wire x_46265;
wire x_46266;
wire x_46267;
wire x_46268;
wire x_46269;
wire x_46270;
wire x_46271;
wire x_46272;
wire x_46273;
wire x_46274;
wire x_46275;
wire x_46276;
wire x_46277;
wire x_46278;
wire x_46279;
wire x_46280;
wire x_46281;
wire x_46282;
wire x_46283;
wire x_46284;
wire x_46285;
wire x_46286;
wire x_46287;
wire x_46288;
wire x_46289;
wire x_46290;
wire x_46291;
wire x_46292;
wire x_46293;
wire x_46294;
wire x_46295;
wire x_46296;
wire x_46297;
wire x_46298;
wire x_46299;
wire x_46300;
wire x_46301;
wire x_46302;
wire x_46303;
wire x_46304;
wire x_46305;
wire x_46306;
wire x_46307;
wire x_46308;
wire x_46309;
wire x_46310;
wire x_46311;
wire x_46312;
wire x_46313;
wire x_46314;
wire x_46315;
wire x_46316;
wire x_46317;
wire x_46318;
wire x_46319;
wire x_46320;
wire x_46321;
wire x_46322;
wire x_46323;
wire x_46324;
wire x_46325;
wire x_46326;
wire x_46327;
wire x_46328;
wire x_46329;
wire x_46330;
wire x_46331;
wire x_46332;
wire x_46333;
wire x_46334;
wire x_46335;
wire x_46336;
wire x_46337;
wire x_46338;
wire x_46339;
wire x_46340;
wire x_46341;
wire x_46342;
wire x_46343;
wire x_46344;
wire x_46345;
wire x_46346;
wire x_46347;
wire x_46348;
wire x_46349;
wire x_46350;
wire x_46351;
wire x_46352;
wire x_46353;
wire x_46354;
wire x_46355;
wire x_46356;
wire x_46357;
wire x_46358;
wire x_46359;
wire x_46360;
wire x_46361;
wire x_46362;
wire x_46363;
wire x_46364;
wire x_46365;
wire x_46366;
wire x_46367;
wire x_46368;
wire x_46369;
wire x_46370;
wire x_46371;
wire x_46372;
wire x_46373;
wire x_46374;
wire x_46375;
wire x_46376;
wire x_46377;
wire x_46378;
wire x_46379;
wire x_46380;
wire x_46381;
wire x_46382;
wire x_46383;
wire x_46384;
wire x_46385;
wire x_46386;
wire x_46387;
wire x_46388;
wire x_46389;
wire x_46390;
wire x_46391;
wire x_46392;
wire x_46393;
wire x_46394;
wire x_46395;
wire x_46396;
wire x_46397;
wire x_46398;
wire x_46399;
wire x_46400;
wire x_46401;
wire x_46402;
wire x_46403;
wire x_46404;
wire x_46405;
wire x_46406;
wire x_46407;
wire x_46408;
wire x_46409;
wire x_46410;
wire x_46411;
wire x_46412;
wire x_46413;
wire x_46414;
wire x_46415;
wire x_46416;
wire x_46417;
wire x_46418;
wire x_46419;
wire x_46420;
wire x_46421;
wire x_46422;
wire x_46423;
wire x_46424;
wire x_46425;
wire x_46426;
wire x_46427;
wire x_46428;
wire x_46429;
wire x_46430;
wire x_46431;
wire x_46432;
wire x_46433;
wire x_46434;
wire x_46435;
wire x_46436;
wire x_46437;
wire x_46438;
wire x_46439;
wire x_46440;
wire x_46441;
wire x_46442;
wire x_46443;
wire x_46444;
wire x_46445;
wire x_46446;
wire x_46447;
wire x_46448;
wire x_46449;
wire x_46450;
wire x_46451;
wire x_46452;
wire x_46453;
wire x_46454;
wire x_46455;
wire x_46456;
wire x_46457;
wire x_46458;
wire x_46459;
wire x_46460;
wire x_46461;
wire x_46462;
wire x_46463;
wire x_46464;
wire x_46465;
wire x_46466;
wire x_46467;
wire x_46468;
wire x_46469;
wire x_46470;
wire x_46471;
wire x_46472;
wire x_46473;
wire x_46474;
wire x_46475;
wire x_46476;
wire x_46477;
wire x_46478;
wire x_46479;
wire x_46480;
wire x_46481;
wire x_46482;
wire x_46483;
wire x_46484;
wire x_46485;
wire x_46486;
wire x_46487;
wire x_46488;
wire x_46489;
wire x_46490;
wire x_46491;
wire x_46492;
wire x_46493;
wire x_46494;
wire x_46495;
wire x_46496;
wire x_46497;
wire x_46498;
wire x_46499;
wire x_46500;
wire x_46501;
wire x_46502;
wire x_46503;
wire x_46504;
wire x_46505;
wire x_46506;
wire x_46507;
wire x_46508;
wire x_46509;
wire x_46510;
wire x_46511;
wire x_46512;
wire x_46513;
wire x_46514;
wire x_46515;
wire x_46516;
wire x_46517;
wire x_46518;
wire x_46519;
wire x_46520;
wire x_46521;
wire x_46522;
wire x_46523;
wire x_46524;
wire x_46525;
wire x_46526;
wire x_46527;
wire x_46528;
wire x_46529;
wire x_46530;
wire x_46531;
wire x_46532;
wire x_46533;
wire x_46534;
wire x_46535;
wire x_46536;
wire x_46537;
wire x_46538;
wire x_46539;
wire x_46540;
wire x_46541;
wire x_46542;
wire x_46543;
wire x_46544;
wire x_46545;
wire x_46546;
wire x_46547;
wire x_46548;
wire x_46549;
wire x_46550;
wire x_46551;
wire x_46552;
wire x_46553;
wire x_46554;
wire x_46555;
wire x_46556;
wire x_46557;
wire x_46558;
wire x_46559;
wire x_46560;
wire x_46561;
wire x_46562;
wire x_46563;
wire x_46564;
wire x_46565;
wire x_46566;
wire x_46567;
wire x_46568;
wire x_46569;
wire x_46570;
wire x_46571;
wire x_46572;
wire x_46573;
wire x_46574;
wire x_46575;
wire x_46576;
wire x_46577;
wire x_46578;
wire x_46579;
wire x_46580;
wire x_46581;
wire x_46582;
wire x_46583;
wire x_46584;
wire x_46585;
wire x_46586;
wire x_46587;
wire x_46588;
wire x_46589;
wire x_46590;
wire x_46591;
wire x_46592;
wire x_46593;
wire x_46594;
wire x_46595;
wire x_46596;
wire x_46597;
wire x_46598;
wire x_46599;
wire x_46600;
wire x_46601;
wire x_46602;
wire x_46603;
wire x_46604;
wire x_46605;
wire x_46606;
wire x_46607;
wire x_46608;
wire x_46609;
wire x_46610;
wire x_46611;
wire x_46612;
wire x_46613;
wire x_46614;
wire x_46615;
wire x_46616;
wire x_46617;
wire x_46618;
wire x_46619;
wire x_46620;
wire x_46621;
wire x_46622;
wire x_46623;
wire x_46624;
wire x_46625;
wire x_46626;
wire x_46627;
wire x_46628;
wire x_46629;
wire x_46630;
wire x_46631;
wire x_46632;
wire x_46633;
wire x_46634;
wire x_46635;
wire x_46636;
wire x_46637;
wire x_46638;
wire x_46639;
wire x_46640;
wire x_46641;
wire x_46642;
wire x_46643;
wire x_46644;
wire x_46645;
wire x_46646;
wire x_46647;
wire x_46648;
wire x_46649;
wire x_46650;
wire x_46651;
wire x_46652;
wire x_46653;
wire x_46654;
wire x_46655;
wire x_46656;
wire x_46657;
wire x_46658;
wire x_46659;
wire x_46660;
wire x_46661;
wire x_46662;
wire x_46663;
wire x_46664;
wire x_46665;
wire x_46666;
wire x_46667;
wire x_46668;
wire x_46669;
wire x_46670;
wire x_46671;
wire x_46672;
wire x_46673;
wire x_46674;
wire x_46675;
wire x_46676;
wire x_46677;
wire x_46678;
wire x_46679;
wire x_46680;
wire x_46681;
wire x_46682;
wire x_46683;
wire x_46684;
wire x_46685;
wire x_46686;
wire x_46687;
wire x_46688;
wire x_46689;
wire x_46690;
wire x_46691;
wire x_46692;
wire x_46693;
wire x_46694;
wire x_46695;
wire x_46696;
wire x_46697;
wire x_46698;
wire x_46699;
wire x_46700;
wire x_46701;
wire x_46702;
wire x_46703;
wire x_46704;
wire x_46705;
wire x_46706;
wire x_46707;
wire x_46708;
wire x_46709;
wire x_46710;
wire x_46711;
wire x_46712;
wire x_46713;
wire x_46714;
wire x_46715;
wire x_46716;
wire x_46717;
wire x_46718;
wire x_46719;
wire x_46720;
wire x_46721;
wire x_46722;
wire x_46723;
wire x_46724;
wire x_46725;
wire x_46726;
wire x_46727;
wire x_46728;
wire x_46729;
wire x_46730;
wire x_46731;
wire x_46732;
wire x_46733;
wire x_46734;
wire x_46735;
wire x_46736;
wire x_46737;
wire x_46738;
wire x_46739;
wire x_46740;
wire x_46741;
wire x_46742;
wire x_46743;
wire x_46744;
wire x_46745;
wire x_46746;
wire x_46747;
wire x_46748;
wire x_46749;
wire x_46750;
wire x_46751;
wire x_46752;
wire x_46753;
wire x_46754;
wire x_46755;
wire x_46756;
wire x_46757;
wire x_46758;
wire x_46759;
wire x_46760;
wire x_46761;
wire x_46762;
wire x_46763;
wire x_46764;
wire x_46765;
wire x_46766;
wire x_46767;
wire x_46768;
wire x_46769;
wire x_46770;
wire x_46771;
wire x_46772;
wire x_46773;
wire x_46774;
wire x_46775;
wire x_46776;
wire x_46777;
wire x_46778;
wire x_46779;
wire x_46780;
wire x_46781;
wire x_46782;
wire x_46783;
wire x_46784;
wire x_46785;
wire x_46786;
wire x_46787;
wire x_46788;
wire x_46789;
wire x_46790;
wire x_46791;
wire x_46792;
wire x_46793;
wire x_46794;
wire x_46795;
wire x_46796;
wire x_46797;
wire x_46798;
wire x_46799;
wire x_46800;
wire x_46801;
wire x_46802;
wire x_46803;
wire x_46804;
wire x_46805;
wire x_46806;
wire x_46807;
wire x_46808;
wire x_46809;
wire x_46810;
wire x_46811;
wire x_46812;
wire x_46813;
wire x_46814;
wire x_46815;
wire x_46816;
wire x_46817;
wire x_46818;
wire x_46819;
wire x_46820;
wire x_46821;
wire x_46822;
wire x_46823;
wire x_46824;
wire x_46825;
wire x_46826;
wire x_46827;
wire x_46828;
wire x_46829;
wire x_46830;
wire x_46831;
wire x_46832;
wire x_46833;
wire x_46834;
wire x_46835;
wire x_46836;
wire x_46837;
wire x_46838;
wire x_46839;
wire x_46840;
wire x_46841;
wire x_46842;
wire x_46843;
wire x_46844;
wire x_46845;
wire x_46846;
wire x_46847;
wire x_46848;
wire x_46849;
wire x_46850;
wire x_46851;
wire x_46852;
wire x_46853;
wire x_46854;
wire x_46855;
wire x_46856;
wire x_46857;
wire x_46858;
wire x_46859;
wire x_46860;
wire x_46861;
wire x_46862;
wire x_46863;
wire x_46864;
wire x_46865;
wire x_46866;
wire x_46867;
wire x_46868;
wire x_46869;
wire x_46870;
wire x_46871;
wire x_46872;
wire x_46873;
wire x_46874;
wire x_46875;
wire x_46876;
wire x_46877;
wire x_46878;
wire x_46879;
wire x_46880;
wire x_46881;
wire x_46882;
wire x_46883;
wire x_46884;
wire x_46885;
wire x_46886;
wire x_46887;
wire x_46888;
wire x_46889;
wire x_46890;
wire x_46891;
wire x_46892;
wire x_46893;
wire x_46894;
wire x_46895;
wire x_46896;
wire x_46897;
wire x_46898;
wire x_46899;
wire x_46900;
wire x_46901;
wire x_46902;
wire x_46903;
wire x_46904;
wire x_46905;
wire x_46906;
wire x_46907;
wire x_46908;
wire x_46909;
wire x_46910;
wire x_46911;
wire x_46912;
wire x_46913;
wire x_46914;
wire x_46915;
wire x_46916;
wire x_46917;
wire x_46918;
wire x_46919;
wire x_46920;
wire x_46921;
wire x_46922;
wire x_46923;
wire x_46924;
wire x_46925;
wire x_46926;
wire x_46927;
wire x_46928;
wire x_46929;
wire x_46930;
wire x_46931;
wire x_46932;
wire x_46933;
wire x_46934;
wire x_46935;
wire x_46936;
wire x_46937;
wire x_46938;
wire x_46939;
wire x_46940;
wire x_46941;
wire x_46942;
wire x_46943;
wire x_46944;
wire x_46945;
wire x_46946;
wire x_46947;
wire x_46948;
wire x_46949;
wire x_46950;
wire x_46951;
wire x_46952;
wire x_46953;
wire x_46954;
wire x_46955;
wire x_46956;
wire x_46957;
wire x_46958;
wire x_46959;
wire x_46960;
wire x_46961;
wire x_46962;
wire x_46963;
wire x_46964;
wire x_46965;
wire x_46966;
wire x_46967;
wire x_46968;
wire x_46969;
wire x_46970;
wire x_46971;
wire x_46972;
wire x_46973;
wire x_46974;
wire x_46975;
wire x_46976;
wire x_46977;
wire x_46978;
wire x_46979;
wire x_46980;
wire x_46981;
wire x_46982;
wire x_46983;
wire x_46984;
wire x_46985;
wire x_46986;
wire x_46987;
wire x_46988;
wire x_46989;
wire x_46990;
wire x_46991;
wire x_46992;
wire x_46993;
wire x_46994;
wire x_46995;
wire x_46996;
wire x_46997;
wire x_46998;
wire x_46999;
wire x_47000;
wire x_47001;
wire x_47002;
wire x_47003;
wire x_47004;
wire x_47005;
wire x_47006;
wire x_47007;
wire x_47008;
wire x_47009;
wire x_47010;
wire x_47011;
wire x_47012;
wire x_47013;
wire x_47014;
wire x_47015;
wire x_47016;
wire x_47017;
wire x_47018;
wire x_47019;
wire x_47020;
wire x_47021;
wire x_47022;
wire x_47023;
wire x_47024;
wire x_47025;
wire x_47026;
wire x_47027;
wire x_47028;
wire x_47029;
wire x_47030;
wire x_47031;
wire x_47032;
wire x_47033;
wire x_47034;
wire x_47035;
wire x_47036;
wire x_47037;
wire x_47038;
wire x_47039;
wire x_47040;
wire x_47041;
wire x_47042;
wire x_47043;
wire x_47044;
wire x_47045;
wire x_47046;
wire x_47047;
wire x_47048;
wire x_47049;
wire x_47050;
wire x_47051;
wire x_47052;
wire x_47053;
wire x_47054;
wire x_47055;
wire x_47056;
wire x_47057;
wire x_47058;
wire x_47059;
wire x_47060;
wire x_47061;
wire x_47062;
wire x_47063;
wire x_47064;
wire x_47065;
wire x_47066;
wire x_47067;
wire x_47068;
wire x_47069;
wire x_47070;
wire x_47071;
wire x_47072;
wire x_47073;
wire x_47074;
wire x_47075;
wire x_47076;
wire x_47077;
wire x_47078;
wire x_47079;
wire x_47080;
wire x_47081;
wire x_47082;
wire x_47083;
wire x_47084;
wire x_47085;
wire x_47086;
wire x_47087;
wire x_47088;
wire x_47089;
wire x_47090;
wire x_47091;
wire x_47092;
wire x_47093;
wire x_47094;
wire x_47095;
wire x_47096;
wire x_47097;
wire x_47098;
wire x_47099;
wire x_47100;
wire x_47101;
wire x_47102;
wire x_47103;
wire x_47104;
wire x_47105;
wire x_47106;
wire x_47107;
wire x_47108;
wire x_47109;
wire x_47110;
wire x_47111;
wire x_47112;
wire x_47113;
wire x_47114;
wire x_47115;
wire x_47116;
wire x_47117;
wire x_47118;
wire x_47119;
wire x_47120;
wire x_47121;
wire x_47122;
wire x_47123;
wire x_47124;
wire x_47125;
wire x_47126;
wire x_47127;
wire x_47128;
wire x_47129;
wire x_47130;
wire x_47131;
wire x_47132;
wire x_47133;
wire x_47134;
wire x_47135;
wire x_47136;
wire x_47137;
wire x_47138;
wire x_47139;
wire x_47140;
wire x_47141;
wire x_47142;
wire x_47143;
wire x_47144;
wire x_47145;
wire x_47146;
wire x_47147;
wire x_47148;
wire x_47149;
wire x_47150;
wire x_47151;
wire x_47152;
wire x_47153;
wire x_47154;
wire x_47155;
wire x_47156;
wire x_47157;
wire x_47158;
wire x_47159;
wire x_47160;
wire x_47161;
wire x_47162;
wire x_47163;
wire x_47164;
wire x_47165;
wire x_47166;
wire x_47167;
wire x_47168;
wire x_47169;
wire x_47170;
wire x_47171;
wire x_47172;
wire x_47173;
wire x_47174;
wire x_47175;
wire x_47176;
wire x_47177;
wire x_47178;
wire x_47179;
wire x_47180;
wire x_47181;
wire x_47182;
wire x_47183;
wire x_47184;
wire x_47185;
wire x_47186;
wire x_47187;
wire x_47188;
wire x_47189;
wire x_47190;
wire x_47191;
wire x_47192;
wire x_47193;
wire x_47194;
wire x_47195;
wire x_47196;
wire x_47197;
wire x_47198;
wire x_47199;
wire x_47200;
wire x_47201;
wire x_47202;
wire x_47203;
wire x_47204;
wire x_47205;
wire x_47206;
wire x_47207;
wire x_47208;
wire x_47209;
wire x_47210;
wire x_47211;
wire x_47212;
wire x_47213;
wire x_47214;
wire x_47215;
wire x_47216;
wire x_47217;
wire x_47218;
wire x_47219;
wire x_47220;
wire x_47221;
wire x_47222;
wire x_47223;
wire x_47224;
wire x_47225;
wire x_47226;
wire x_47227;
wire x_47228;
wire x_47229;
wire x_47230;
wire x_47231;
wire x_47232;
wire x_47233;
wire x_47234;
wire x_47235;
wire x_47236;
wire x_47237;
wire x_47238;
wire x_47239;
wire x_47240;
wire x_47241;
wire x_47242;
wire x_47243;
wire x_47244;
wire x_47245;
wire x_47246;
wire x_47247;
wire x_47248;
wire x_47249;
wire x_47250;
wire x_47251;
wire x_47252;
wire x_47253;
wire x_47254;
wire x_47255;
wire x_47256;
wire x_47257;
wire x_47258;
wire x_47259;
wire x_47260;
wire x_47261;
wire x_47262;
wire x_47263;
wire x_47264;
wire x_47265;
wire x_47266;
wire x_47267;
wire x_47268;
wire x_47269;
wire x_47270;
wire x_47271;
wire x_47272;
wire x_47273;
wire x_47274;
wire x_47275;
wire x_47276;
wire x_47277;
wire x_47278;
wire x_47279;
wire x_47280;
wire x_47281;
wire x_47282;
wire x_47283;
wire x_47284;
wire x_47285;
wire x_47286;
wire x_47287;
wire x_47288;
wire x_47289;
wire x_47290;
wire x_47291;
wire x_47292;
wire x_47293;
wire x_47294;
wire x_47295;
wire x_47296;
wire x_47297;
wire x_47298;
wire x_47299;
wire x_47300;
wire x_47301;
wire x_47302;
wire x_47303;
wire x_47304;
wire x_47305;
wire x_47306;
wire x_47307;
wire x_47308;
wire x_47309;
wire x_47310;
wire x_47311;
wire x_47312;
wire x_47313;
wire x_47314;
wire x_47315;
wire x_47316;
wire x_47317;
wire x_47318;
wire x_47319;
wire x_47320;
wire x_47321;
wire x_47322;
wire x_47323;
wire x_47324;
wire x_47325;
wire x_47326;
wire x_47327;
wire x_47328;
wire x_47329;
wire x_47330;
wire x_47331;
wire x_47332;
wire x_47333;
wire x_47334;
wire x_47335;
wire x_47336;
wire x_47337;
wire x_47338;
wire x_47339;
wire x_47340;
wire x_47341;
wire x_47342;
wire x_47343;
wire x_47344;
wire x_47345;
wire x_47346;
wire x_47347;
wire x_47348;
wire x_47349;
wire x_47350;
wire x_47351;
wire x_47352;
wire x_47353;
wire x_47354;
wire x_47355;
wire x_47356;
wire x_47357;
wire x_47358;
wire x_47359;
wire x_47360;
wire x_47361;
wire x_47362;
wire x_47363;
wire x_47364;
wire x_47365;
wire x_47366;
wire x_47367;
wire x_47368;
wire x_47369;
wire x_47370;
wire x_47371;
wire x_47372;
wire x_47373;
wire x_47374;
wire x_47375;
wire x_47376;
wire x_47377;
wire x_47378;
wire x_47379;
wire x_47380;
wire x_47381;
wire x_47382;
wire x_47383;
wire x_47384;
wire x_47385;
wire x_47386;
wire x_47387;
wire x_47388;
wire x_47389;
wire x_47390;
wire x_47391;
wire x_47392;
wire x_47393;
wire x_47394;
wire x_47395;
wire x_47396;
wire x_47397;
wire x_47398;
wire x_47399;
wire x_47400;
wire x_47401;
wire x_47402;
wire x_47403;
wire x_47404;
wire x_47405;
wire x_47406;
wire x_47407;
wire x_47408;
wire x_47409;
wire x_47410;
wire x_47411;
wire x_47412;
wire x_47413;
wire x_47414;
wire x_47415;
wire x_47416;
wire x_47417;
wire x_47418;
wire x_47419;
wire x_47420;
wire x_47421;
wire x_47422;
wire x_47423;
wire x_47424;
wire x_47425;
wire x_47426;
wire x_47427;
wire x_47428;
wire x_47429;
wire x_47430;
wire x_47431;
wire x_47432;
wire x_47433;
wire x_47434;
wire x_47435;
wire x_47436;
wire x_47437;
wire x_47438;
wire x_47439;
wire x_47440;
wire x_47441;
wire x_47442;
wire x_47443;
wire x_47444;
wire x_47445;
wire x_47446;
wire x_47447;
wire x_47448;
wire x_47449;
wire x_47450;
wire x_47451;
wire x_47452;
wire x_47453;
wire x_47454;
wire x_47455;
wire x_47456;
wire x_47457;
wire x_47458;
wire x_47459;
wire x_47460;
wire x_47461;
wire x_47462;
wire x_47463;
wire x_47464;
wire x_47465;
wire x_47466;
wire x_47467;
wire x_47468;
wire x_47469;
wire x_47470;
wire x_47471;
wire x_47472;
wire x_47473;
wire x_47474;
wire x_47475;
wire x_47476;
wire x_47477;
wire x_47478;
wire x_47479;
wire x_47480;
wire x_47481;
wire x_47482;
wire x_47483;
wire x_47484;
wire x_47485;
wire x_47486;
wire x_47487;
wire x_47488;
wire x_47489;
wire x_47490;
wire x_47491;
wire x_47492;
wire x_47493;
wire x_47494;
wire x_47495;
wire x_47496;
wire x_47497;
wire x_47498;
wire x_47499;
wire x_47500;
wire x_47501;
wire x_47502;
wire x_47503;
wire x_47504;
wire x_47505;
wire x_47506;
wire x_47507;
wire x_47508;
wire x_47509;
wire x_47510;
wire x_47511;
wire x_47512;
wire x_47513;
wire x_47514;
wire x_47515;
wire x_47516;
wire x_47517;
wire x_47518;
wire x_47519;
wire x_47520;
wire x_47521;
wire x_47522;
wire x_47523;
wire x_47524;
wire x_47525;
wire x_47526;
wire x_47527;
wire x_47528;
wire x_47529;
wire x_47530;
wire x_47531;
wire x_47532;
wire x_47533;
wire x_47534;
wire x_47535;
wire x_47536;
wire x_47537;
wire x_47538;
wire x_47539;
wire x_47540;
wire x_47541;
wire x_47542;
wire x_47543;
wire x_47544;
wire x_47545;
wire x_47546;
wire x_47547;
wire x_47548;
wire x_47549;
wire x_47550;
wire x_47551;
wire x_47552;
wire x_47553;
wire x_47554;
wire x_47555;
wire x_47556;
wire x_47557;
wire x_47558;
wire x_47559;
wire x_47560;
wire x_47561;
wire x_47562;
wire x_47563;
wire x_47564;
wire x_47565;
wire x_47566;
wire x_47567;
wire x_47568;
wire x_47569;
wire x_47570;
wire x_47571;
wire x_47572;
wire x_47573;
wire x_47574;
wire x_47575;
wire x_47576;
wire x_47577;
wire x_47578;
wire x_47579;
wire x_47580;
wire x_47581;
wire x_47582;
wire x_47583;
wire x_47584;
wire x_47585;
wire x_47586;
wire x_47587;
wire x_47588;
wire x_47589;
wire x_47590;
wire x_47591;
wire x_47592;
wire x_47593;
wire x_47594;
wire x_47595;
wire x_47596;
wire x_47597;
wire x_47598;
wire x_47599;
wire x_47600;
wire x_47601;
wire x_47602;
wire x_47603;
wire x_47604;
wire x_47605;
wire x_47606;
wire x_47607;
wire x_47608;
wire x_47609;
wire x_47610;
wire x_47611;
wire x_47612;
wire x_47613;
wire x_47614;
wire x_47615;
wire x_47616;
wire x_47617;
wire x_47618;
wire x_47619;
wire x_47620;
wire x_47621;
wire x_47622;
wire x_47623;
wire x_47624;
wire x_47625;
wire x_47626;
wire x_47627;
wire x_47628;
wire x_47629;
wire x_47630;
wire x_47631;
wire x_47632;
wire x_47633;
wire x_47634;
wire x_47635;
wire x_47636;
wire x_47637;
wire x_47638;
wire x_47639;
wire x_47640;
wire x_47641;
wire x_47642;
wire x_47643;
wire x_47644;
wire x_47645;
wire x_47646;
wire x_47647;
wire x_47648;
wire x_47649;
wire x_47650;
wire x_47651;
wire x_47652;
wire x_47653;
wire x_47654;
wire x_47655;
wire x_47656;
wire x_47657;
wire x_47658;
wire x_47659;
wire x_47660;
wire x_47661;
wire x_47662;
wire x_47663;
wire x_47664;
wire x_47665;
wire x_47666;
wire x_47667;
wire x_47668;
wire x_47669;
wire x_47670;
wire x_47671;
wire x_47672;
wire x_47673;
wire x_47674;
wire x_47675;
wire x_47676;
wire x_47677;
wire x_47678;
wire x_47679;
wire x_47680;
wire x_47681;
wire x_47682;
wire x_47683;
wire x_47684;
wire x_47685;
wire x_47686;
wire x_47687;
wire x_47688;
wire x_47689;
wire x_47690;
wire x_47691;
wire x_47692;
wire x_47693;
wire x_47694;
wire x_47695;
wire x_47696;
wire x_47697;
wire x_47698;
wire x_47699;
wire x_47700;
wire x_47701;
wire x_47702;
wire x_47703;
wire x_47704;
wire x_47705;
wire x_47706;
wire x_47707;
wire x_47708;
wire x_47709;
wire x_47710;
wire x_47711;
wire x_47712;
wire x_47713;
wire x_47714;
wire x_47715;
wire x_47716;
wire x_47717;
wire x_47718;
wire x_47719;
wire x_47720;
wire x_47721;
wire x_47722;
wire x_47723;
wire x_47724;
wire x_47725;
wire x_47726;
wire x_47727;
wire x_47728;
wire x_47729;
wire x_47730;
wire x_47731;
wire x_47732;
wire x_47733;
wire x_47734;
wire x_47735;
wire x_47736;
wire x_47737;
wire x_47738;
wire x_47739;
wire x_47740;
wire x_47741;
wire x_47742;
wire x_47743;
wire x_47744;
wire x_47745;
wire x_47746;
wire x_47747;
wire x_47748;
wire x_47749;
wire x_47750;
wire x_47751;
wire x_47752;
wire x_47753;
wire x_47754;
wire x_47755;
wire x_47756;
wire x_47757;
wire x_47758;
wire x_47759;
wire x_47760;
wire x_47761;
wire x_47762;
wire x_47763;
wire x_47764;
wire x_47765;
wire x_47766;
wire x_47767;
wire x_47768;
wire x_47769;
wire x_47770;
wire x_47771;
wire x_47772;
wire x_47773;
wire x_47774;
wire x_47775;
wire x_47776;
wire x_47777;
wire x_47778;
wire x_47779;
wire x_47780;
wire x_47781;
wire x_47782;
wire x_47783;
wire x_47784;
wire x_47785;
wire x_47786;
wire x_47787;
wire x_47788;
wire x_47789;
wire x_47790;
wire x_47791;
wire x_47792;
wire x_47793;
wire x_47794;
wire x_47795;
wire x_47796;
wire x_47797;
wire x_47798;
wire x_47799;
wire x_47800;
wire x_47801;
wire x_47802;
wire x_47803;
wire x_47804;
wire x_47805;
wire x_47806;
wire x_47807;
wire x_47808;
wire x_47809;
wire x_47810;
wire x_47811;
wire x_47812;
wire x_47813;
wire x_47814;
wire x_47815;
wire x_47816;
wire x_47817;
wire x_47818;
wire x_47819;
wire x_47820;
wire x_47821;
wire x_47822;
wire x_47823;
wire x_47824;
wire x_47825;
wire x_47826;
wire x_47827;
wire x_47828;
wire x_47829;
wire x_47830;
wire x_47831;
wire x_47832;
wire x_47833;
wire x_47834;
wire x_47835;
wire x_47836;
wire x_47837;
wire x_47838;
wire x_47839;
wire x_47840;
wire x_47841;
wire x_47842;
wire x_47843;
wire x_47844;
wire x_47845;
wire x_47846;
wire x_47847;
wire x_47848;
wire x_47849;
wire x_47850;
wire x_47851;
wire x_47852;
wire x_47853;
wire x_47854;
wire x_47855;
wire x_47856;
wire x_47857;
wire x_47858;
wire x_47859;
wire x_47860;
wire x_47861;
wire x_47862;
wire x_47863;
wire x_47864;
wire x_47865;
wire x_47866;
wire x_47867;
wire x_47868;
wire x_47869;
wire x_47870;
wire x_47871;
wire x_47872;
wire x_47873;
wire x_47874;
wire x_47875;
wire x_47876;
wire x_47877;
wire x_47878;
wire x_47879;
wire x_47880;
wire x_47881;
wire x_47882;
wire x_47883;
wire x_47884;
wire x_47885;
wire x_47886;
wire x_47887;
wire x_47888;
wire x_47889;
wire x_47890;
wire x_47891;
wire x_47892;
wire x_47893;
wire x_47894;
wire x_47895;
wire x_47896;
wire x_47897;
wire x_47898;
wire x_47899;
wire x_47900;
wire x_47901;
wire x_47902;
wire x_47903;
wire x_47904;
wire x_47905;
wire x_47906;
wire x_47907;
wire x_47908;
wire x_47909;
wire x_47910;
wire x_47911;
wire x_47912;
wire x_47913;
wire x_47914;
wire x_47915;
wire x_47916;
wire x_47917;
wire x_47918;
wire x_47919;
wire x_47920;
wire x_47921;
wire x_47922;
wire x_47923;
wire x_47924;
wire x_47925;
wire x_47926;
wire x_47927;
wire x_47928;
wire x_47929;
wire x_47930;
wire x_47931;
wire x_47932;
wire x_47933;
wire x_47934;
wire x_47935;
wire x_47936;
wire x_47937;
wire x_47938;
wire x_47939;
wire x_47940;
wire x_47941;
wire x_47942;
wire x_47943;
wire x_47944;
wire x_47945;
wire x_47946;
wire x_47947;
wire x_47948;
wire x_47949;
wire x_47950;
wire x_47951;
wire x_47952;
wire x_47953;
wire x_47954;
wire x_47955;
wire x_47956;
wire x_47957;
wire x_47958;
wire x_47959;
wire x_47960;
wire x_47961;
wire x_47962;
wire x_47963;
wire x_47964;
wire x_47965;
wire x_47966;
wire x_47967;
wire x_47968;
wire x_47969;
wire x_47970;
wire x_47971;
wire x_47972;
wire x_47973;
wire x_47974;
wire x_47975;
wire x_47976;
wire x_47977;
wire x_47978;
wire x_47979;
wire x_47980;
wire x_47981;
wire x_47982;
wire x_47983;
wire x_47984;
wire x_47985;
wire x_47986;
wire x_47987;
wire x_47988;
wire x_47989;
wire x_47990;
wire x_47991;
wire x_47992;
wire x_47993;
wire x_47994;
wire x_47995;
wire x_47996;
wire x_47997;
wire x_47998;
wire x_47999;
wire x_48000;
wire x_48001;
wire x_48002;
wire x_48003;
wire x_48004;
wire x_48005;
wire x_48006;
wire x_48007;
wire x_48008;
wire x_48009;
wire x_48010;
wire x_48011;
wire x_48012;
wire x_48013;
wire x_48014;
wire x_48015;
wire x_48016;
wire x_48017;
wire x_48018;
wire x_48019;
wire x_48020;
wire x_48021;
wire x_48022;
wire x_48023;
wire x_48024;
wire x_48025;
wire x_48026;
wire x_48027;
wire x_48028;
wire x_48029;
wire x_48030;
wire x_48031;
wire x_48032;
wire x_48033;
wire x_48034;
wire x_48035;
wire x_48036;
wire x_48037;
wire x_48038;
wire x_48039;
wire x_48040;
wire x_48041;
wire x_48042;
wire x_48043;
wire x_48044;
wire x_48045;
wire x_48046;
wire x_48047;
wire x_48048;
wire x_48049;
wire x_48050;
wire x_48051;
wire x_48052;
wire x_48053;
wire x_48054;
wire x_48055;
wire x_48056;
wire x_48057;
wire x_48058;
wire x_48059;
wire x_48060;
wire x_48061;
wire x_48062;
wire x_48063;
wire x_48064;
wire x_48065;
wire x_48066;
wire x_48067;
wire x_48068;
wire x_48069;
wire x_48070;
wire x_48071;
wire x_48072;
wire x_48073;
wire x_48074;
wire x_48075;
wire x_48076;
wire x_48077;
wire x_48078;
wire x_48079;
wire x_48080;
wire x_48081;
wire x_48082;
wire x_48083;
wire x_48084;
wire x_48085;
wire x_48086;
wire x_48087;
wire x_48088;
wire x_48089;
wire x_48090;
wire x_48091;
wire x_48092;
wire x_48093;
wire x_48094;
wire x_48095;
wire x_48096;
wire x_48097;
wire x_48098;
wire x_48099;
wire x_48100;
wire x_48101;
wire x_48102;
wire x_48103;
wire x_48104;
wire x_48105;
wire x_48106;
wire x_48107;
wire x_48108;
wire x_48109;
wire x_48110;
wire x_48111;
wire x_48112;
wire x_48113;
wire x_48114;
wire x_48115;
wire x_48116;
wire x_48117;
wire x_48118;
wire x_48119;
wire x_48120;
wire x_48121;
wire x_48122;
wire x_48123;
wire x_48124;
wire x_48125;
wire x_48126;
wire x_48127;
wire x_48128;
wire x_48129;
wire x_48130;
wire x_48131;
wire x_48132;
wire x_48133;
wire x_48134;
wire x_48135;
wire x_48136;
wire x_48137;
wire x_48138;
wire x_48139;
wire x_48140;
wire x_48141;
wire x_48142;
wire x_48143;
wire x_48144;
wire x_48145;
wire x_48146;
wire x_48147;
wire x_48148;
wire x_48149;
wire x_48150;
wire x_48151;
wire x_48152;
wire x_48153;
wire x_48154;
wire x_48155;
wire x_48156;
wire x_48157;
wire x_48158;
wire x_48159;
wire x_48160;
wire x_48161;
wire x_48162;
wire x_48163;
wire x_48164;
wire x_48165;
wire x_48166;
wire x_48167;
wire x_48168;
wire x_48169;
wire x_48170;
wire x_48171;
wire x_48172;
wire x_48173;
wire x_48174;
wire x_48175;
wire x_48176;
wire x_48177;
wire x_48178;
wire x_48179;
wire x_48180;
wire x_48181;
wire x_48182;
wire x_48183;
wire x_48184;
wire x_48185;
wire x_48186;
wire x_48187;
wire x_48188;
wire x_48189;
wire x_48190;
wire x_48191;
wire x_48192;
wire x_48193;
wire x_48194;
wire x_48195;
wire x_48196;
wire x_48197;
wire x_48198;
wire x_48199;
wire x_48200;
wire x_48201;
wire x_48202;
wire x_48203;
wire x_48204;
wire x_48205;
wire x_48206;
wire x_48207;
wire x_48208;
wire x_48209;
wire x_48210;
wire x_48211;
wire x_48212;
wire x_48213;
wire x_48214;
wire x_48215;
wire x_48216;
wire x_48217;
wire x_48218;
wire x_48219;
wire x_48220;
wire x_48221;
wire x_48222;
wire x_48223;
wire x_48224;
wire x_48225;
wire x_48226;
wire x_48227;
wire x_48228;
wire x_48229;
wire x_48230;
wire x_48231;
wire x_48232;
wire x_48233;
wire x_48234;
wire x_48235;
wire x_48236;
wire x_48237;
wire x_48238;
wire x_48239;
wire x_48240;
wire x_48241;
wire x_48242;
wire x_48243;
wire x_48244;
wire x_48245;
wire x_48246;
wire x_48247;
wire x_48248;
wire x_48249;
wire x_48250;
wire x_48251;
wire x_48252;
wire x_48253;
wire x_48254;
wire x_48255;
wire x_48256;
wire x_48257;
wire x_48258;
wire x_48259;
wire x_48260;
wire x_48261;
wire x_48262;
wire x_48263;
wire x_48264;
wire x_48265;
wire x_48266;
wire x_48267;
wire x_48268;
wire x_48269;
wire x_48270;
wire x_48271;
wire x_48272;
wire x_48273;
wire x_48274;
wire x_48275;
wire x_48276;
wire x_48277;
wire x_48278;
wire x_48279;
wire x_48280;
wire x_48281;
wire x_48282;
wire x_48283;
wire x_48284;
wire x_48285;
wire x_48286;
wire x_48287;
wire x_48288;
wire x_48289;
wire x_48290;
wire x_48291;
wire x_48292;
wire x_48293;
wire x_48294;
wire x_48295;
wire x_48296;
wire x_48297;
wire x_48298;
wire x_48299;
wire x_48300;
wire x_48301;
wire x_48302;
wire x_48303;
wire x_48304;
wire x_48305;
wire x_48306;
wire x_48307;
wire x_48308;
wire x_48309;
wire x_48310;
wire x_48311;
wire x_48312;
wire x_48313;
wire x_48314;
wire x_48315;
wire x_48316;
wire x_48317;
wire x_48318;
wire x_48319;
wire x_48320;
wire x_48321;
wire x_48322;
wire x_48323;
wire x_48324;
wire x_48325;
wire x_48326;
wire x_48327;
wire x_48328;
wire x_48329;
wire x_48330;
wire x_48331;
wire x_48332;
wire x_48333;
wire x_48334;
wire x_48335;
wire x_48336;
wire x_48337;
wire x_48338;
wire x_48339;
wire x_48340;
wire x_48341;
wire x_48342;
wire x_48343;
wire x_48344;
wire x_48345;
wire x_48346;
wire x_48347;
wire x_48348;
wire x_48349;
wire x_48350;
wire x_48351;
wire x_48352;
wire x_48353;
wire x_48354;
wire x_48355;
wire x_48356;
wire x_48357;
wire x_48358;
wire x_48359;
wire x_48360;
wire x_48361;
wire x_48362;
wire x_48363;
wire x_48364;
wire x_48365;
wire x_48366;
wire x_48367;
wire x_48368;
wire x_48369;
wire x_48370;
wire x_48371;
wire x_48372;
wire x_48373;
wire x_48374;
wire x_48375;
wire x_48376;
wire x_48377;
wire x_48378;
wire x_48379;
wire x_48380;
wire x_48381;
wire x_48382;
wire x_48383;
wire x_48384;
wire x_48385;
wire x_48386;
wire x_48387;
wire x_48388;
wire x_48389;
wire x_48390;
wire x_48391;
wire x_48392;
wire x_48393;
wire x_48394;
wire x_48395;
wire x_48396;
wire x_48397;
wire x_48398;
wire x_48399;
wire x_48400;
wire x_48401;
wire x_48402;
wire x_48403;
wire x_48404;
wire x_48405;
wire x_48406;
wire x_48407;
wire x_48408;
wire x_48409;
wire x_48410;
wire x_48411;
wire x_48412;
wire x_48413;
wire x_48414;
wire x_48415;
wire x_48416;
wire x_48417;
wire x_48418;
wire x_48419;
wire x_48420;
wire x_48421;
wire x_48422;
wire x_48423;
wire x_48424;
wire x_48425;
wire x_48426;
wire x_48427;
wire x_48428;
wire x_48429;
wire x_48430;
wire x_48431;
wire x_48432;
wire x_48433;
wire x_48434;
wire x_48435;
wire x_48436;
wire x_48437;
wire x_48438;
wire x_48439;
wire x_48440;
wire x_48441;
wire x_48442;
wire x_48443;
wire x_48444;
wire x_48445;
wire x_48446;
wire x_48447;
wire x_48448;
wire x_48449;
wire x_48450;
wire x_48451;
wire x_48452;
wire x_48453;
wire x_48454;
wire x_48455;
wire x_48456;
wire x_48457;
wire x_48458;
wire x_48459;
wire x_48460;
wire x_48461;
wire x_48462;
wire x_48463;
wire x_48464;
wire x_48465;
wire x_48466;
wire x_48467;
wire x_48468;
wire x_48469;
wire x_48470;
wire x_48471;
wire x_48472;
wire x_48473;
wire x_48474;
wire x_48475;
wire x_48476;
wire x_48477;
wire x_48478;
wire x_48479;
wire x_48480;
wire x_48481;
wire x_48482;
wire x_48483;
wire x_48484;
wire x_48485;
wire x_48486;
wire x_48487;
wire x_48488;
wire x_48489;
wire x_48490;
wire x_48491;
wire x_48492;
wire x_48493;
wire x_48494;
wire x_48495;
wire x_48496;
wire x_48497;
wire x_48498;
wire x_48499;
wire x_48500;
wire x_48501;
wire x_48502;
wire x_48503;
wire x_48504;
wire x_48505;
wire x_48506;
wire x_48507;
wire x_48508;
wire x_48509;
wire x_48510;
wire x_48511;
wire x_48512;
wire x_48513;
wire x_48514;
wire x_48515;
wire x_48516;
wire x_48517;
wire x_48518;
wire x_48519;
wire x_48520;
wire x_48521;
wire x_48522;
wire x_48523;
wire x_48524;
wire x_48525;
wire x_48526;
wire x_48527;
wire x_48528;
wire x_48529;
wire x_48530;
wire x_48531;
wire x_48532;
wire x_48533;
wire x_48534;
wire x_48535;
wire x_48536;
wire x_48537;
wire x_48538;
wire x_48539;
wire x_48540;
wire x_48541;
wire x_48542;
wire x_48543;
wire x_48544;
wire x_48545;
wire x_48546;
wire x_48547;
wire x_48548;
wire x_48549;
wire x_48550;
wire x_48551;
wire x_48552;
wire x_48553;
wire x_48554;
wire x_48555;
wire x_48556;
wire x_48557;
wire x_48558;
wire x_48559;
wire x_48560;
wire x_48561;
wire x_48562;
wire x_48563;
wire x_48564;
wire x_48565;
wire x_48566;
wire x_48567;
wire x_48568;
wire x_48569;
wire x_48570;
wire x_48571;
wire x_48572;
wire x_48573;
wire x_48574;
wire x_48575;
wire x_48576;
wire x_48577;
wire x_48578;
wire x_48579;
wire x_48580;
wire x_48581;
wire x_48582;
wire x_48583;
wire x_48584;
wire x_48585;
wire x_48586;
wire x_48587;
wire x_48588;
wire x_48589;
wire x_48590;
wire x_48591;
wire x_48592;
wire x_48593;
wire x_48594;
wire x_48595;
wire x_48596;
wire x_48597;
wire x_48598;
wire x_48599;
wire x_48600;
wire x_48601;
wire x_48602;
wire x_48603;
wire x_48604;
wire x_48605;
wire x_48606;
wire x_48607;
wire x_48608;
wire x_48609;
wire x_48610;
wire x_48611;
wire x_48612;
wire x_48613;
wire x_48614;
wire x_48615;
wire x_48616;
wire x_48617;
wire x_48618;
wire x_48619;
wire x_48620;
wire x_48621;
wire x_48622;
wire x_48623;
wire x_48624;
wire x_48625;
wire x_48626;
wire x_48627;
wire x_48628;
wire x_48629;
wire x_48630;
wire x_48631;
wire x_48632;
wire x_48633;
wire x_48634;
wire x_48635;
wire x_48636;
wire x_48637;
wire x_48638;
wire x_48639;
wire x_48640;
wire x_48641;
wire x_48642;
wire x_48643;
wire x_48644;
wire x_48645;
wire x_48646;
wire x_48647;
wire x_48648;
wire x_48649;
wire x_48650;
wire x_48651;
wire x_48652;
wire x_48653;
wire x_48654;
wire x_48655;
wire x_48656;
wire x_48657;
wire x_48658;
wire x_48659;
wire x_48660;
wire x_48661;
wire x_48662;
wire x_48663;
wire x_48664;
wire x_48665;
wire x_48666;
wire x_48667;
wire x_48668;
wire x_48669;
wire x_48670;
wire x_48671;
wire x_48672;
wire x_48673;
wire x_48674;
wire x_48675;
wire x_48676;
wire x_48677;
wire x_48678;
wire x_48679;
wire x_48680;
wire x_48681;
wire x_48682;
wire x_48683;
wire x_48684;
wire x_48685;
wire x_48686;
wire x_48687;
wire x_48688;
wire x_48689;
wire x_48690;
wire x_48691;
wire x_48692;
wire x_48693;
wire x_48694;
wire x_48695;
wire x_48696;
wire x_48697;
wire x_48698;
wire x_48699;
wire x_48700;
wire x_48701;
wire x_48702;
wire x_48703;
wire x_48704;
wire x_48705;
wire x_48706;
wire x_48707;
wire x_48708;
wire x_48709;
wire x_48710;
wire x_48711;
wire x_48712;
wire x_48713;
wire x_48714;
wire x_48715;
wire x_48716;
wire x_48717;
wire x_48718;
wire x_48719;
wire x_48720;
wire x_48721;
wire x_48722;
wire x_48723;
wire x_48724;
wire x_48725;
wire x_48726;
wire x_48727;
wire x_48728;
wire x_48729;
wire x_48730;
wire x_48731;
wire x_48732;
wire x_48733;
wire x_48734;
wire x_48735;
wire x_48736;
wire x_48737;
wire x_48738;
wire x_48739;
wire x_48740;
wire x_48741;
wire x_48742;
wire x_48743;
wire x_48744;
wire x_48745;
wire x_48746;
wire x_48747;
wire x_48748;
wire x_48749;
wire x_48750;
wire x_48751;
wire x_48752;
wire x_48753;
wire x_48754;
wire x_48755;
wire x_48756;
wire x_48757;
wire x_48758;
wire x_48759;
wire x_48760;
wire x_48761;
wire x_48762;
wire x_48763;
wire x_48764;
wire x_48765;
wire x_48766;
wire x_48767;
wire x_48768;
wire x_48769;
wire x_48770;
wire x_48771;
wire x_48772;
wire x_48773;
wire x_48774;
wire x_48775;
wire x_48776;
wire x_48777;
wire x_48778;
wire x_48779;
wire x_48780;
wire x_48781;
wire x_48782;
wire x_48783;
wire x_48784;
wire x_48785;
wire x_48786;
wire x_48787;
wire x_48788;
wire x_48789;
wire x_48790;
wire x_48791;
wire x_48792;
wire x_48793;
wire x_48794;
wire x_48795;
wire x_48796;
wire x_48797;
wire x_48798;
wire x_48799;
wire x_48800;
wire x_48801;
wire x_48802;
wire x_48803;
wire x_48804;
wire x_48805;
wire x_48806;
wire x_48807;
wire x_48808;
wire x_48809;
wire x_48810;
wire x_48811;
wire x_48812;
wire x_48813;
wire x_48814;
wire x_48815;
wire x_48816;
wire x_48817;
wire x_48818;
wire x_48819;
wire x_48820;
wire x_48821;
wire x_48822;
wire x_48823;
wire x_48824;
wire x_48825;
wire x_48826;
wire x_48827;
wire x_48828;
wire x_48829;
wire x_48830;
wire x_48831;
wire x_48832;
wire x_48833;
wire x_48834;
wire x_48835;
wire x_48836;
wire x_48837;
wire x_48838;
wire x_48839;
wire x_48840;
wire x_48841;
wire x_48842;
wire x_48843;
wire x_48844;
wire x_48845;
wire x_48846;
wire x_48847;
wire x_48848;
wire x_48849;
wire x_48850;
wire x_48851;
wire x_48852;
wire x_48853;
wire x_48854;
wire x_48855;
wire x_48856;
wire x_48857;
wire x_48858;
wire x_48859;
wire x_48860;
wire x_48861;
wire x_48862;
wire x_48863;
wire x_48864;
wire x_48865;
wire x_48866;
wire x_48867;
wire x_48868;
wire x_48869;
wire x_48870;
wire x_48871;
wire x_48872;
wire x_48873;
wire x_48874;
wire x_48875;
wire x_48876;
wire x_48877;
wire x_48878;
wire x_48879;
wire x_48880;
wire x_48881;
wire x_48882;
wire x_48883;
wire x_48884;
wire x_48885;
wire x_48886;
wire x_48887;
wire x_48888;
wire x_48889;
wire x_48890;
wire x_48891;
wire x_48892;
wire x_48893;
wire x_48894;
wire x_48895;
wire x_48896;
wire x_48897;
wire x_48898;
wire x_48899;
wire x_48900;
wire x_48901;
wire x_48902;
wire x_48903;
wire x_48904;
wire x_48905;
wire x_48906;
wire x_48907;
wire x_48908;
wire x_48909;
wire x_48910;
wire x_48911;
wire x_48912;
wire x_48913;
wire x_48914;
wire x_48915;
wire x_48916;
wire x_48917;
wire x_48918;
wire x_48919;
wire x_48920;
wire x_48921;
wire x_48922;
wire x_48923;
wire x_48924;
wire x_48925;
wire x_48926;
wire x_48927;
wire x_48928;
wire x_48929;
wire x_48930;
wire x_48931;
wire x_48932;
wire x_48933;
wire x_48934;
wire x_48935;
wire x_48936;
wire x_48937;
wire x_48938;
wire x_48939;
wire x_48940;
wire x_48941;
wire x_48942;
wire x_48943;
wire x_48944;
wire x_48945;
wire x_48946;
wire x_48947;
wire x_48948;
wire x_48949;
wire x_48950;
wire x_48951;
wire x_48952;
wire x_48953;
wire x_48954;
wire x_48955;
wire x_48956;
wire x_48957;
wire x_48958;
wire x_48959;
wire x_48960;
wire x_48961;
wire x_48962;
wire x_48963;
wire x_48964;
wire x_48965;
wire x_48966;
wire x_48967;
wire x_48968;
wire x_48969;
wire x_48970;
wire x_48971;
wire x_48972;
wire x_48973;
wire x_48974;
wire x_48975;
wire x_48976;
wire x_48977;
wire x_48978;
wire x_48979;
wire x_48980;
wire x_48981;
wire x_48982;
wire x_48983;
wire x_48984;
wire x_48985;
wire x_48986;
wire x_48987;
wire x_48988;
wire x_48989;
wire x_48990;
wire x_48991;
wire x_48992;
wire x_48993;
wire x_48994;
wire x_48995;
wire x_48996;
wire x_48997;
wire x_48998;
wire x_48999;
wire x_49000;
wire x_49001;
wire x_49002;
wire x_49003;
wire x_49004;
wire x_49005;
wire x_49006;
wire x_49007;
wire x_49008;
wire x_49009;
wire x_49010;
wire x_49011;
wire x_49012;
wire x_49013;
wire x_49014;
wire x_49015;
wire x_49016;
wire x_49017;
wire x_49018;
wire x_49019;
wire x_49020;
wire x_49021;
wire x_49022;
wire x_49023;
wire x_49024;
wire x_49025;
wire x_49026;
wire x_49027;
wire x_49028;
wire x_49029;
wire x_49030;
wire x_49031;
wire x_49032;
wire x_49033;
wire x_49034;
wire x_49035;
wire x_49036;
wire x_49037;
wire x_49038;
wire x_49039;
wire x_49040;
wire x_49041;
wire x_49042;
wire x_49043;
wire x_49044;
wire x_49045;
wire x_49046;
wire x_49047;
wire x_49048;
wire x_49049;
wire x_49050;
wire x_49051;
wire x_49052;
wire x_49053;
wire x_49054;
wire x_49055;
wire x_49056;
wire x_49057;
wire x_49058;
wire x_49059;
wire x_49060;
wire x_49061;
wire x_49062;
wire x_49063;
wire x_49064;
wire x_49065;
wire x_49066;
wire x_49067;
wire x_49068;
wire x_49069;
wire x_49070;
wire x_49071;
wire x_49072;
wire x_49073;
wire x_49074;
wire x_49075;
wire x_49076;
wire x_49077;
wire x_49078;
wire x_49079;
wire x_49080;
wire x_49081;
wire x_49082;
wire x_49083;
wire x_49084;
wire x_49085;
wire x_49086;
wire x_49087;
wire x_49088;
wire x_49089;
wire x_49090;
wire x_49091;
wire x_49092;
wire x_49093;
wire x_49094;
wire x_49095;
wire x_49096;
wire x_49097;
wire x_49098;
wire x_49099;
wire x_49100;
wire x_49101;
wire x_49102;
wire x_49103;
wire x_49104;
wire x_49105;
wire x_49106;
wire x_49107;
wire x_49108;
wire x_49109;
wire x_49110;
wire x_49111;
wire x_49112;
wire x_49113;
wire x_49114;
wire x_49115;
wire x_49116;
wire x_49117;
wire x_49118;
wire x_49119;
wire x_49120;
wire x_49121;
wire x_49122;
wire x_49123;
wire x_49124;
wire x_49125;
wire x_49126;
wire x_49127;
wire x_49128;
wire x_49129;
wire x_49130;
wire x_49131;
wire x_49132;
wire x_49133;
wire x_49134;
wire x_49135;
wire x_49136;
wire x_49137;
wire x_49138;
wire x_49139;
wire x_49140;
wire x_49141;
wire x_49142;
wire x_49143;
wire x_49144;
wire x_49145;
wire x_49146;
wire x_49147;
wire x_49148;
wire x_49149;
wire x_49150;
wire x_49151;
wire x_49152;
wire x_49153;
wire x_49154;
wire x_49155;
wire x_49156;
wire x_49157;
wire x_49158;
wire x_49159;
wire x_49160;
wire x_49161;
wire x_49162;
wire x_49163;
wire x_49164;
wire x_49165;
wire x_49166;
wire x_49167;
wire x_49168;
wire x_49169;
wire x_49170;
wire x_49171;
wire x_49172;
wire x_49173;
wire x_49174;
wire x_49175;
wire x_49176;
wire x_49177;
wire x_49178;
wire x_49179;
wire x_49180;
wire x_49181;
wire x_49182;
wire x_49183;
wire x_49184;
wire x_49185;
wire x_49186;
wire x_49187;
wire x_49188;
wire x_49189;
wire x_49190;
wire x_49191;
wire x_49192;
wire x_49193;
wire x_49194;
wire x_49195;
wire x_49196;
wire x_49197;
wire x_49198;
wire x_49199;
wire x_49200;
wire x_49201;
wire x_49202;
wire x_49203;
wire x_49204;
wire x_49205;
wire x_49206;
wire x_49207;
wire x_49208;
wire x_49209;
wire x_49210;
wire x_49211;
wire x_49212;
wire x_49213;
wire x_49214;
wire x_49215;
wire x_49216;
wire x_49217;
wire x_49218;
wire x_49219;
wire x_49220;
wire x_49221;
wire x_49222;
wire x_49223;
wire x_49224;
wire x_49225;
wire x_49226;
wire x_49227;
wire x_49228;
wire x_49229;
wire x_49230;
wire x_49231;
wire x_49232;
wire x_49233;
wire x_49234;
wire x_49235;
wire x_49236;
wire x_49237;
wire x_49238;
wire x_49239;
wire x_49240;
wire x_49241;
wire x_49242;
wire x_49243;
wire x_49244;
wire x_49245;
wire x_49246;
wire x_49247;
wire x_49248;
wire x_49249;
wire x_49250;
wire x_49251;
wire x_49252;
wire x_49253;
wire x_49254;
wire x_49255;
wire x_49256;
wire x_49257;
wire x_49258;
wire x_49259;
wire x_49260;
wire x_49261;
wire x_49262;
wire x_49263;
wire x_49264;
wire x_49265;
wire x_49266;
wire x_49267;
wire x_49268;
wire x_49269;
wire x_49270;
wire x_49271;
wire x_49272;
wire x_49273;
wire x_49274;
wire x_49275;
wire x_49276;
wire x_49277;
wire x_49278;
wire x_49279;
wire x_49280;
wire x_49281;
wire x_49282;
wire x_49283;
wire x_49284;
wire x_49285;
wire x_49286;
wire x_49287;
wire x_49288;
wire x_49289;
wire x_49290;
wire x_49291;
wire x_49292;
wire x_49293;
wire x_49294;
wire x_49295;
wire x_49296;
wire x_49297;
wire x_49298;
wire x_49299;
wire x_49300;
wire x_49301;
wire x_49302;
wire x_49303;
wire x_49304;
wire x_49305;
wire x_49306;
wire x_49307;
wire x_49308;
wire x_49309;
wire x_49310;
wire x_49311;
wire x_49312;
wire x_49313;
wire x_49314;
wire x_49315;
wire x_49316;
wire x_49317;
wire x_49318;
wire x_49319;
wire x_49320;
wire x_49321;
wire x_49322;
wire x_49323;
wire x_49324;
wire x_49325;
wire x_49326;
wire x_49327;
wire x_49328;
wire x_49329;
wire x_49330;
wire x_49331;
wire x_49332;
wire x_49333;
wire x_49334;
wire x_49335;
wire x_49336;
wire x_49337;
wire x_49338;
wire x_49339;
wire x_49340;
wire x_49341;
wire x_49342;
wire x_49343;
wire x_49344;
wire x_49345;
wire x_49346;
wire x_49347;
wire x_49348;
wire x_49349;
wire x_49350;
wire x_49351;
wire x_49352;
wire x_49353;
wire x_49354;
wire x_49355;
wire x_49356;
wire x_49357;
wire x_49358;
wire x_49359;
wire x_49360;
wire x_49361;
wire x_49362;
wire x_49363;
wire x_49364;
wire x_49365;
wire x_49366;
wire x_49367;
wire x_49368;
wire x_49369;
wire x_49370;
wire x_49371;
wire x_49372;
wire x_49373;
wire x_49374;
wire x_49375;
wire x_49376;
wire x_49377;
wire x_49378;
wire x_49379;
wire x_49380;
wire x_49381;
wire x_49382;
wire x_49383;
wire x_49384;
wire x_49385;
wire x_49386;
wire x_49387;
wire x_49388;
wire x_49389;
wire x_49390;
wire x_49391;
wire x_49392;
wire x_49393;
wire x_49394;
wire x_49395;
wire x_49396;
wire x_49397;
wire x_49398;
wire x_49399;
wire x_49400;
wire x_49401;
wire x_49402;
wire x_49403;
wire x_49404;
wire x_49405;
wire x_49406;
wire x_49407;
wire x_49408;
wire x_49409;
wire x_49410;
wire x_49411;
wire x_49412;
wire x_49413;
wire x_49414;
wire x_49415;
wire x_49416;
wire x_49417;
wire x_49418;
wire x_49419;
wire x_49420;
wire x_49421;
wire x_49422;
wire x_49423;
wire x_49424;
wire x_49425;
wire x_49426;
wire x_49427;
wire x_49428;
wire x_49429;
wire x_49430;
wire x_49431;
wire x_49432;
wire x_49433;
wire x_49434;
wire x_49435;
wire x_49436;
wire x_49437;
wire x_49438;
wire x_49439;
wire x_49440;
wire x_49441;
wire x_49442;
wire x_49443;
wire x_49444;
wire x_49445;
wire x_49446;
wire x_49447;
wire x_49448;
wire x_49449;
wire x_49450;
wire x_49451;
wire x_49452;
wire x_49453;
wire x_49454;
wire x_49455;
wire x_49456;
wire x_49457;
wire x_49458;
wire x_49459;
wire x_49460;
wire x_49461;
wire x_49462;
wire x_49463;
wire x_49464;
wire x_49465;
wire x_49466;
wire x_49467;
wire x_49468;
wire x_49469;
wire x_49470;
wire x_49471;
wire x_49472;
wire x_49473;
wire x_49474;
wire x_49475;
wire x_49476;
wire x_49477;
wire x_49478;
wire x_49479;
wire x_49480;
wire x_49481;
wire x_49482;
wire x_49483;
wire x_49484;
wire x_49485;
wire x_49486;
wire x_49487;
wire x_49488;
wire x_49489;
wire x_49490;
wire x_49491;
wire x_49492;
wire x_49493;
wire x_49494;
wire x_49495;
wire x_49496;
wire x_49497;
wire x_49498;
wire x_49499;
wire x_49500;
wire x_49501;
wire x_49502;
wire x_49503;
wire x_49504;
wire x_49505;
wire x_49506;
wire x_49507;
wire x_49508;
wire x_49509;
wire x_49510;
wire x_49511;
wire x_49512;
wire x_49513;
wire x_49514;
wire x_49515;
wire x_49516;
wire x_49517;
wire x_49518;
wire x_49519;
wire x_49520;
wire x_49521;
wire x_49522;
wire x_49523;
wire x_49524;
wire x_49525;
wire x_49526;
wire x_49527;
wire x_49528;
wire x_49529;
wire x_49530;
wire x_49531;
wire x_49532;
wire x_49533;
wire x_49534;
wire x_49535;
wire x_49536;
wire x_49537;
wire x_49538;
wire x_49539;
wire x_49540;
wire x_49541;
wire x_49542;
wire x_49543;
wire x_49544;
wire x_49545;
wire x_49546;
wire x_49547;
wire x_49548;
wire x_49549;
wire x_49550;
wire x_49551;
wire x_49552;
wire x_49553;
wire x_49554;
wire x_49555;
wire x_49556;
wire x_49557;
wire x_49558;
wire x_49559;
wire x_49560;
wire x_49561;
wire x_49562;
wire x_49563;
wire x_49564;
wire x_49565;
wire x_49566;
wire x_49567;
wire x_49568;
wire x_49569;
wire x_49570;
wire x_49571;
wire x_49572;
wire x_49573;
wire x_49574;
wire x_49575;
wire x_49576;
wire x_49577;
wire x_49578;
wire x_49579;
wire x_49580;
wire x_49581;
wire x_49582;
wire x_49583;
wire x_49584;
wire x_49585;
wire x_49586;
wire x_49587;
wire x_49588;
wire x_49589;
wire x_49590;
wire x_49591;
wire x_49592;
wire x_49593;
wire x_49594;
wire x_49595;
wire x_49596;
wire x_49597;
wire x_49598;
wire x_49599;
wire x_49600;
wire x_49601;
wire x_49602;
wire x_49603;
wire x_49604;
wire x_49605;
wire x_49606;
wire x_49607;
wire x_49608;
wire x_49609;
wire x_49610;
wire x_49611;
wire x_49612;
wire x_49613;
wire x_49614;
wire x_49615;
wire x_49616;
wire x_49617;
wire x_49618;
wire x_49619;
wire x_49620;
wire x_49621;
wire x_49622;
wire x_49623;
wire x_49624;
wire x_49625;
wire x_49626;
wire x_49627;
wire x_49628;
wire x_49629;
wire x_49630;
wire x_49631;
wire x_49632;
wire x_49633;
wire x_49634;
wire x_49635;
wire x_49636;
wire x_49637;
wire x_49638;
wire x_49639;
wire x_49640;
wire x_49641;
wire x_49642;
wire x_49643;
wire x_49644;
wire x_49645;
wire x_49646;
wire x_49647;
wire x_49648;
wire x_49649;
wire x_49650;
wire x_49651;
wire x_49652;
wire x_49653;
wire x_49654;
wire x_49655;
wire x_49656;
wire x_49657;
wire x_49658;
wire x_49659;
wire x_49660;
wire x_49661;
wire x_49662;
wire x_49663;
wire x_49664;
wire x_49665;
wire x_49666;
wire x_49667;
wire x_49668;
wire x_49669;
wire x_49670;
wire x_49671;
wire x_49672;
wire x_49673;
wire x_49674;
wire x_49675;
wire x_49676;
wire x_49677;
wire x_49678;
wire x_49679;
wire x_49680;
wire x_49681;
wire x_49682;
wire x_49683;
wire x_49684;
wire x_49685;
wire x_49686;
wire x_49687;
wire x_49688;
wire x_49689;
wire x_49690;
wire x_49691;
wire x_49692;
wire x_49693;
wire x_49694;
wire x_49695;
wire x_49696;
wire x_49697;
wire x_49698;
wire x_49699;
wire x_49700;
wire x_49701;
wire x_49702;
wire x_49703;
wire x_49704;
wire x_49705;
wire x_49706;
wire x_49707;
wire x_49708;
wire x_49709;
wire x_49710;
wire x_49711;
wire x_49712;
wire x_49713;
wire x_49714;
wire x_49715;
wire x_49716;
wire x_49717;
wire x_49718;
wire x_49719;
wire x_49720;
wire x_49721;
wire x_49722;
wire x_49723;
wire x_49724;
wire x_49725;
wire x_49726;
wire x_49727;
wire x_49728;
wire x_49729;
wire x_49730;
wire x_49731;
wire x_49732;
wire x_49733;
wire x_49734;
wire x_49735;
wire x_49736;
wire x_49737;
wire x_49738;
wire x_49739;
wire x_49740;
wire x_49741;
wire x_49742;
wire x_49743;
wire x_49744;
wire x_49745;
wire x_49746;
wire x_49747;
wire x_49748;
wire x_49749;
wire x_49750;
wire x_49751;
wire x_49752;
wire x_49753;
wire x_49754;
wire x_49755;
wire x_49756;
wire x_49757;
wire x_49758;
wire x_49759;
wire x_49760;
wire x_49761;
wire x_49762;
wire x_49763;
wire x_49764;
wire x_49765;
wire x_49766;
wire x_49767;
wire x_49768;
wire x_49769;
wire x_49770;
wire x_49771;
wire x_49772;
wire x_49773;
wire x_49774;
wire x_49775;
wire x_49776;
wire x_49777;
wire x_49778;
wire x_49779;
wire x_49780;
wire x_49781;
wire x_49782;
wire x_49783;
wire x_49784;
wire x_49785;
wire x_49786;
wire x_49787;
wire x_49788;
wire x_49789;
wire x_49790;
wire x_49791;
wire x_49792;
wire x_49793;
wire x_49794;
wire x_49795;
wire x_49796;
wire x_49797;
wire x_49798;
wire x_49799;
wire x_49800;
wire x_49801;
wire x_49802;
wire x_49803;
wire x_49804;
wire x_49805;
wire x_49806;
wire x_49807;
wire x_49808;
wire x_49809;
wire x_49810;
wire x_49811;
wire x_49812;
wire x_49813;
wire x_49814;
wire x_49815;
wire x_49816;
wire x_49817;
wire x_49818;
wire x_49819;
wire x_49820;
wire x_49821;
wire x_49822;
wire x_49823;
wire x_49824;
wire x_49825;
wire x_49826;
wire x_49827;
wire x_49828;
wire x_49829;
wire x_49830;
wire x_49831;
wire x_49832;
wire x_49833;
wire x_49834;
wire x_49835;
wire x_49836;
wire x_49837;
wire x_49838;
wire x_49839;
wire x_49840;
wire x_49841;
wire x_49842;
wire x_49843;
wire x_49844;
wire x_49845;
wire x_49846;
wire x_49847;
wire x_49848;
wire x_49849;
wire x_49850;
wire x_49851;
wire x_49852;
wire x_49853;
wire x_49854;
wire x_49855;
wire x_49856;
wire x_49857;
wire x_49858;
wire x_49859;
wire x_49860;
wire x_49861;
wire x_49862;
wire x_49863;
wire x_49864;
wire x_49865;
wire x_49866;
wire x_49867;
wire x_49868;
wire x_49869;
wire x_49870;
wire x_49871;
wire x_49872;
wire x_49873;
wire x_49874;
wire x_49875;
wire x_49876;
wire x_49877;
wire x_49878;
wire x_49879;
wire x_49880;
wire x_49881;
wire x_49882;
wire x_49883;
wire x_49884;
wire x_49885;
wire x_49886;
wire x_49887;
wire x_49888;
wire x_49889;
wire x_49890;
wire x_49891;
wire x_49892;
wire x_49893;
wire x_49894;
wire x_49895;
wire x_49896;
wire x_49897;
wire x_49898;
wire x_49899;
wire x_49900;
wire x_49901;
wire x_49902;
wire x_49903;
wire x_49904;
wire x_49905;
wire x_49906;
wire x_49907;
wire x_49908;
wire x_49909;
wire x_49910;
wire x_49911;
wire x_49912;
wire x_49913;
wire x_49914;
wire x_49915;
wire x_49916;
wire x_49917;
wire x_49918;
wire x_49919;
wire x_49920;
wire x_49921;
wire x_49922;
wire x_49923;
wire x_49924;
wire x_49925;
wire x_49926;
wire x_49927;
wire x_49928;
wire x_49929;
wire x_49930;
wire x_49931;
wire x_49932;
wire x_49933;
wire x_49934;
wire x_49935;
wire x_49936;
wire x_49937;
wire x_49938;
wire x_49939;
wire x_49940;
wire x_49941;
wire x_49942;
wire x_49943;
wire x_49944;
wire x_49945;
wire x_49946;
wire x_49947;
wire x_49948;
wire x_49949;
wire x_49950;
wire x_49951;
wire x_49952;
wire x_49953;
wire x_49954;
wire x_49955;
wire x_49956;
wire x_49957;
wire x_49958;
wire x_49959;
wire x_49960;
wire x_49961;
wire x_49962;
wire x_49963;
wire x_49964;
wire x_49965;
wire x_49966;
wire x_49967;
wire x_49968;
wire x_49969;
wire x_49970;
wire x_49971;
wire x_49972;
wire x_49973;
wire x_49974;
wire x_49975;
wire x_49976;
wire x_49977;
wire x_49978;
wire x_49979;
wire x_49980;
wire x_49981;
wire x_49982;
wire x_49983;
wire x_49984;
wire x_49985;
wire x_49986;
wire x_49987;
wire x_49988;
wire x_49989;
wire x_49990;
wire x_49991;
wire x_49992;
wire x_49993;
wire x_49994;
wire x_49995;
wire x_49996;
wire x_49997;
wire x_49998;
wire x_49999;
wire x_50000;
wire x_50001;
wire x_50002;
wire x_50003;
wire x_50004;
wire x_50005;
wire x_50006;
wire x_50007;
wire x_50008;
wire x_50009;
wire x_50010;
wire x_50011;
wire x_50012;
wire x_50013;
wire x_50014;
wire x_50015;
wire x_50016;
wire x_50017;
wire x_50018;
wire x_50019;
wire x_50020;
wire x_50021;
wire x_50022;
wire x_50023;
wire x_50024;
wire x_50025;
wire x_50026;
wire x_50027;
wire x_50028;
wire x_50029;
wire x_50030;
wire x_50031;
wire x_50032;
wire x_50033;
wire x_50034;
wire x_50035;
wire x_50036;
wire x_50037;
wire x_50038;
wire x_50039;
wire x_50040;
wire x_50041;
wire x_50042;
wire x_50043;
wire x_50044;
wire x_50045;
wire x_50046;
wire x_50047;
wire x_50048;
wire x_50049;
wire x_50050;
wire x_50051;
wire x_50052;
wire x_50053;
wire x_50054;
wire x_50055;
wire x_50056;
wire x_50057;
wire x_50058;
wire x_50059;
wire x_50060;
wire x_50061;
wire x_50062;
wire x_50063;
wire x_50064;
wire x_50065;
wire x_50066;
wire x_50067;
wire x_50068;
wire x_50069;
wire x_50070;
wire x_50071;
wire x_50072;
wire x_50073;
wire x_50074;
wire x_50075;
wire x_50076;
wire x_50077;
wire x_50078;
wire x_50079;
wire x_50080;
wire x_50081;
wire x_50082;
wire x_50083;
wire x_50084;
wire x_50085;
wire x_50086;
wire x_50087;
wire x_50088;
wire x_50089;
wire x_50090;
wire x_50091;
wire x_50092;
wire x_50093;
wire x_50094;
wire x_50095;
wire x_50096;
wire x_50097;
wire x_50098;
wire x_50099;
wire x_50100;
wire x_50101;
wire x_50102;
wire x_50103;
wire x_50104;
wire x_50105;
wire x_50106;
wire x_50107;
wire x_50108;
wire x_50109;
wire x_50110;
wire x_50111;
wire x_50112;
wire x_50113;
wire x_50114;
wire x_50115;
wire x_50116;
wire x_50117;
wire x_50118;
wire x_50119;
wire x_50120;
wire x_50121;
wire x_50122;
wire x_50123;
wire x_50124;
wire x_50125;
wire x_50126;
wire x_50127;
wire x_50128;
wire x_50129;
wire x_50130;
wire x_50131;
wire x_50132;
wire x_50133;
wire x_50134;
wire x_50135;
wire x_50136;
wire x_50137;
wire x_50138;
wire x_50139;
wire x_50140;
wire x_50141;
wire x_50142;
wire x_50143;
wire x_50144;
wire x_50145;
wire x_50146;
wire x_50147;
wire x_50148;
wire x_50149;
wire x_50150;
wire x_50151;
wire x_50152;
wire x_50153;
wire x_50154;
wire x_50155;
wire x_50156;
wire x_50157;
wire x_50158;
wire x_50159;
wire x_50160;
wire x_50161;
wire x_50162;
wire x_50163;
wire x_50164;
wire x_50165;
wire x_50166;
wire x_50167;
wire x_50168;
wire x_50169;
wire x_50170;
wire x_50171;
wire x_50172;
wire x_50173;
wire x_50174;
wire x_50175;
wire x_50176;
wire x_50177;
wire x_50178;
wire x_50179;
wire x_50180;
wire x_50181;
wire x_50182;
wire x_50183;
wire x_50184;
wire x_50185;
wire x_50186;
wire x_50187;
wire x_50188;
wire x_50189;
wire x_50190;
wire x_50191;
wire x_50192;
wire x_50193;
wire x_50194;
wire x_50195;
wire x_50196;
wire x_50197;
wire x_50198;
wire x_50199;
wire x_50200;
wire x_50201;
wire x_50202;
wire x_50203;
wire x_50204;
wire x_50205;
wire x_50206;
wire x_50207;
wire x_50208;
wire x_50209;
wire x_50210;
wire x_50211;
wire x_50212;
wire x_50213;
wire x_50214;
wire x_50215;
wire x_50216;
wire x_50217;
wire x_50218;
wire x_50219;
wire x_50220;
wire x_50221;
wire x_50222;
wire x_50223;
wire x_50224;
wire x_50225;
wire x_50226;
wire x_50227;
wire x_50228;
wire x_50229;
wire x_50230;
wire x_50231;
wire x_50232;
wire x_50233;
wire x_50234;
wire x_50235;
wire x_50236;
wire x_50237;
wire x_50238;
wire x_50239;
wire x_50240;
wire x_50241;
wire x_50242;
wire x_50243;
wire x_50244;
wire x_50245;
wire x_50246;
wire x_50247;
wire x_50248;
wire x_50249;
wire x_50250;
wire x_50251;
wire x_50252;
wire x_50253;
wire x_50254;
wire x_50255;
wire x_50256;
wire x_50257;
wire x_50258;
wire x_50259;
wire x_50260;
wire x_50261;
wire x_50262;
wire x_50263;
wire x_50264;
wire x_50265;
wire x_50266;
wire x_50267;
wire x_50268;
wire x_50269;
wire x_50270;
wire x_50271;
wire x_50272;
wire x_50273;
wire x_50274;
wire x_50275;
wire x_50276;
wire x_50277;
wire x_50278;
wire x_50279;
wire x_50280;
wire x_50281;
wire x_50282;
wire x_50283;
wire x_50284;
wire x_50285;
wire x_50286;
wire x_50287;
wire x_50288;
wire x_50289;
wire x_50290;
wire x_50291;
wire x_50292;
wire x_50293;
wire x_50294;
wire x_50295;
wire x_50296;
wire x_50297;
wire x_50298;
wire x_50299;
wire x_50300;
wire x_50301;
wire x_50302;
wire x_50303;
wire x_50304;
wire x_50305;
wire x_50306;
wire x_50307;
wire x_50308;
wire x_50309;
wire x_50310;
wire x_50311;
wire x_50312;
wire x_50313;
wire x_50314;
wire x_50315;
wire x_50316;
wire x_50317;
wire x_50318;
wire x_50319;
wire x_50320;
wire x_50321;
wire x_50322;
wire x_50323;
wire x_50324;
wire x_50325;
wire x_50326;
wire x_50327;
wire x_50328;
wire x_50329;
wire x_50330;
wire x_50331;
wire x_50332;
wire x_50333;
wire x_50334;
wire x_50335;
wire x_50336;
wire x_50337;
wire x_50338;
wire x_50339;
wire x_50340;
wire x_50341;
wire x_50342;
wire x_50343;
wire x_50344;
wire x_50345;
wire x_50346;
wire x_50347;
wire x_50348;
wire x_50349;
wire x_50350;
wire x_50351;
wire x_50352;
wire x_50353;
wire x_50354;
wire x_50355;
wire x_50356;
wire x_50357;
wire x_50358;
wire x_50359;
wire x_50360;
wire x_50361;
wire x_50362;
wire x_50363;
wire x_50364;
wire x_50365;
wire x_50366;
wire x_50367;
wire x_50368;
wire x_50369;
wire x_50370;
wire x_50371;
wire x_50372;
wire x_50373;
wire x_50374;
wire x_50375;
wire x_50376;
wire x_50377;
wire x_50378;
wire x_50379;
wire x_50380;
wire x_50381;
wire x_50382;
wire x_50383;
wire x_50384;
wire x_50385;
wire x_50386;
wire x_50387;
wire x_50388;
wire x_50389;
wire x_50390;
wire x_50391;
wire x_50392;
wire x_50393;
wire x_50394;
wire x_50395;
wire x_50396;
wire x_50397;
wire x_50398;
wire x_50399;
wire x_50400;
wire x_50401;
wire x_50402;
wire x_50403;
wire x_50404;
wire x_50405;
wire x_50406;
wire x_50407;
wire x_50408;
wire x_50409;
wire x_50410;
wire x_50411;
wire x_50412;
wire x_50413;
wire x_50414;
wire x_50415;
wire x_50416;
wire x_50417;
wire x_50418;
wire x_50419;
wire x_50420;
wire x_50421;
wire x_50422;
wire x_50423;
wire x_50424;
wire x_50425;
wire x_50426;
wire x_50427;
wire x_50428;
wire x_50429;
wire x_50430;
wire x_50431;
wire x_50432;
wire x_50433;
wire x_50434;
wire x_50435;
wire x_50436;
wire x_50437;
wire x_50438;
wire x_50439;
wire x_50440;
wire x_50441;
wire x_50442;
wire x_50443;
wire x_50444;
wire x_50445;
wire x_50446;
wire x_50447;
wire x_50448;
wire x_50449;
wire x_50450;
wire x_50451;
wire x_50452;
wire x_50453;
wire x_50454;
wire x_50455;
wire x_50456;
wire x_50457;
wire x_50458;
wire x_50459;
wire x_50460;
wire x_50461;
wire x_50462;
wire x_50463;
wire x_50464;
wire x_50465;
wire x_50466;
wire x_50467;
wire x_50468;
wire x_50469;
wire x_50470;
wire x_50471;
wire x_50472;
wire x_50473;
wire x_50474;
wire x_50475;
wire x_50476;
wire x_50477;
wire x_50478;
wire x_50479;
wire x_50480;
wire x_50481;
wire x_50482;
wire x_50483;
wire x_50484;
wire x_50485;
wire x_50486;
wire x_50487;
wire x_50488;
wire x_50489;
wire x_50490;
wire x_50491;
wire x_50492;
wire x_50493;
wire x_50494;
wire x_50495;
wire x_50496;
wire x_50497;
wire x_50498;
wire x_50499;
wire x_50500;
wire x_50501;
wire x_50502;
wire x_50503;
wire x_50504;
wire x_50505;
wire x_50506;
wire x_50507;
wire x_50508;
wire x_50509;
wire x_50510;
wire x_50511;
wire x_50512;
wire x_50513;
wire x_50514;
wire x_50515;
wire x_50516;
wire x_50517;
wire x_50518;
wire x_50519;
wire x_50520;
wire x_50521;
wire x_50522;
wire x_50523;
wire x_50524;
wire x_50525;
wire x_50526;
wire x_50527;
wire x_50528;
wire x_50529;
wire x_50530;
wire x_50531;
wire x_50532;
wire x_50533;
wire x_50534;
wire x_50535;
wire x_50536;
wire x_50537;
wire x_50538;
wire x_50539;
wire x_50540;
wire x_50541;
wire x_50542;
wire x_50543;
wire x_50544;
wire x_50545;
wire x_50546;
wire x_50547;
wire x_50548;
wire x_50549;
wire x_50550;
wire x_50551;
wire x_50552;
wire x_50553;
wire x_50554;
wire x_50555;
wire x_50556;
wire x_50557;
wire x_50558;
wire x_50559;
wire x_50560;
wire x_50561;
wire x_50562;
wire x_50563;
wire x_50564;
wire x_50565;
wire x_50566;
wire x_50567;
wire x_50568;
wire x_50569;
wire x_50570;
wire x_50571;
wire x_50572;
wire x_50573;
wire x_50574;
wire x_50575;
wire x_50576;
wire x_50577;
wire x_50578;
wire x_50579;
wire x_50580;
wire x_50581;
wire x_50582;
wire x_50583;
wire x_50584;
wire x_50585;
wire x_50586;
wire x_50587;
wire x_50588;
wire x_50589;
wire x_50590;
wire x_50591;
wire x_50592;
wire x_50593;
wire x_50594;
wire x_50595;
wire x_50596;
wire x_50597;
wire x_50598;
wire x_50599;
wire x_50600;
wire x_50601;
wire x_50602;
wire x_50603;
wire x_50604;
wire x_50605;
wire x_50606;
wire x_50607;
wire x_50608;
wire x_50609;
wire x_50610;
wire x_50611;
wire x_50612;
wire x_50613;
wire x_50614;
wire x_50615;
wire x_50616;
wire x_50617;
wire x_50618;
wire x_50619;
wire x_50620;
wire x_50621;
wire x_50622;
wire x_50623;
wire x_50624;
wire x_50625;
wire x_50626;
wire x_50627;
wire x_50628;
wire x_50629;
wire x_50630;
wire x_50631;
wire x_50632;
wire x_50633;
wire x_50634;
wire x_50635;
wire x_50636;
wire x_50637;
wire x_50638;
wire x_50639;
wire x_50640;
wire x_50641;
wire x_50642;
wire x_50643;
wire x_50644;
wire x_50645;
wire x_50646;
wire x_50647;
wire x_50648;
wire x_50649;
wire x_50650;
wire x_50651;
wire x_50652;
wire x_50653;
wire x_50654;
wire x_50655;
wire x_50656;
wire x_50657;
wire x_50658;
wire x_50659;
wire x_50660;
wire x_50661;
wire x_50662;
wire x_50663;
wire x_50664;
wire x_50665;
wire x_50666;
wire x_50667;
wire x_50668;
wire x_50669;
wire x_50670;
wire x_50671;
wire x_50672;
wire x_50673;
wire x_50674;
wire x_50675;
wire x_50676;
wire x_50677;
wire x_50678;
wire x_50679;
wire x_50680;
wire x_50681;
wire x_50682;
wire x_50683;
wire x_50684;
wire x_50685;
wire x_50686;
wire x_50687;
wire x_50688;
wire x_50689;
wire x_50690;
wire x_50691;
wire x_50692;
wire x_50693;
wire x_50694;
wire x_50695;
wire x_50696;
wire x_50697;
wire x_50698;
wire x_50699;
wire x_50700;
wire x_50701;
wire x_50702;
wire x_50703;
wire x_50704;
wire x_50705;
wire x_50706;
wire x_50707;
wire x_50708;
wire x_50709;
wire x_50710;
wire x_50711;
wire x_50712;
wire x_50713;
wire x_50714;
wire x_50715;
wire x_50716;
wire x_50717;
wire x_50718;
wire x_50719;
wire x_50720;
wire x_50721;
wire x_50722;
wire x_50723;
wire x_50724;
wire x_50725;
wire x_50726;
wire x_50727;
wire x_50728;
wire x_50729;
wire x_50730;
wire x_50731;
wire x_50732;
wire x_50733;
wire x_50734;
wire x_50735;
wire x_50736;
wire x_50737;
wire x_50738;
wire x_50739;
wire x_50740;
wire x_50741;
wire x_50742;
wire x_50743;
wire x_50744;
wire x_50745;
wire x_50746;
wire x_50747;
wire x_50748;
wire x_50749;
wire x_50750;
wire x_50751;
wire x_50752;
wire x_50753;
wire x_50754;
wire x_50755;
wire x_50756;
wire x_50757;
wire x_50758;
wire x_50759;
wire x_50760;
wire x_50761;
wire x_50762;
wire x_50763;
wire x_50764;
wire x_50765;
wire x_50766;
wire x_50767;
wire x_50768;
wire x_50769;
wire x_50770;
wire x_50771;
wire x_50772;
wire x_50773;
wire x_50774;
wire x_50775;
wire x_50776;
wire x_50777;
wire x_50778;
wire x_50779;
wire x_50780;
wire x_50781;
wire x_50782;
wire x_50783;
wire x_50784;
wire x_50785;
wire x_50786;
wire x_50787;
wire x_50788;
wire x_50789;
wire x_50790;
wire x_50791;
wire x_50792;
wire x_50793;
wire x_50794;
wire x_50795;
wire x_50796;
wire x_50797;
wire x_50798;
wire x_50799;
wire x_50800;
wire x_50801;
wire x_50802;
wire x_50803;
wire x_50804;
wire x_50805;
wire x_50806;
wire x_50807;
wire x_50808;
wire x_50809;
wire x_50810;
wire x_50811;
wire x_50812;
wire x_50813;
wire x_50814;
wire x_50815;
wire x_50816;
wire x_50817;
wire x_50818;
wire x_50819;
wire x_50820;
wire x_50821;
wire x_50822;
wire x_50823;
wire x_50824;
wire x_50825;
wire x_50826;
wire x_50827;
wire x_50828;
wire x_50829;
wire x_50830;
wire x_50831;
wire x_50832;
wire x_50833;
wire x_50834;
wire x_50835;
wire x_50836;
wire x_50837;
wire x_50838;
wire x_50839;
wire x_50840;
wire x_50841;
wire x_50842;
wire x_50843;
wire x_50844;
wire x_50845;
wire x_50846;
wire x_50847;
wire x_50848;
wire x_50849;
wire x_50850;
wire x_50851;
wire x_50852;
wire x_50853;
wire x_50854;
wire x_50855;
wire x_50856;
wire x_50857;
wire x_50858;
wire x_50859;
wire x_50860;
wire x_50861;
wire x_50862;
wire x_50863;
wire x_50864;
wire x_50865;
wire x_50866;
wire x_50867;
wire x_50868;
wire x_50869;
wire x_50870;
wire x_50871;
wire x_50872;
wire x_50873;
wire x_50874;
wire x_50875;
wire x_50876;
wire x_50877;
wire x_50878;
wire x_50879;
wire x_50880;
wire x_50881;
wire x_50882;
wire x_50883;
wire x_50884;
wire x_50885;
wire x_50886;
wire x_50887;
wire x_50888;
wire x_50889;
wire x_50890;
wire x_50891;
wire x_50892;
wire x_50893;
wire x_50894;
wire x_50895;
wire x_50896;
wire x_50897;
wire x_50898;
wire x_50899;
wire x_50900;
wire x_50901;
wire x_50902;
wire x_50903;
wire x_50904;
wire x_50905;
wire x_50906;
wire x_50907;
wire x_50908;
wire x_50909;
wire x_50910;
wire x_50911;
wire x_50912;
wire x_50913;
wire x_50914;
wire x_50915;
wire x_50916;
wire x_50917;
wire x_50918;
wire x_50919;
wire x_50920;
wire x_50921;
wire x_50922;
wire x_50923;
wire x_50924;
wire x_50925;
wire x_50926;
wire x_50927;
wire x_50928;
wire x_50929;
wire x_50930;
wire x_50931;
wire x_50932;
wire x_50933;
wire x_50934;
wire x_50935;
wire x_50936;
wire x_50937;
wire x_50938;
wire x_50939;
wire x_50940;
wire x_50941;
wire x_50942;
wire x_50943;
wire x_50944;
wire x_50945;
wire x_50946;
wire x_50947;
wire x_50948;
wire x_50949;
wire x_50950;
wire x_50951;
wire x_50952;
wire x_50953;
wire x_50954;
wire x_50955;
wire x_50956;
wire x_50957;
wire x_50958;
wire x_50959;
wire x_50960;
wire x_50961;
wire x_50962;
wire x_50963;
wire x_50964;
wire x_50965;
wire x_50966;
wire x_50967;
wire x_50968;
wire x_50969;
wire x_50970;
wire x_50971;
wire x_50972;
wire x_50973;
wire x_50974;
wire x_50975;
wire x_50976;
wire x_50977;
wire x_50978;
wire x_50979;
wire x_50980;
wire x_50981;
wire x_50982;
wire x_50983;
wire x_50984;
wire x_50985;
wire x_50986;
wire x_50987;
wire x_50988;
wire x_50989;
wire x_50990;
wire x_50991;
wire x_50992;
wire x_50993;
wire x_50994;
wire x_50995;
wire x_50996;
wire x_50997;
wire x_50998;
wire x_50999;
wire x_51000;
wire x_51001;
wire x_51002;
wire x_51003;
wire x_51004;
wire x_51005;
wire x_51006;
wire x_51007;
wire x_51008;
wire x_51009;
wire x_51010;
wire x_51011;
wire x_51012;
wire x_51013;
wire x_51014;
wire x_51015;
wire x_51016;
wire x_51017;
wire x_51018;
wire x_51019;
wire x_51020;
wire x_51021;
wire x_51022;
wire x_51023;
wire x_51024;
wire x_51025;
wire x_51026;
wire x_51027;
wire x_51028;
wire x_51029;
wire x_51030;
wire x_51031;
wire x_51032;
wire x_51033;
wire x_51034;
wire x_51035;
wire x_51036;
wire x_51037;
wire x_51038;
wire x_51039;
wire x_51040;
wire x_51041;
wire x_51042;
wire x_51043;
wire x_51044;
wire x_51045;
wire x_51046;
wire x_51047;
wire x_51048;
wire x_51049;
wire x_51050;
wire x_51051;
wire x_51052;
wire x_51053;
wire x_51054;
wire x_51055;
wire x_51056;
wire x_51057;
wire x_51058;
wire x_51059;
wire x_51060;
wire x_51061;
wire x_51062;
wire x_51063;
wire x_51064;
wire x_51065;
wire x_51066;
wire x_51067;
wire x_51068;
wire x_51069;
wire x_51070;
wire x_51071;
wire x_51072;
wire x_51073;
wire x_51074;
wire x_51075;
wire x_51076;
wire x_51077;
wire x_51078;
wire x_51079;
wire x_51080;
wire x_51081;
wire x_51082;
wire x_51083;
wire x_51084;
wire x_51085;
wire x_51086;
wire x_51087;
wire x_51088;
wire x_51089;
wire x_51090;
wire x_51091;
wire x_51092;
wire x_51093;
wire x_51094;
wire x_51095;
wire x_51096;
wire x_51097;
wire x_51098;
wire x_51099;
wire x_51100;
wire x_51101;
wire x_51102;
wire x_51103;
wire x_51104;
wire x_51105;
wire x_51106;
wire x_51107;
wire x_51108;
wire x_51109;
wire x_51110;
wire x_51111;
wire x_51112;
wire x_51113;
wire x_51114;
wire x_51115;
wire x_51116;
wire x_51117;
wire x_51118;
wire x_51119;
wire x_51120;
wire x_51121;
wire x_51122;
wire x_51123;
wire x_51124;
wire x_51125;
wire x_51126;
wire x_51127;
wire x_51128;
wire x_51129;
wire x_51130;
wire x_51131;
wire x_51132;
wire x_51133;
wire x_51134;
wire x_51135;
wire x_51136;
wire x_51137;
wire x_51138;
wire x_51139;
wire x_51140;
wire x_51141;
wire x_51142;
wire x_51143;
wire x_51144;
wire x_51145;
wire x_51146;
wire x_51147;
wire x_51148;
wire x_51149;
wire x_51150;
wire x_51151;
wire x_51152;
wire x_51153;
wire x_51154;
wire x_51155;
wire x_51156;
wire x_51157;
wire x_51158;
wire x_51159;
wire x_51160;
wire x_51161;
wire x_51162;
wire x_51163;
wire x_51164;
wire x_51165;
wire x_51166;
wire x_51167;
wire x_51168;
wire x_51169;
wire x_51170;
wire x_51171;
wire x_51172;
wire x_51173;
wire x_51174;
wire x_51175;
wire x_51176;
wire x_51177;
wire x_51178;
wire x_51179;
wire x_51180;
wire x_51181;
wire x_51182;
wire x_51183;
wire x_51184;
wire x_51185;
wire x_51186;
wire x_51187;
wire x_51188;
wire x_51189;
wire x_51190;
wire x_51191;
wire x_51192;
wire x_51193;
wire x_51194;
wire x_51195;
wire x_51196;
wire x_51197;
wire x_51198;
wire x_51199;
wire x_51200;
wire x_51201;
wire x_51202;
wire x_51203;
wire x_51204;
wire x_51205;
wire x_51206;
wire x_51207;
wire x_51208;
wire x_51209;
wire x_51210;
wire x_51211;
wire x_51212;
wire x_51213;
wire x_51214;
wire x_51215;
wire x_51216;
wire x_51217;
wire x_51218;
wire x_51219;
wire x_51220;
wire x_51221;
wire x_51222;
wire x_51223;
wire x_51224;
wire x_51225;
wire x_51226;
wire x_51227;
wire x_51228;
wire x_51229;
wire x_51230;
wire x_51231;
wire x_51232;
wire x_51233;
wire x_51234;
wire x_51235;
wire x_51236;
wire x_51237;
wire x_51238;
wire x_51239;
wire x_51240;
wire x_51241;
wire x_51242;
wire x_51243;
wire x_51244;
wire x_51245;
wire x_51246;
wire x_51247;
wire x_51248;
wire x_51249;
wire x_51250;
wire x_51251;
wire x_51252;
wire x_51253;
wire x_51254;
wire x_51255;
wire x_51256;
wire x_51257;
wire x_51258;
wire x_51259;
wire x_51260;
wire x_51261;
wire x_51262;
wire x_51263;
wire x_51264;
wire x_51265;
wire x_51266;
wire x_51267;
wire x_51268;
wire x_51269;
wire x_51270;
wire x_51271;
wire x_51272;
wire x_51273;
wire x_51274;
wire x_51275;
wire x_51276;
wire x_51277;
wire x_51278;
wire x_51279;
wire x_51280;
wire x_51281;
wire x_51282;
wire x_51283;
wire x_51284;
wire x_51285;
wire x_51286;
wire x_51287;
wire x_51288;
wire x_51289;
wire x_51290;
wire x_51291;
wire x_51292;
wire x_51293;
wire x_51294;
wire x_51295;
wire x_51296;
wire x_51297;
wire x_51298;
wire x_51299;
wire x_51300;
wire x_51301;
wire x_51302;
wire x_51303;
wire x_51304;
wire x_51305;
wire x_51306;
wire x_51307;
wire x_51308;
wire x_51309;
wire x_51310;
wire x_51311;
wire x_51312;
wire x_51313;
wire x_51314;
wire x_51315;
wire x_51316;
wire x_51317;
wire x_51318;
wire x_51319;
wire x_51320;
wire x_51321;
wire x_51322;
wire x_51323;
wire x_51324;
wire x_51325;
wire x_51326;
wire x_51327;
wire x_51328;
wire x_51329;
wire x_51330;
wire x_51331;
wire x_51332;
wire x_51333;
wire x_51334;
wire x_51335;
wire x_51336;
wire x_51337;
wire x_51338;
wire x_51339;
wire x_51340;
wire x_51341;
wire x_51342;
wire x_51343;
wire x_51344;
wire x_51345;
wire x_51346;
wire x_51347;
wire x_51348;
wire x_51349;
wire x_51350;
wire x_51351;
wire x_51352;
wire x_51353;
wire x_51354;
wire x_51355;
wire x_51356;
wire x_51357;
wire x_51358;
wire x_51359;
wire x_51360;
wire x_51361;
wire x_51362;
wire x_51363;
wire x_51364;
wire x_51365;
wire x_51366;
wire x_51367;
wire x_51368;
wire x_51369;
wire x_51370;
wire x_51371;
wire x_51372;
wire x_51373;
wire x_51374;
wire x_51375;
wire x_51376;
wire x_51377;
wire x_51378;
wire x_51379;
wire x_51380;
wire x_51381;
wire x_51382;
wire x_51383;
wire x_51384;
wire x_51385;
wire x_51386;
wire x_51387;
wire x_51388;
wire x_51389;
wire x_51390;
wire x_51391;
wire x_51392;
wire x_51393;
wire x_51394;
wire x_51395;
wire x_51396;
wire x_51397;
wire x_51398;
wire x_51399;
wire x_51400;
wire x_51401;
wire x_51402;
wire x_51403;
wire x_51404;
wire x_51405;
wire x_51406;
wire x_51407;
wire x_51408;
wire x_51409;
wire x_51410;
wire x_51411;
wire x_51412;
wire x_51413;
wire x_51414;
wire x_51415;
wire x_51416;
wire x_51417;
wire x_51418;
wire x_51419;
wire x_51420;
wire x_51421;
wire x_51422;
wire x_51423;
wire x_51424;
wire x_51425;
wire x_51426;
wire x_51427;
wire x_51428;
wire x_51429;
wire x_51430;
wire x_51431;
wire x_51432;
wire x_51433;
wire x_51434;
wire x_51435;
wire x_51436;
wire x_51437;
wire x_51438;
wire x_51439;
wire x_51440;
wire x_51441;
wire x_51442;
wire x_51443;
wire x_51444;
wire x_51445;
wire x_51446;
wire x_51447;
wire x_51448;
wire x_51449;
wire x_51450;
wire x_51451;
wire x_51452;
wire x_51453;
wire x_51454;
wire x_51455;
wire x_51456;
wire x_51457;
wire x_51458;
wire x_51459;
wire x_51460;
wire x_51461;
wire x_51462;
wire x_51463;
wire x_51464;
wire x_51465;
wire x_51466;
wire x_51467;
wire x_51468;
wire x_51469;
wire x_51470;
wire x_51471;
wire x_51472;
wire x_51473;
wire x_51474;
wire x_51475;
wire x_51476;
wire x_51477;
wire x_51478;
wire x_51479;
wire x_51480;
wire x_51481;
wire x_51482;
wire x_51483;
wire x_51484;
wire x_51485;
wire x_51486;
wire x_51487;
wire x_51488;
wire x_51489;
wire x_51490;
wire x_51491;
wire x_51492;
wire x_51493;
wire x_51494;
wire x_51495;
wire x_51496;
wire x_51497;
wire x_51498;
wire x_51499;
wire x_51500;
wire x_51501;
wire x_51502;
wire x_51503;
wire x_51504;
wire x_51505;
wire x_51506;
wire x_51507;
wire x_51508;
wire x_51509;
wire x_51510;
wire x_51511;
wire x_51512;
wire x_51513;
wire x_51514;
wire x_51515;
wire x_51516;
wire x_51517;
wire x_51518;
wire x_51519;
wire x_51520;
wire x_51521;
wire x_51522;
wire x_51523;
wire x_51524;
wire x_51525;
wire x_51526;
wire x_51527;
wire x_51528;
wire x_51529;
wire x_51530;
wire x_51531;
wire x_51532;
wire x_51533;
wire x_51534;
wire x_51535;
wire x_51536;
wire x_51537;
wire x_51538;
wire x_51539;
wire x_51540;
wire x_51541;
wire x_51542;
wire x_51543;
wire x_51544;
wire x_51545;
wire x_51546;
wire x_51547;
wire x_51548;
wire x_51549;
wire x_51550;
wire x_51551;
wire x_51552;
wire x_51553;
wire x_51554;
wire x_51555;
wire x_51556;
wire x_51557;
wire x_51558;
wire x_51559;
wire x_51560;
wire x_51561;
wire x_51562;
wire x_51563;
wire x_51564;
wire x_51565;
wire x_51566;
wire x_51567;
wire x_51568;
wire x_51569;
wire x_51570;
wire x_51571;
wire x_51572;
wire x_51573;
wire x_51574;
wire x_51575;
wire x_51576;
wire x_51577;
wire x_51578;
wire x_51579;
wire x_51580;
wire x_51581;
wire x_51582;
wire x_51583;
wire x_51584;
wire x_51585;
wire x_51586;
wire x_51587;
wire x_51588;
wire x_51589;
wire x_51590;
wire x_51591;
wire x_51592;
wire x_51593;
wire x_51594;
wire x_51595;
wire x_51596;
wire x_51597;
wire x_51598;
wire x_51599;
wire x_51600;
wire x_51601;
wire x_51602;
wire x_51603;
wire x_51604;
wire x_51605;
wire x_51606;
wire x_51607;
wire x_51608;
wire x_51609;
wire x_51610;
wire x_51611;
wire x_51612;
wire x_51613;
wire x_51614;
wire x_51615;
wire x_51616;
wire x_51617;
wire x_51618;
wire x_51619;
wire x_51620;
wire x_51621;
wire x_51622;
wire x_51623;
wire x_51624;
wire x_51625;
wire x_51626;
wire x_51627;
wire x_51628;
wire x_51629;
wire x_51630;
wire x_51631;
wire x_51632;
wire x_51633;
wire x_51634;
wire x_51635;
wire x_51636;
wire x_51637;
wire x_51638;
wire x_51639;
wire x_51640;
wire x_51641;
wire x_51642;
wire x_51643;
wire x_51644;
wire x_51645;
wire x_51646;
wire x_51647;
wire x_51648;
wire x_51649;
wire x_51650;
wire x_51651;
wire x_51652;
wire x_51653;
wire x_51654;
wire x_51655;
wire x_51656;
wire x_51657;
wire x_51658;
wire x_51659;
wire x_51660;
wire x_51661;
wire x_51662;
wire x_51663;
wire x_51664;
wire x_51665;
wire x_51666;
wire x_51667;
wire x_51668;
wire x_51669;
wire x_51670;
wire x_51671;
wire x_51672;
wire x_51673;
wire x_51674;
wire x_51675;
wire x_51676;
wire x_51677;
wire x_51678;
wire x_51679;
wire x_51680;
wire x_51681;
wire x_51682;
wire x_51683;
wire x_51684;
wire x_51685;
wire x_51686;
wire x_51687;
wire x_51688;
wire x_51689;
wire x_51690;
wire x_51691;
wire x_51692;
wire x_51693;
wire x_51694;
wire x_51695;
wire x_51696;
wire x_51697;
wire x_51698;
wire x_51699;
wire x_51700;
wire x_51701;
wire x_51702;
wire x_51703;
wire x_51704;
wire x_51705;
wire x_51706;
wire x_51707;
wire x_51708;
wire x_51709;
wire x_51710;
wire x_51711;
wire x_51712;
wire x_51713;
wire x_51714;
wire x_51715;
wire x_51716;
wire x_51717;
wire x_51718;
wire x_51719;
wire x_51720;
wire x_51721;
wire x_51722;
wire x_51723;
wire x_51724;
wire x_51725;
wire x_51726;
wire x_51727;
wire x_51728;
wire x_51729;
wire x_51730;
wire x_51731;
wire x_51732;
wire x_51733;
wire x_51734;
wire x_51735;
wire x_51736;
wire x_51737;
wire x_51738;
wire x_51739;
wire x_51740;
wire x_51741;
wire x_51742;
wire x_51743;
wire x_51744;
wire x_51745;
wire x_51746;
wire x_51747;
wire x_51748;
wire x_51749;
wire x_51750;
wire x_51751;
wire x_51752;
wire x_51753;
wire x_51754;
wire x_51755;
wire x_51756;
wire x_51757;
wire x_51758;
wire x_51759;
wire x_51760;
wire x_51761;
wire x_51762;
wire x_51763;
wire x_51764;
wire x_51765;
wire x_51766;
wire x_51767;
wire x_51768;
wire x_51769;
wire x_51770;
wire x_51771;
wire x_51772;
wire x_51773;
wire x_51774;
wire x_51775;
wire x_51776;
wire x_51777;
wire x_51778;
wire x_51779;
wire x_51780;
wire x_51781;
wire x_51782;
wire x_51783;
wire x_51784;
wire x_51785;
wire x_51786;
wire x_51787;
wire x_51788;
wire x_51789;
wire x_51790;
wire x_51791;
wire x_51792;
wire x_51793;
wire x_51794;
wire x_51795;
wire x_51796;
wire x_51797;
wire x_51798;
wire x_51799;
wire x_51800;
wire x_51801;
wire x_51802;
wire x_51803;
wire x_51804;
wire x_51805;
wire x_51806;
wire x_51807;
wire x_51808;
wire x_51809;
wire x_51810;
wire x_51811;
wire x_51812;
wire x_51813;
wire x_51814;
wire x_51815;
wire x_51816;
wire x_51817;
wire x_51818;
wire x_51819;
wire x_51820;
wire x_51821;
wire x_51822;
wire x_51823;
wire x_51824;
wire x_51825;
wire x_51826;
wire x_51827;
wire x_51828;
wire x_51829;
wire x_51830;
wire x_51831;
wire x_51832;
wire x_51833;
wire x_51834;
wire x_51835;
wire x_51836;
wire x_51837;
wire x_51838;
wire x_51839;
wire x_51840;
wire x_51841;
wire x_51842;
wire x_51843;
wire x_51844;
wire x_51845;
wire x_51846;
wire x_51847;
wire x_51848;
wire x_51849;
wire x_51850;
wire x_51851;
wire x_51852;
wire x_51853;
wire x_51854;
wire x_51855;
wire x_51856;
wire x_51857;
wire x_51858;
wire x_51859;
wire x_51860;
wire x_51861;
wire x_51862;
wire x_51863;
wire x_51864;
wire x_51865;
wire x_51866;
wire x_51867;
wire x_51868;
wire x_51869;
wire x_51870;
wire x_51871;
wire x_51872;
wire x_51873;
wire x_51874;
wire x_51875;
wire x_51876;
wire x_51877;
wire x_51878;
wire x_51879;
wire x_51880;
wire x_51881;
wire x_51882;
wire x_51883;
wire x_51884;
wire x_51885;
wire x_51886;
wire x_51887;
wire x_51888;
wire x_51889;
wire x_51890;
wire x_51891;
wire x_51892;
wire x_51893;
wire x_51894;
wire x_51895;
wire x_51896;
wire x_51897;
wire x_51898;
wire x_51899;
wire x_51900;
wire x_51901;
wire x_51902;
wire x_51903;
wire x_51904;
wire x_51905;
wire x_51906;
wire x_51907;
wire x_51908;
wire x_51909;
wire x_51910;
wire x_51911;
wire x_51912;
wire x_51913;
wire x_51914;
wire x_51915;
wire x_51916;
wire x_51917;
wire x_51918;
wire x_51919;
wire x_51920;
wire x_51921;
wire x_51922;
wire x_51923;
wire x_51924;
wire x_51925;
wire x_51926;
wire x_51927;
wire x_51928;
wire x_51929;
wire x_51930;
wire x_51931;
wire x_51932;
wire x_51933;
wire x_51934;
wire x_51935;
wire x_51936;
wire x_51937;
wire x_51938;
wire x_51939;
wire x_51940;
wire x_51941;
wire x_51942;
wire x_51943;
wire x_51944;
wire x_51945;
wire x_51946;
wire x_51947;
wire x_51948;
wire x_51949;
wire x_51950;
wire x_51951;
wire x_51952;
wire x_51953;
wire x_51954;
wire x_51955;
wire x_51956;
wire x_51957;
wire x_51958;
wire x_51959;
wire x_51960;
wire x_51961;
wire x_51962;
wire x_51963;
wire x_51964;
wire x_51965;
wire x_51966;
wire x_51967;
wire x_51968;
wire x_51969;
wire x_51970;
wire x_51971;
wire x_51972;
wire x_51973;
wire x_51974;
wire x_51975;
wire x_51976;
wire x_51977;
wire x_51978;
wire x_51979;
wire x_51980;
wire x_51981;
wire x_51982;
wire x_51983;
wire x_51984;
wire x_51985;
wire x_51986;
wire x_51987;
wire x_51988;
wire x_51989;
wire x_51990;
wire x_51991;
wire x_51992;
wire x_51993;
wire x_51994;
wire x_51995;
wire x_51996;
wire x_51997;
wire x_51998;
wire x_51999;
wire x_52000;
wire x_52001;
wire x_52002;
wire x_52003;
wire x_52004;
wire x_52005;
wire x_52006;
wire x_52007;
wire x_52008;
wire x_52009;
wire x_52010;
wire x_52011;
wire x_52012;
wire x_52013;
wire x_52014;
wire x_52015;
wire x_52016;
wire x_52017;
wire x_52018;
wire x_52019;
wire x_52020;
wire x_52021;
wire x_52022;
wire x_52023;
wire x_52024;
wire x_52025;
wire x_52026;
wire x_52027;
wire x_52028;
wire x_52029;
wire x_52030;
wire x_52031;
wire x_52032;
wire x_52033;
wire x_52034;
wire x_52035;
wire x_52036;
wire x_52037;
wire x_52038;
wire x_52039;
wire x_52040;
wire x_52041;
wire x_52042;
wire x_52043;
wire x_52044;
wire x_52045;
wire x_52046;
wire x_52047;
wire x_52048;
wire x_52049;
wire x_52050;
wire x_52051;
wire x_52052;
wire x_52053;
wire x_52054;
wire x_52055;
wire x_52056;
wire x_52057;
wire x_52058;
wire x_52059;
wire x_52060;
wire x_52061;
wire x_52062;
wire x_52063;
wire x_52064;
wire x_52065;
wire x_52066;
wire x_52067;
wire x_52068;
wire x_52069;
wire x_52070;
wire x_52071;
wire x_52072;
wire x_52073;
wire x_52074;
wire x_52075;
wire x_52076;
wire x_52077;
wire x_52078;
wire x_52079;
wire x_52080;
wire x_52081;
wire x_52082;
wire x_52083;
wire x_52084;
wire x_52085;
wire x_52086;
wire x_52087;
wire x_52088;
wire x_52089;
wire x_52090;
wire x_52091;
wire x_52092;
wire x_52093;
wire x_52094;
wire x_52095;
wire x_52096;
wire x_52097;
wire x_52098;
wire x_52099;
wire x_52100;
wire x_52101;
wire x_52102;
wire x_52103;
wire x_52104;
wire x_52105;
wire x_52106;
wire x_52107;
wire x_52108;
wire x_52109;
wire x_52110;
wire x_52111;
wire x_52112;
wire x_52113;
wire x_52114;
wire x_52115;
wire x_52116;
wire x_52117;
wire x_52118;
wire x_52119;
wire x_52120;
wire x_52121;
wire x_52122;
wire x_52123;
wire x_52124;
wire x_52125;
wire x_52126;
wire x_52127;
wire x_52128;
wire x_52129;
wire x_52130;
wire x_52131;
wire x_52132;
wire x_52133;
wire x_52134;
wire x_52135;
wire x_52136;
wire x_52137;
wire x_52138;
wire x_52139;
wire x_52140;
wire x_52141;
wire x_52142;
wire x_52143;
wire x_52144;
wire x_52145;
wire x_52146;
wire x_52147;
wire x_52148;
wire x_52149;
wire x_52150;
wire x_52151;
wire x_52152;
wire x_52153;
wire x_52154;
wire x_52155;
wire x_52156;
wire x_52157;
wire x_52158;
wire x_52159;
wire x_52160;
wire x_52161;
wire x_52162;
wire x_52163;
wire x_52164;
wire x_52165;
wire x_52166;
wire x_52167;
wire x_52168;
wire x_52169;
wire x_52170;
wire x_52171;
wire x_52172;
wire x_52173;
wire x_52174;
wire x_52175;
wire x_52176;
wire x_52177;
wire x_52178;
wire x_52179;
wire x_52180;
wire x_52181;
wire x_52182;
wire x_52183;
wire x_52184;
wire x_52185;
wire x_52186;
wire x_52187;
wire x_52188;
wire x_52189;
wire x_52190;
wire x_52191;
wire x_52192;
wire x_52193;
wire x_52194;
wire x_52195;
wire x_52196;
wire x_52197;
wire x_52198;
wire x_52199;
wire x_52200;
wire x_52201;
wire x_52202;
wire x_52203;
wire x_52204;
wire x_52205;
wire x_52206;
wire x_52207;
wire x_52208;
wire x_52209;
wire x_52210;
wire x_52211;
wire x_52212;
wire x_52213;
wire x_52214;
wire x_52215;
wire x_52216;
wire x_52217;
wire x_52218;
wire x_52219;
wire x_52220;
wire x_52221;
wire x_52222;
wire x_52223;
wire x_52224;
wire x_52225;
wire x_52226;
wire x_52227;
wire x_52228;
wire x_52229;
wire x_52230;
wire x_52231;
wire x_52232;
wire x_52233;
wire x_52234;
wire x_52235;
wire x_52236;
wire x_52237;
wire x_52238;
wire x_52239;
wire x_52240;
wire x_52241;
wire x_52242;
wire x_52243;
wire x_52244;
wire x_52245;
wire x_52246;
wire x_52247;
wire x_52248;
wire x_52249;
wire x_52250;
wire x_52251;
wire x_52252;
wire x_52253;
wire x_52254;
wire x_52255;
wire x_52256;
wire x_52257;
wire x_52258;
wire x_52259;
wire x_52260;
wire x_52261;
wire x_52262;
wire x_52263;
wire x_52264;
wire x_52265;
wire x_52266;
wire x_52267;
wire x_52268;
wire x_52269;
wire x_52270;
wire x_52271;
wire x_52272;
wire x_52273;
wire x_52274;
wire x_52275;
wire x_52276;
wire x_52277;
wire x_52278;
wire x_52279;
wire x_52280;
wire x_52281;
wire x_52282;
wire x_52283;
wire x_52284;
wire x_52285;
wire x_52286;
wire x_52287;
wire x_52288;
wire x_52289;
wire x_52290;
wire x_52291;
wire x_52292;
wire x_52293;
wire x_52294;
wire x_52295;
wire x_52296;
wire x_52297;
wire x_52298;
wire x_52299;
wire x_52300;
wire x_52301;
wire x_52302;
wire x_52303;
wire x_52304;
wire x_52305;
wire x_52306;
wire x_52307;
wire x_52308;
wire x_52309;
wire x_52310;
wire x_52311;
wire x_52312;
wire x_52313;
wire x_52314;
wire x_52315;
wire x_52316;
wire x_52317;
wire x_52318;
wire x_52319;
wire x_52320;
wire x_52321;
wire x_52322;
wire x_52323;
wire x_52324;
wire x_52325;
wire x_52326;
wire x_52327;
wire x_52328;
wire x_52329;
wire x_52330;
wire x_52331;
wire x_52332;
wire x_52333;
wire x_52334;
wire x_52335;
wire x_52336;
wire x_52337;
wire x_52338;
wire x_52339;
wire x_52340;
wire x_52341;
wire x_52342;
wire x_52343;
wire x_52344;
wire x_52345;
wire x_52346;
wire x_52347;
wire x_52348;
wire x_52349;
wire x_52350;
wire x_52351;
wire x_52352;
wire x_52353;
wire x_52354;
wire x_52355;
wire x_52356;
wire x_52357;
wire x_52358;
wire x_52359;
wire x_52360;
wire x_52361;
wire x_52362;
wire x_52363;
wire x_52364;
wire x_52365;
wire x_52366;
wire x_52367;
wire x_52368;
wire x_52369;
wire x_52370;
wire x_52371;
wire x_52372;
wire x_52373;
wire x_52374;
wire x_52375;
wire x_52376;
wire x_52377;
wire x_52378;
wire x_52379;
wire x_52380;
wire x_52381;
wire x_52382;
wire x_52383;
wire x_52384;
wire x_52385;
wire x_52386;
wire x_52387;
wire x_52388;
wire x_52389;
wire x_52390;
wire x_52391;
wire x_52392;
wire x_52393;
wire x_52394;
wire x_52395;
wire x_52396;
wire x_52397;
wire x_52398;
wire x_52399;
wire x_52400;
wire x_52401;
wire x_52402;
wire x_52403;
wire x_52404;
wire x_52405;
wire x_52406;
wire x_52407;
wire x_52408;
wire x_52409;
wire x_52410;
wire x_52411;
wire x_52412;
wire x_52413;
wire x_52414;
wire x_52415;
wire x_52416;
wire x_52417;
wire x_52418;
wire x_52419;
wire x_52420;
wire x_52421;
wire x_52422;
wire x_52423;
wire x_52424;
wire x_52425;
wire x_52426;
wire x_52427;
wire x_52428;
wire x_52429;
wire x_52430;
wire x_52431;
wire x_52432;
wire x_52433;
wire x_52434;
wire x_52435;
wire x_52436;
wire x_52437;
wire x_52438;
wire x_52439;
wire x_52440;
wire x_52441;
wire x_52442;
wire x_52443;
wire x_52444;
wire x_52445;
wire x_52446;
wire x_52447;
wire x_52448;
wire x_52449;
wire x_52450;
wire x_52451;
wire x_52452;
wire x_52453;
wire x_52454;
wire x_52455;
wire x_52456;
wire x_52457;
wire x_52458;
wire x_52459;
wire x_52460;
wire x_52461;
wire x_52462;
wire x_52463;
wire x_52464;
wire x_52465;
wire x_52466;
wire x_52467;
wire x_52468;
wire x_52469;
wire x_52470;
wire x_52471;
wire x_52472;
wire x_52473;
wire x_52474;
wire x_52475;
wire x_52476;
wire x_52477;
wire x_52478;
wire x_52479;
wire x_52480;
wire x_52481;
wire x_52482;
wire x_52483;
wire x_52484;
wire x_52485;
wire x_52486;
wire x_52487;
wire x_52488;
wire x_52489;
wire x_52490;
wire x_52491;
wire x_52492;
wire x_52493;
wire x_52494;
wire x_52495;
wire x_52496;
wire x_52497;
wire x_52498;
wire x_52499;
wire x_52500;
wire x_52501;
wire x_52502;
wire x_52503;
wire x_52504;
wire x_52505;
wire x_52506;
wire x_52507;
wire x_52508;
wire x_52509;
wire x_52510;
wire x_52511;
wire x_52512;
wire x_52513;
wire x_52514;
wire x_52515;
wire x_52516;
wire x_52517;
wire x_52518;
wire x_52519;
wire x_52520;
wire x_52521;
wire x_52522;
wire x_52523;
wire x_52524;
wire x_52525;
wire x_52526;
wire x_52527;
wire x_52528;
wire x_52529;
wire x_52530;
wire x_52531;
wire x_52532;
wire x_52533;
wire x_52534;
wire x_52535;
wire x_52536;
wire x_52537;
wire x_52538;
wire x_52539;
wire x_52540;
wire x_52541;
wire x_52542;
wire x_52543;
wire x_52544;
wire x_52545;
wire x_52546;
wire x_52547;
wire x_52548;
wire x_52549;
wire x_52550;
wire x_52551;
wire x_52552;
wire x_52553;
wire x_52554;
wire x_52555;
wire x_52556;
wire x_52557;
wire x_52558;
wire x_52559;
wire x_52560;
wire x_52561;
wire x_52562;
wire x_52563;
wire x_52564;
wire x_52565;
wire x_52566;
wire x_52567;
wire x_52568;
wire x_52569;
wire x_52570;
wire x_52571;
wire x_52572;
wire x_52573;
wire x_52574;
wire x_52575;
wire x_52576;
wire x_52577;
wire x_52578;
wire x_52579;
wire x_52580;
wire x_52581;
wire x_52582;
wire x_52583;
wire x_52584;
wire x_52585;
wire x_52586;
wire x_52587;
wire x_52588;
wire x_52589;
wire x_52590;
wire x_52591;
wire x_52592;
wire x_52593;
wire x_52594;
wire x_52595;
wire x_52596;
wire x_52597;
wire x_52598;
wire x_52599;
wire x_52600;
wire x_52601;
wire x_52602;
wire x_52603;
wire x_52604;
wire x_52605;
wire x_52606;
wire x_52607;
wire x_52608;
wire x_52609;
wire x_52610;
wire x_52611;
wire x_52612;
wire x_52613;
wire x_52614;
wire x_52615;
wire x_52616;
wire x_52617;
wire x_52618;
wire x_52619;
wire x_52620;
wire x_52621;
wire x_52622;
wire x_52623;
wire x_52624;
wire x_52625;
wire x_52626;
wire x_52627;
wire x_52628;
wire x_52629;
wire x_52630;
wire x_52631;
wire x_52632;
wire x_52633;
wire x_52634;
wire x_52635;
wire x_52636;
wire x_52637;
wire x_52638;
wire x_52639;
wire x_52640;
wire x_52641;
wire x_52642;
wire x_52643;
wire x_52644;
wire x_52645;
wire x_52646;
wire x_52647;
wire x_52648;
wire x_52649;
wire x_52650;
wire x_52651;
wire x_52652;
wire x_52653;
wire x_52654;
wire x_52655;
wire x_52656;
wire x_52657;
wire x_52658;
wire x_52659;
wire x_52660;
wire x_52661;
wire x_52662;
wire x_52663;
wire x_52664;
wire x_52665;
wire x_52666;
wire x_52667;
wire x_52668;
wire x_52669;
wire x_52670;
wire x_52671;
wire x_52672;
wire x_52673;
wire x_52674;
wire x_52675;
wire x_52676;
wire x_52677;
wire x_52678;
wire x_52679;
wire x_52680;
wire x_52681;
wire x_52682;
wire x_52683;
wire x_52684;
wire x_52685;
wire x_52686;
wire x_52687;
wire x_52688;
wire x_52689;
wire x_52690;
wire x_52691;
wire x_52692;
wire x_52693;
wire x_52694;
wire x_52695;
wire x_52696;
wire x_52697;
wire x_52698;
wire x_52699;
wire x_52700;
wire x_52701;
wire x_52702;
wire x_52703;
wire x_52704;
wire x_52705;
wire x_52706;
wire x_52707;
wire x_52708;
wire x_52709;
wire x_52710;
wire x_52711;
wire x_52712;
wire x_52713;
wire x_52714;
wire x_52715;
wire x_52716;
wire x_52717;
wire x_52718;
wire x_52719;
wire x_52720;
wire x_52721;
wire x_52722;
wire x_52723;
wire x_52724;
wire x_52725;
wire x_52726;
wire x_52727;
wire x_52728;
wire x_52729;
wire x_52730;
wire x_52731;
wire x_52732;
wire x_52733;
wire x_52734;
wire x_52735;
wire x_52736;
wire x_52737;
wire x_52738;
wire x_52739;
wire x_52740;
wire x_52741;
wire x_52742;
wire x_52743;
wire x_52744;
wire x_52745;
wire x_52746;
wire x_52747;
wire x_52748;
wire x_52749;
wire x_52750;
wire x_52751;
wire x_52752;
wire x_52753;
wire x_52754;
wire x_52755;
wire x_52756;
wire x_52757;
wire x_52758;
wire x_52759;
wire x_52760;
wire x_52761;
wire x_52762;
wire x_52763;
wire x_52764;
wire x_52765;
wire x_52766;
wire x_52767;
wire x_52768;
wire x_52769;
wire x_52770;
wire x_52771;
wire x_52772;
wire x_52773;
wire x_52774;
wire x_52775;
wire x_52776;
wire x_52777;
wire x_52778;
wire x_52779;
wire x_52780;
wire x_52781;
wire x_52782;
wire x_52783;
wire x_52784;
wire x_52785;
wire x_52786;
wire x_52787;
wire x_52788;
wire x_52789;
wire x_52790;
wire x_52791;
wire x_52792;
wire x_52793;
wire x_52794;
wire x_52795;
wire x_52796;
wire x_52797;
wire x_52798;
wire x_52799;
wire x_52800;
wire x_52801;
wire x_52802;
wire x_52803;
wire x_52804;
wire x_52805;
wire x_52806;
wire x_52807;
wire x_52808;
wire x_52809;
wire x_52810;
wire x_52811;
wire x_52812;
wire x_52813;
wire x_52814;
wire x_52815;
wire x_52816;
wire x_52817;
wire x_52818;
wire x_52819;
wire x_52820;
wire x_52821;
wire x_52822;
wire x_52823;
wire x_52824;
wire x_52825;
wire x_52826;
wire x_52827;
wire x_52828;
wire x_52829;
wire x_52830;
wire x_52831;
wire x_52832;
wire x_52833;
wire x_52834;
wire x_52835;
wire x_52836;
wire x_52837;
wire x_52838;
wire x_52839;
wire x_52840;
wire x_52841;
wire x_52842;
wire x_52843;
wire x_52844;
wire x_52845;
wire x_52846;
wire x_52847;
wire x_52848;
wire x_52849;
wire x_52850;
wire x_52851;
wire x_52852;
wire x_52853;
wire x_52854;
wire x_52855;
wire x_52856;
wire x_52857;
wire x_52858;
wire x_52859;
wire x_52860;
wire x_52861;
wire x_52862;
wire x_52863;
wire x_52864;
wire x_52865;
wire x_52866;
wire x_52867;
wire x_52868;
wire x_52869;
wire x_52870;
wire x_52871;
wire x_52872;
wire x_52873;
wire x_52874;
wire x_52875;
wire x_52876;
wire x_52877;
wire x_52878;
wire x_52879;
wire x_52880;
wire x_52881;
wire x_52882;
wire x_52883;
wire x_52884;
wire x_52885;
wire x_52886;
wire x_52887;
wire x_52888;
wire x_52889;
wire x_52890;
wire x_52891;
wire x_52892;
wire x_52893;
wire x_52894;
wire x_52895;
wire x_52896;
wire x_52897;
wire x_52898;
wire x_52899;
wire x_52900;
wire x_52901;
wire x_52902;
wire x_52903;
wire x_52904;
wire x_52905;
wire x_52906;
wire x_52907;
wire x_52908;
wire x_52909;
wire x_52910;
wire x_52911;
wire x_52912;
wire x_52913;
wire x_52914;
wire x_52915;
wire x_52916;
wire x_52917;
wire x_52918;
wire x_52919;
wire x_52920;
wire x_52921;
wire x_52922;
wire x_52923;
wire x_52924;
wire x_52925;
wire x_52926;
wire x_52927;
wire x_52928;
wire x_52929;
wire x_52930;
wire x_52931;
wire x_52932;
wire x_52933;
wire x_52934;
wire x_52935;
wire x_52936;
wire x_52937;
wire x_52938;
wire x_52939;
wire x_52940;
wire x_52941;
wire x_52942;
wire x_52943;
wire x_52944;
wire x_52945;
wire x_52946;
wire x_52947;
wire x_52948;
wire x_52949;
wire x_52950;
wire x_52951;
wire x_52952;
wire x_52953;
wire x_52954;
wire x_52955;
wire x_52956;
wire x_52957;
wire x_52958;
wire x_52959;
wire x_52960;
wire x_52961;
wire x_52962;
wire x_52963;
wire x_52964;
wire x_52965;
wire x_52966;
wire x_52967;
wire x_52968;
wire x_52969;
wire x_52970;
wire x_52971;
wire x_52972;
wire x_52973;
wire x_52974;
wire x_52975;
wire x_52976;
wire x_52977;
wire x_52978;
wire x_52979;
wire x_52980;
wire x_52981;
wire x_52982;
wire x_52983;
wire x_52984;
wire x_52985;
wire x_52986;
wire x_52987;
wire x_52988;
wire x_52989;
wire x_52990;
wire x_52991;
wire x_52992;
wire x_52993;
wire x_52994;
wire x_52995;
wire x_52996;
wire x_52997;
wire x_52998;
wire x_52999;
wire x_53000;
wire x_53001;
wire x_53002;
wire x_53003;
wire x_53004;
wire x_53005;
wire x_53006;
wire x_53007;
wire x_53008;
wire x_53009;
wire x_53010;
wire x_53011;
wire x_53012;
wire x_53013;
wire x_53014;
wire x_53015;
wire x_53016;
wire x_53017;
wire x_53018;
wire x_53019;
wire x_53020;
wire x_53021;
wire x_53022;
wire x_53023;
wire x_53024;
wire x_53025;
wire x_53026;
wire x_53027;
wire x_53028;
wire x_53029;
wire x_53030;
wire x_53031;
wire x_53032;
wire x_53033;
wire x_53034;
wire x_53035;
wire x_53036;
wire x_53037;
wire x_53038;
wire x_53039;
wire x_53040;
wire x_53041;
wire x_53042;
wire x_53043;
wire x_53044;
wire x_53045;
wire x_53046;
wire x_53047;
wire x_53048;
wire x_53049;
wire x_53050;
wire x_53051;
wire x_53052;
wire x_53053;
wire x_53054;
wire x_53055;
wire x_53056;
wire x_53057;
wire x_53058;
wire x_53059;
wire x_53060;
wire x_53061;
wire x_53062;
wire x_53063;
wire x_53064;
wire x_53065;
wire x_53066;
wire x_53067;
wire x_53068;
wire x_53069;
wire x_53070;
wire x_53071;
wire x_53072;
wire x_53073;
wire x_53074;
wire x_53075;
wire x_53076;
wire x_53077;
wire x_53078;
wire x_53079;
wire x_53080;
wire x_53081;
wire x_53082;
wire x_53083;
wire x_53084;
wire x_53085;
wire x_53086;
wire x_53087;
wire x_53088;
wire x_53089;
wire x_53090;
wire x_53091;
wire x_53092;
wire x_53093;
wire x_53094;
wire x_53095;
wire x_53096;
wire x_53097;
wire x_53098;
wire x_53099;
wire x_53100;
wire x_53101;
wire x_53102;
wire x_53103;
wire x_53104;
wire x_53105;
wire x_53106;
wire x_53107;
wire x_53108;
wire x_53109;
wire x_53110;
wire x_53111;
wire x_53112;
wire x_53113;
wire x_53114;
wire x_53115;
wire x_53116;
wire x_53117;
wire x_53118;
wire x_53119;
wire x_53120;
wire x_53121;
wire x_53122;
wire x_53123;
wire x_53124;
wire x_53125;
wire x_53126;
wire x_53127;
wire x_53128;
wire x_53129;
wire x_53130;
wire x_53131;
wire x_53132;
wire x_53133;
wire x_53134;
wire x_53135;
wire x_53136;
wire x_53137;
wire x_53138;
wire x_53139;
wire x_53140;
wire x_53141;
wire x_53142;
wire x_53143;
wire x_53144;
wire x_53145;
wire x_53146;
wire x_53147;
wire x_53148;
wire x_53149;
wire x_53150;
wire x_53151;
wire x_53152;
wire x_53153;
wire x_53154;
wire x_53155;
wire x_53156;
wire x_53157;
wire x_53158;
wire x_53159;
wire x_53160;
wire x_53161;
wire x_53162;
wire x_53163;
wire x_53164;
wire x_53165;
wire x_53166;
wire x_53167;
wire x_53168;
wire x_53169;
wire x_53170;
wire x_53171;
wire x_53172;
wire x_53173;
wire x_53174;
wire x_53175;
wire x_53176;
wire x_53177;
wire x_53178;
wire x_53179;
wire x_53180;
wire x_53181;
wire x_53182;
wire x_53183;
wire x_53184;
wire x_53185;
wire x_53186;
wire x_53187;
wire x_53188;
wire x_53189;
wire x_53190;
wire x_53191;
wire x_53192;
wire x_53193;
wire x_53194;
wire x_53195;
wire x_53196;
wire x_53197;
wire x_53198;
wire x_53199;
wire x_53200;
wire x_53201;
wire x_53202;
wire x_53203;
wire x_53204;
wire x_53205;
wire x_53206;
wire x_53207;
wire x_53208;
wire x_53209;
wire x_53210;
wire x_53211;
wire x_53212;
wire x_53213;
wire x_53214;
wire x_53215;
wire x_53216;
wire x_53217;
wire x_53218;
wire x_53219;
wire x_53220;
wire x_53221;
wire x_53222;
wire x_53223;
wire x_53224;
wire x_53225;
wire x_53226;
wire x_53227;
wire x_53228;
wire x_53229;
wire x_53230;
wire x_53231;
wire x_53232;
wire x_53233;
wire x_53234;
wire x_53235;
wire x_53236;
wire x_53237;
wire x_53238;
wire x_53239;
wire x_53240;
wire x_53241;
wire x_53242;
wire x_53243;
wire x_53244;
wire x_53245;
wire x_53246;
wire x_53247;
wire x_53248;
wire x_53249;
wire x_53250;
wire x_53251;
wire x_53252;
wire x_53253;
wire x_53254;
wire x_53255;
wire x_53256;
wire x_53257;
wire x_53258;
wire x_53259;
wire x_53260;
wire x_53261;
wire x_53262;
wire x_53263;
wire x_53264;
wire x_53265;
wire x_53266;
wire x_53267;
wire x_53268;
wire x_53269;
wire x_53270;
wire x_53271;
wire x_53272;
wire x_53273;
wire x_53274;
wire x_53275;
wire x_53276;
wire x_53277;
wire x_53278;
wire x_53279;
wire x_53280;
wire x_53281;
wire x_53282;
wire x_53283;
wire x_53284;
wire x_53285;
wire x_53286;
wire x_53287;
wire x_53288;
wire x_53289;
wire x_53290;
wire x_53291;
wire x_53292;
wire x_53293;
wire x_53294;
wire x_53295;
wire x_53296;
wire x_53297;
wire x_53298;
wire x_53299;
wire x_53300;
wire x_53301;
wire x_53302;
wire x_53303;
wire x_53304;
wire x_53305;
wire x_53306;
wire x_53307;
wire x_53308;
wire x_53309;
wire x_53310;
wire x_53311;
wire x_53312;
wire x_53313;
wire x_53314;
wire x_53315;
wire x_53316;
wire x_53317;
wire x_53318;
wire x_53319;
wire x_53320;
wire x_53321;
wire x_53322;
wire x_53323;
wire x_53324;
wire x_53325;
wire x_53326;
wire x_53327;
wire x_53328;
wire x_53329;
wire x_53330;
wire x_53331;
wire x_53332;
wire x_53333;
wire x_53334;
wire x_53335;
wire x_53336;
wire x_53337;
wire x_53338;
wire x_53339;
wire x_53340;
wire x_53341;
wire x_53342;
wire x_53343;
wire x_53344;
wire x_53345;
wire x_53346;
wire x_53347;
wire x_53348;
wire x_53349;
wire x_53350;
wire x_53351;
wire x_53352;
wire x_53353;
wire x_53354;
wire x_53355;
wire x_53356;
wire x_53357;
wire x_53358;
wire x_53359;
wire x_53360;
wire x_53361;
wire x_53362;
wire x_53363;
wire x_53364;
wire x_53365;
wire x_53366;
wire x_53367;
wire x_53368;
wire x_53369;
wire x_53370;
wire x_53371;
wire x_53372;
wire x_53373;
wire x_53374;
wire x_53375;
wire x_53376;
wire x_53377;
wire x_53378;
wire x_53379;
wire x_53380;
wire x_53381;
wire x_53382;
wire x_53383;
wire x_53384;
wire x_53385;
wire x_53386;
wire x_53387;
wire x_53388;
wire x_53389;
wire x_53390;
wire x_53391;
wire x_53392;
wire x_53393;
wire x_53394;
wire x_53395;
wire x_53396;
wire x_53397;
wire x_53398;
wire x_53399;
wire x_53400;
wire x_53401;
wire x_53402;
wire x_53403;
wire x_53404;
wire x_53405;
wire x_53406;
wire x_53407;
wire x_53408;
wire x_53409;
wire x_53410;
wire x_53411;
wire x_53412;
wire x_53413;
wire x_53414;
wire x_53415;
wire x_53416;
wire x_53417;
wire x_53418;
wire x_53419;
wire x_53420;
wire x_53421;
wire x_53422;
wire x_53423;
wire x_53424;
wire x_53425;
wire x_53426;
wire x_53427;
wire x_53428;
wire x_53429;
wire x_53430;
wire x_53431;
wire x_53432;
wire x_53433;
wire x_53434;
wire x_53435;
wire x_53436;
wire x_53437;
wire x_53438;
wire x_53439;
wire x_53440;
wire x_53441;
wire x_53442;
wire x_53443;
wire x_53444;
wire x_53445;
wire x_53446;
wire x_53447;
wire x_53448;
wire x_53449;
wire x_53450;
wire x_53451;
wire x_53452;
wire x_53453;
wire x_53454;
wire x_53455;
wire x_53456;
wire x_53457;
wire x_53458;
wire x_53459;
wire x_53460;
wire x_53461;
wire x_53462;
wire x_53463;
wire x_53464;
wire x_53465;
wire x_53466;
wire x_53467;
wire x_53468;
wire x_53469;
wire x_53470;
wire x_53471;
wire x_53472;
wire x_53473;
wire x_53474;
wire x_53475;
wire x_53476;
wire x_53477;
wire x_53478;
wire x_53479;
wire x_53480;
wire x_53481;
wire x_53482;
wire x_53483;
wire x_53484;
wire x_53485;
wire x_53486;
wire x_53487;
wire x_53488;
wire x_53489;
wire x_53490;
wire x_53491;
wire x_53492;
wire x_53493;
wire x_53494;
wire x_53495;
wire x_53496;
wire x_53497;
wire x_53498;
wire x_53499;
wire x_53500;
wire x_53501;
wire x_53502;
wire x_53503;
wire x_53504;
wire x_53505;
wire x_53506;
wire x_53507;
wire x_53508;
wire x_53509;
wire x_53510;
wire x_53511;
wire x_53512;
wire x_53513;
wire x_53514;
wire x_53515;
wire x_53516;
wire x_53517;
wire x_53518;
wire x_53519;
wire x_53520;
wire x_53521;
wire x_53522;
wire x_53523;
wire x_53524;
wire x_53525;
wire x_53526;
wire x_53527;
wire x_53528;
wire x_53529;
wire x_53530;
wire x_53531;
wire x_53532;
wire x_53533;
wire x_53534;
wire x_53535;
wire x_53536;
wire x_53537;
wire x_53538;
wire x_53539;
wire x_53540;
wire x_53541;
wire x_53542;
wire x_53543;
wire x_53544;
wire x_53545;
wire x_53546;
wire x_53547;
wire x_53548;
wire x_53549;
wire x_53550;
wire x_53551;
wire x_53552;
wire x_53553;
wire x_53554;
wire x_53555;
wire x_53556;
wire x_53557;
wire x_53558;
wire x_53559;
wire x_53560;
wire x_53561;
wire x_53562;
wire x_53563;
wire x_53564;
wire x_53565;
wire x_53566;
wire x_53567;
wire x_53568;
wire x_53569;
wire x_53570;
wire x_53571;
wire x_53572;
wire x_53573;
wire x_53574;
wire x_53575;
wire x_53576;
wire x_53577;
wire x_53578;
wire x_53579;
wire x_53580;
wire x_53581;
wire x_53582;
wire x_53583;
wire x_53584;
wire x_53585;
wire x_53586;
wire x_53587;
wire x_53588;
wire x_53589;
wire x_53590;
wire x_53591;
wire x_53592;
wire x_53593;
wire x_53594;
wire x_53595;
wire x_53596;
wire x_53597;
wire x_53598;
wire x_53599;
wire x_53600;
wire x_53601;
wire x_53602;
wire x_53603;
wire x_53604;
wire x_53605;
wire x_53606;
wire x_53607;
wire x_53608;
wire x_53609;
wire x_53610;
wire x_53611;
wire x_53612;
wire x_53613;
wire x_53614;
wire x_53615;
wire x_53616;
wire x_53617;
wire x_53618;
wire x_53619;
wire x_53620;
wire x_53621;
wire x_53622;
wire x_53623;
wire x_53624;
wire x_53625;
wire x_53626;
wire x_53627;
wire x_53628;
wire x_53629;
wire x_53630;
wire x_53631;
wire x_53632;
wire x_53633;
wire x_53634;
wire x_53635;
wire x_53636;
wire x_53637;
wire x_53638;
wire x_53639;
wire x_53640;
wire x_53641;
wire x_53642;
wire x_53643;
wire x_53644;
wire x_53645;
wire x_53646;
wire x_53647;
wire x_53648;
wire x_53649;
wire x_53650;
wire x_53651;
wire x_53652;
wire x_53653;
wire x_53654;
wire x_53655;
wire x_53656;
wire x_53657;
wire x_53658;
wire x_53659;
wire x_53660;
wire x_53661;
wire x_53662;
wire x_53663;
wire x_53664;
wire x_53665;
wire x_53666;
wire x_53667;
wire x_53668;
wire x_53669;
wire x_53670;
wire x_53671;
wire x_53672;
wire x_53673;
wire x_53674;
wire x_53675;
wire x_53676;
wire x_53677;
wire x_53678;
wire x_53679;
wire x_53680;
wire x_53681;
wire x_53682;
wire x_53683;
wire x_53684;
wire x_53685;
wire x_53686;
wire x_53687;
wire x_53688;
wire x_53689;
wire x_53690;
wire x_53691;
wire x_53692;
wire x_53693;
wire x_53694;
wire x_53695;
wire x_53696;
wire x_53697;
wire x_53698;
wire x_53699;
wire x_53700;
wire x_53701;
wire x_53702;
wire x_53703;
wire x_53704;
wire x_53705;
wire x_53706;
wire x_53707;
wire x_53708;
wire x_53709;
wire x_53710;
wire x_53711;
wire x_53712;
wire x_53713;
wire x_53714;
wire x_53715;
wire x_53716;
wire x_53717;
wire x_53718;
wire x_53719;
wire x_53720;
wire x_53721;
wire x_53722;
wire x_53723;
wire x_53724;
wire x_53725;
wire x_53726;
wire x_53727;
wire x_53728;
wire x_53729;
wire x_53730;
wire x_53731;
wire x_53732;
wire x_53733;
wire x_53734;
wire x_53735;
wire x_53736;
wire x_53737;
wire x_53738;
wire x_53739;
wire x_53740;
wire x_53741;
wire x_53742;
wire x_53743;
wire x_53744;
wire x_53745;
wire x_53746;
wire x_53747;
wire x_53748;
wire x_53749;
wire x_53750;
wire x_53751;
wire x_53752;
wire x_53753;
wire x_53754;
wire x_53755;
wire x_53756;
wire x_53757;
wire x_53758;
wire x_53759;
wire x_53760;
wire x_53761;
wire x_53762;
wire x_53763;
wire x_53764;
wire x_53765;
wire x_53766;
wire x_53767;
wire x_53768;
wire x_53769;
wire x_53770;
wire x_53771;
wire x_53772;
wire x_53773;
wire x_53774;
wire x_53775;
wire x_53776;
wire x_53777;
wire x_53778;
wire x_53779;
wire x_53780;
wire x_53781;
wire x_53782;
wire x_53783;
wire x_53784;
wire x_53785;
wire x_53786;
wire x_53787;
wire x_53788;
wire x_53789;
wire x_53790;
wire x_53791;
wire x_53792;
wire x_53793;
wire x_53794;
wire x_53795;
wire x_53796;
wire x_53797;
wire x_53798;
wire x_53799;
wire x_53800;
wire x_53801;
wire x_53802;
wire x_53803;
wire x_53804;
wire x_53805;
wire x_53806;
wire x_53807;
wire x_53808;
wire x_53809;
wire x_53810;
wire x_53811;
wire x_53812;
wire x_53813;
wire x_53814;
wire x_53815;
wire x_53816;
wire x_53817;
wire x_53818;
wire x_53819;
wire x_53820;
wire x_53821;
wire x_53822;
wire x_53823;
wire x_53824;
wire x_53825;
wire x_53826;
wire x_53827;
wire x_53828;
wire x_53829;
wire x_53830;
wire x_53831;
wire x_53832;
wire x_53833;
wire x_53834;
wire x_53835;
wire x_53836;
wire x_53837;
wire x_53838;
wire x_53839;
wire x_53840;
wire x_53841;
wire x_53842;
wire x_53843;
wire x_53844;
wire x_53845;
wire x_53846;
wire x_53847;
wire x_53848;
wire x_53849;
wire x_53850;
wire x_53851;
wire x_53852;
wire x_53853;
wire x_53854;
wire x_53855;
wire x_53856;
wire x_53857;
wire x_53858;
wire x_53859;
wire x_53860;
wire x_53861;
wire x_53862;
wire x_53863;
wire x_53864;
wire x_53865;
wire x_53866;
wire x_53867;
wire x_53868;
wire x_53869;
wire x_53870;
wire x_53871;
wire x_53872;
wire x_53873;
wire x_53874;
wire x_53875;
wire x_53876;
wire x_53877;
wire x_53878;
wire x_53879;
wire x_53880;
wire x_53881;
wire x_53882;
wire x_53883;
wire x_53884;
wire x_53885;
wire x_53886;
wire x_53887;
wire x_53888;
wire x_53889;
wire x_53890;
wire x_53891;
wire x_53892;
wire x_53893;
wire x_53894;
wire x_53895;
wire x_53896;
wire x_53897;
wire x_53898;
wire x_53899;
wire x_53900;
wire x_53901;
wire x_53902;
wire x_53903;
wire x_53904;
wire x_53905;
wire x_53906;
wire x_53907;
wire x_53908;
wire x_53909;
wire x_53910;
wire x_53911;
wire x_53912;
wire x_53913;
wire x_53914;
wire x_53915;
wire x_53916;
wire x_53917;
wire x_53918;
wire x_53919;
wire x_53920;
wire x_53921;
wire x_53922;
wire x_53923;
wire x_53924;
wire x_53925;
wire x_53926;
wire x_53927;
wire x_53928;
wire x_53929;
wire x_53930;
wire x_53931;
wire x_53932;
wire x_53933;
wire x_53934;
wire x_53935;
wire x_53936;
wire x_53937;
wire x_53938;
wire x_53939;
wire x_53940;
wire x_53941;
wire x_53942;
wire x_53943;
wire x_53944;
wire x_53945;
wire x_53946;
wire x_53947;
wire x_53948;
wire x_53949;
wire x_53950;
wire x_53951;
wire x_53952;
wire x_53953;
wire x_53954;
wire x_53955;
wire x_53956;
wire x_53957;
wire x_53958;
wire x_53959;
wire x_53960;
wire x_53961;
wire x_53962;
wire x_53963;
wire x_53964;
wire x_53965;
wire x_53966;
wire x_53967;
wire x_53968;
wire x_53969;
wire x_53970;
wire x_53971;
wire x_53972;
wire x_53973;
wire x_53974;
wire x_53975;
wire x_53976;
wire x_53977;
wire x_53978;
wire x_53979;
wire x_53980;
wire x_53981;
wire x_53982;
wire x_53983;
wire x_53984;
wire x_53985;
wire x_53986;
wire x_53987;
wire x_53988;
wire x_53989;
wire x_53990;
wire x_53991;
wire x_53992;
wire x_53993;
wire x_53994;
wire x_53995;
wire x_53996;
wire x_53997;
wire x_53998;
wire x_53999;
wire x_54000;
wire x_54001;
wire x_54002;
wire x_54003;
wire x_54004;
wire x_54005;
wire x_54006;
wire x_54007;
wire x_54008;
wire x_54009;
wire x_54010;
wire x_54011;
wire x_54012;
wire x_54013;
wire x_54014;
wire x_54015;
wire x_54016;
wire x_54017;
wire x_54018;
wire x_54019;
wire x_54020;
wire x_54021;
wire x_54022;
wire x_54023;
wire x_54024;
wire x_54025;
wire x_54026;
wire x_54027;
wire x_54028;
wire x_54029;
wire x_54030;
wire x_54031;
wire x_54032;
wire x_54033;
wire x_54034;
wire x_54035;
wire x_54036;
wire x_54037;
wire x_54038;
wire x_54039;
wire x_54040;
wire x_54041;
wire x_54042;
wire x_54043;
wire x_54044;
wire x_54045;
wire x_54046;
wire x_54047;
wire x_54048;
wire x_54049;
wire x_54050;
wire x_54051;
wire x_54052;
wire x_54053;
wire x_54054;
wire x_54055;
wire x_54056;
wire x_54057;
wire x_54058;
wire x_54059;
wire x_54060;
wire x_54061;
wire x_54062;
wire x_54063;
wire x_54064;
wire x_54065;
wire x_54066;
wire x_54067;
wire x_54068;
wire x_54069;
wire x_54070;
wire x_54071;
wire x_54072;
wire x_54073;
wire x_54074;
wire x_54075;
wire x_54076;
wire x_54077;
wire x_54078;
wire x_54079;
wire x_54080;
wire x_54081;
wire x_54082;
wire x_54083;
wire x_54084;
wire x_54085;
wire x_54086;
wire x_54087;
wire x_54088;
wire x_54089;
wire x_54090;
wire x_54091;
wire x_54092;
wire x_54093;
wire x_54094;
wire x_54095;
wire x_54096;
wire x_54097;
wire x_54098;
wire x_54099;
wire x_54100;
wire x_54101;
wire x_54102;
wire x_54103;
wire x_54104;
wire x_54105;
wire x_54106;
wire x_54107;
wire x_54108;
wire x_54109;
wire x_54110;
wire x_54111;
wire x_54112;
wire x_54113;
wire x_54114;
wire x_54115;
wire x_54116;
wire x_54117;
wire x_54118;
wire x_54119;
wire x_54120;
wire x_54121;
wire x_54122;
wire x_54123;
wire x_54124;
wire x_54125;
wire x_54126;
wire x_54127;
wire x_54128;
wire x_54129;
wire x_54130;
wire x_54131;
wire x_54132;
wire x_54133;
wire x_54134;
wire x_54135;
wire x_54136;
wire x_54137;
wire x_54138;
wire x_54139;
wire x_54140;
wire x_54141;
wire x_54142;
wire x_54143;
wire x_54144;
wire x_54145;
wire x_54146;
wire x_54147;
wire x_54148;
wire x_54149;
wire x_54150;
wire x_54151;
wire x_54152;
wire x_54153;
wire x_54154;
wire x_54155;
wire x_54156;
wire x_54157;
wire x_54158;
wire x_54159;
wire x_54160;
wire x_54161;
wire x_54162;
wire x_54163;
wire x_54164;
wire x_54165;
wire x_54166;
wire x_54167;
wire x_54168;
wire x_54169;
wire x_54170;
wire x_54171;
wire x_54172;
wire x_54173;
wire x_54174;
wire x_54175;
wire x_54176;
wire x_54177;
wire x_54178;
wire x_54179;
wire x_54180;
wire x_54181;
wire x_54182;
wire x_54183;
wire x_54184;
wire x_54185;
wire x_54186;
wire x_54187;
wire x_54188;
wire x_54189;
wire x_54190;
wire x_54191;
wire x_54192;
wire x_54193;
wire x_54194;
wire x_54195;
wire x_54196;
wire x_54197;
wire x_54198;
wire x_54199;
wire x_54200;
wire x_54201;
wire x_54202;
wire x_54203;
wire x_54204;
wire x_54205;
wire x_54206;
wire x_54207;
wire x_54208;
wire x_54209;
wire x_54210;
wire x_54211;
wire x_54212;
wire x_54213;
wire x_54214;
wire x_54215;
wire x_54216;
wire x_54217;
wire x_54218;
wire x_54219;
wire x_54220;
wire x_54221;
wire x_54222;
wire x_54223;
wire x_54224;
wire x_54225;
wire x_54226;
wire x_54227;
wire x_54228;
wire x_54229;
wire x_54230;
wire x_54231;
wire x_54232;
wire x_54233;
wire x_54234;
wire x_54235;
wire x_54236;
wire x_54237;
wire x_54238;
wire x_54239;
wire x_54240;
wire x_54241;
wire x_54242;
wire x_54243;
wire x_54244;
wire x_54245;
wire x_54246;
wire x_54247;
wire x_54248;
wire x_54249;
wire x_54250;
wire x_54251;
wire x_54252;
wire x_54253;
wire x_54254;
wire x_54255;
wire x_54256;
wire x_54257;
wire x_54258;
wire x_54259;
wire x_54260;
wire x_54261;
wire x_54262;
wire x_54263;
wire x_54264;
wire x_54265;
wire x_54266;
wire x_54267;
wire x_54268;
wire x_54269;
wire x_54270;
wire x_54271;
wire x_54272;
wire x_54273;
wire x_54274;
wire x_54275;
wire x_54276;
wire x_54277;
wire x_54278;
wire x_54279;
wire x_54280;
wire x_54281;
wire x_54282;
wire x_54283;
wire x_54284;
wire x_54285;
wire x_54286;
wire x_54287;
wire x_54288;
wire x_54289;
wire x_54290;
wire x_54291;
wire x_54292;
wire x_54293;
wire x_54294;
wire x_54295;
wire x_54296;
wire x_54297;
wire x_54298;
wire x_54299;
wire x_54300;
wire x_54301;
wire x_54302;
wire x_54303;
wire x_54304;
wire x_54305;
wire x_54306;
wire x_54307;
wire x_54308;
wire x_54309;
wire x_54310;
wire x_54311;
wire x_54312;
wire x_54313;
wire x_54314;
wire x_54315;
wire x_54316;
wire x_54317;
wire x_54318;
wire x_54319;
wire x_54320;
wire x_54321;
wire x_54322;
wire x_54323;
wire x_54324;
wire x_54325;
wire x_54326;
wire x_54327;
wire x_54328;
wire x_54329;
wire x_54330;
wire x_54331;
wire x_54332;
wire x_54333;
wire x_54334;
wire x_54335;
wire x_54336;
wire x_54337;
wire x_54338;
wire x_54339;
wire x_54340;
wire x_54341;
wire x_54342;
wire x_54343;
wire x_54344;
wire x_54345;
wire x_54346;
wire x_54347;
wire x_54348;
wire x_54349;
wire x_54350;
wire x_54351;
wire x_54352;
wire x_54353;
wire x_54354;
wire x_54355;
wire x_54356;
wire x_54357;
wire x_54358;
wire x_54359;
wire x_54360;
wire x_54361;
wire x_54362;
wire x_54363;
wire x_54364;
wire x_54365;
wire x_54366;
wire x_54367;
wire x_54368;
wire x_54369;
wire x_54370;
wire x_54371;
wire x_54372;
wire x_54373;
wire x_54374;
wire x_54375;
wire x_54376;
wire x_54377;
wire x_54378;
wire x_54379;
wire x_54380;
wire x_54381;
wire x_54382;
wire x_54383;
wire x_54384;
wire x_54385;
wire x_54386;
wire x_54387;
wire x_54388;
wire x_54389;
wire x_54390;
wire x_54391;
wire x_54392;
wire x_54393;
wire x_54394;
wire x_54395;
wire x_54396;
wire x_54397;
wire x_54398;
wire x_54399;
wire x_54400;
wire x_54401;
wire x_54402;
wire x_54403;
wire x_54404;
wire x_54405;
wire x_54406;
wire x_54407;
wire x_54408;
wire x_54409;
wire x_54410;
wire x_54411;
wire x_54412;
wire x_54413;
wire x_54414;
wire x_54415;
wire x_54416;
wire x_54417;
wire x_54418;
wire x_54419;
wire x_54420;
wire x_54421;
wire x_54422;
wire x_54423;
wire x_54424;
wire x_54425;
wire x_54426;
wire x_54427;
wire x_54428;
wire x_54429;
wire x_54430;
wire x_54431;
wire x_54432;
wire x_54433;
wire x_54434;
wire x_54435;
wire x_54436;
wire x_54437;
wire x_54438;
wire x_54439;
wire x_54440;
wire x_54441;
wire x_54442;
wire x_54443;
wire x_54444;
wire x_54445;
wire x_54446;
wire x_54447;
wire x_54448;
wire x_54449;
wire x_54450;
wire x_54451;
wire x_54452;
wire x_54453;
wire x_54454;
wire x_54455;
wire x_54456;
wire x_54457;
wire x_54458;
wire x_54459;
wire x_54460;
wire x_54461;
wire x_54462;
wire x_54463;
wire x_54464;
wire x_54465;
wire x_54466;
wire x_54467;
wire x_54468;
wire x_54469;
wire x_54470;
wire x_54471;
wire x_54472;
wire x_54473;
wire x_54474;
wire x_54475;
wire x_54476;
wire x_54477;
wire x_54478;
wire x_54479;
wire x_54480;
wire x_54481;
wire x_54482;
wire x_54483;
wire x_54484;
wire x_54485;
wire x_54486;
wire x_54487;
wire x_54488;
wire x_54489;
wire x_54490;
wire x_54491;
wire x_54492;
wire x_54493;
wire x_54494;
wire x_54495;
wire x_54496;
wire x_54497;
wire x_54498;
wire x_54499;
wire x_54500;
wire x_54501;
wire x_54502;
wire x_54503;
wire x_54504;
wire x_54505;
wire x_54506;
wire x_54507;
wire x_54508;
wire x_54509;
wire x_54510;
wire x_54511;
wire x_54512;
wire x_54513;
wire x_54514;
wire x_54515;
wire x_54516;
wire x_54517;
wire x_54518;
wire x_54519;
wire x_54520;
wire x_54521;
wire x_54522;
wire x_54523;
wire x_54524;
wire x_54525;
wire x_54526;
wire x_54527;
wire x_54528;
wire x_54529;
wire x_54530;
wire x_54531;
wire x_54532;
wire x_54533;
wire x_54534;
wire x_54535;
wire x_54536;
wire x_54537;
wire x_54538;
wire x_54539;
wire x_54540;
wire x_54541;
wire x_54542;
wire x_54543;
wire x_54544;
wire x_54545;
wire x_54546;
wire x_54547;
wire x_54548;
wire x_54549;
wire x_54550;
wire x_54551;
wire x_54552;
wire x_54553;
wire x_54554;
wire x_54555;
wire x_54556;
wire x_54557;
wire x_54558;
wire x_54559;
wire x_54560;
wire x_54561;
wire x_54562;
wire x_54563;
wire x_54564;
wire x_54565;
wire x_54566;
wire x_54567;
wire x_54568;
wire x_54569;
wire x_54570;
wire x_54571;
wire x_54572;
wire x_54573;
wire x_54574;
wire x_54575;
wire x_54576;
wire x_54577;
wire x_54578;
wire x_54579;
wire x_54580;
wire x_54581;
wire x_54582;
wire x_54583;
wire x_54584;
wire x_54585;
wire x_54586;
wire x_54587;
wire x_54588;
wire x_54589;
wire x_54590;
wire x_54591;
wire x_54592;
wire x_54593;
wire x_54594;
wire x_54595;
wire x_54596;
wire x_54597;
wire x_54598;
wire x_54599;
wire x_54600;
wire x_54601;
wire x_54602;
wire x_54603;
wire x_54604;
wire x_54605;
wire x_54606;
wire x_54607;
wire x_54608;
wire x_54609;
wire x_54610;
wire x_54611;
wire x_54612;
wire x_54613;
wire x_54614;
wire x_54615;
wire x_54616;
wire x_54617;
wire x_54618;
wire x_54619;
wire x_54620;
wire x_54621;
wire x_54622;
wire x_54623;
wire x_54624;
wire x_54625;
wire x_54626;
wire x_54627;
wire x_54628;
wire x_54629;
wire x_54630;
wire x_54631;
wire x_54632;
wire x_54633;
wire x_54634;
wire x_54635;
wire x_54636;
wire x_54637;
wire x_54638;
wire x_54639;
wire x_54640;
wire x_54641;
wire x_54642;
wire x_54643;
wire x_54644;
wire x_54645;
wire x_54646;
wire x_54647;
wire x_54648;
wire x_54649;
wire x_54650;
wire x_54651;
wire x_54652;
wire x_54653;
wire x_54654;
wire x_54655;
wire x_54656;
wire x_54657;
wire x_54658;
wire x_54659;
wire x_54660;
wire x_54661;
wire x_54662;
wire x_54663;
wire x_54664;
wire x_54665;
wire x_54666;
wire x_54667;
wire x_54668;
wire x_54669;
wire x_54670;
wire x_54671;
wire x_54672;
wire x_54673;
wire x_54674;
wire x_54675;
wire x_54676;
wire x_54677;
wire x_54678;
wire x_54679;
wire x_54680;
wire x_54681;
wire x_54682;
wire x_54683;
wire x_54684;
wire x_54685;
wire x_54686;
wire x_54687;
wire x_54688;
wire x_54689;
wire x_54690;
wire x_54691;
wire x_54692;
wire x_54693;
wire x_54694;
wire x_54695;
wire x_54696;
wire x_54697;
wire x_54698;
wire x_54699;
wire x_54700;
wire x_54701;
wire x_54702;
wire x_54703;
wire x_54704;
wire x_54705;
wire x_54706;
wire x_54707;
wire x_54708;
wire x_54709;
wire x_54710;
wire x_54711;
wire x_54712;
wire x_54713;
wire x_54714;
wire x_54715;
wire x_54716;
wire x_54717;
wire x_54718;
wire x_54719;
wire x_54720;
wire x_54721;
wire x_54722;
wire x_54723;
wire x_54724;
wire x_54725;
wire x_54726;
wire x_54727;
wire x_54728;
wire x_54729;
wire x_54730;
wire x_54731;
wire x_54732;
wire x_54733;
wire x_54734;
wire x_54735;
wire x_54736;
wire x_54737;
wire x_54738;
wire x_54739;
wire x_54740;
wire x_54741;
wire x_54742;
wire x_54743;
wire x_54744;
wire x_54745;
wire x_54746;
wire x_54747;
wire x_54748;
wire x_54749;
wire x_54750;
wire x_54751;
wire x_54752;
wire x_54753;
wire x_54754;
wire x_54755;
wire x_54756;
wire x_54757;
wire x_54758;
wire x_54759;
wire x_54760;
wire x_54761;
wire x_54762;
wire x_54763;
wire x_54764;
wire x_54765;
wire x_54766;
wire x_54767;
wire x_54768;
wire x_54769;
wire x_54770;
wire x_54771;
wire x_54772;
wire x_54773;
wire x_54774;
wire x_54775;
wire x_54776;
wire x_54777;
wire x_54778;
wire x_54779;
wire x_54780;
wire x_54781;
wire x_54782;
wire x_54783;
wire x_54784;
wire x_54785;
wire x_54786;
wire x_54787;
wire x_54788;
wire x_54789;
wire x_54790;
wire x_54791;
wire x_54792;
wire x_54793;
wire x_54794;
wire x_54795;
wire x_54796;
wire x_54797;
wire x_54798;
wire x_54799;
wire x_54800;
wire x_54801;
wire x_54802;
wire x_54803;
wire x_54804;
wire x_54805;
wire x_54806;
wire x_54807;
wire x_54808;
wire x_54809;
wire x_54810;
wire x_54811;
wire x_54812;
wire x_54813;
wire x_54814;
wire x_54815;
wire x_54816;
wire x_54817;
wire x_54818;
wire x_54819;
wire x_54820;
wire x_54821;
wire x_54822;
wire x_54823;
wire x_54824;
wire x_54825;
wire x_54826;
wire x_54827;
wire x_54828;
wire x_54829;
wire x_54830;
wire x_54831;
wire x_54832;
wire x_54833;
wire x_54834;
wire x_54835;
wire x_54836;
wire x_54837;
wire x_54838;
wire x_54839;
wire x_54840;
wire x_54841;
wire x_54842;
wire x_54843;
wire x_54844;
wire x_54845;
wire x_54846;
wire x_54847;
wire x_54848;
wire x_54849;
wire x_54850;
wire x_54851;
wire x_54852;
wire x_54853;
wire x_54854;
wire x_54855;
wire x_54856;
wire x_54857;
wire x_54858;
wire x_54859;
wire x_54860;
wire x_54861;
wire x_54862;
wire x_54863;
wire x_54864;
wire x_54865;
wire x_54866;
wire x_54867;
wire x_54868;
wire x_54869;
wire x_54870;
wire x_54871;
wire x_54872;
wire x_54873;
wire x_54874;
wire x_54875;
wire x_54876;
wire x_54877;
wire x_54878;
wire x_54879;
wire x_54880;
wire x_54881;
wire x_54882;
wire x_54883;
wire x_54884;
wire x_54885;
wire x_54886;
wire x_54887;
wire x_54888;
wire x_54889;
wire x_54890;
wire x_54891;
wire x_54892;
wire x_54893;
wire x_54894;
wire x_54895;
wire x_54896;
wire x_54897;
wire x_54898;
wire x_54899;
wire x_54900;
wire x_54901;
wire x_54902;
wire x_54903;
wire x_54904;
wire x_54905;
wire x_54906;
wire x_54907;
wire x_54908;
wire x_54909;
wire x_54910;
wire x_54911;
wire x_54912;
wire x_54913;
wire x_54914;
wire x_54915;
wire x_54916;
wire x_54917;
wire x_54918;
wire x_54919;
wire x_54920;
wire x_54921;
wire x_54922;
wire x_54923;
wire x_54924;
wire x_54925;
wire x_54926;
wire x_54927;
wire x_54928;
wire x_54929;
wire x_54930;
wire x_54931;
wire x_54932;
wire x_54933;
wire x_54934;
wire x_54935;
wire x_54936;
wire x_54937;
wire x_54938;
wire x_54939;
wire x_54940;
wire x_54941;
wire x_54942;
wire x_54943;
wire x_54944;
wire x_54945;
wire x_54946;
wire x_54947;
wire x_54948;
wire x_54949;
wire x_54950;
wire x_54951;
wire x_54952;
wire x_54953;
wire x_54954;
wire x_54955;
wire x_54956;
wire x_54957;
wire x_54958;
wire x_54959;
wire x_54960;
wire x_54961;
wire x_54962;
wire x_54963;
wire x_54964;
wire x_54965;
wire x_54966;
wire x_54967;
wire x_54968;
wire x_54969;
wire x_54970;
wire x_54971;
wire x_54972;
wire x_54973;
wire x_54974;
wire x_54975;
wire x_54976;
wire x_54977;
wire x_54978;
wire x_54979;
wire x_54980;
wire x_54981;
wire x_54982;
wire x_54983;
wire x_54984;
wire x_54985;
wire x_54986;
wire x_54987;
wire x_54988;
wire x_54989;
wire x_54990;
wire x_54991;
wire x_54992;
wire x_54993;
wire x_54994;
wire x_54995;
wire x_54996;
wire x_54997;
wire x_54998;
wire x_54999;
wire x_55000;
wire x_55001;
wire x_55002;
wire x_55003;
wire x_55004;
wire x_55005;
wire x_55006;
wire x_55007;
wire x_55008;
wire x_55009;
wire x_55010;
wire x_55011;
wire x_55012;
wire x_55013;
wire x_55014;
wire x_55015;
wire x_55016;
wire x_55017;
wire x_55018;
wire x_55019;
wire x_55020;
wire x_55021;
wire x_55022;
wire x_55023;
wire x_55024;
wire x_55025;
wire x_55026;
wire x_55027;
wire x_55028;
wire x_55029;
wire x_55030;
wire x_55031;
wire x_55032;
wire x_55033;
wire x_55034;
wire x_55035;
wire x_55036;
wire x_55037;
wire x_55038;
wire x_55039;
wire x_55040;
wire x_55041;
wire x_55042;
wire x_55043;
wire x_55044;
wire x_55045;
wire x_55046;
wire x_55047;
wire x_55048;
wire x_55049;
wire x_55050;
wire x_55051;
wire x_55052;
wire x_55053;
wire x_55054;
wire x_55055;
wire x_55056;
wire x_55057;
wire x_55058;
wire x_55059;
wire x_55060;
wire x_55061;
wire x_55062;
wire x_55063;
wire x_55064;
wire x_55065;
wire x_55066;
wire x_55067;
wire x_55068;
wire x_55069;
wire x_55070;
wire x_55071;
wire x_55072;
wire x_55073;
wire x_55074;
wire x_55075;
wire x_55076;
wire x_55077;
wire x_55078;
wire x_55079;
wire x_55080;
wire x_55081;
wire x_55082;
wire x_55083;
wire x_55084;
wire x_55085;
wire x_55086;
wire x_55087;
wire x_55088;
wire x_55089;
wire x_55090;
wire x_55091;
wire x_55092;
wire x_55093;
wire x_55094;
wire x_55095;
wire x_55096;
wire x_55097;
wire x_55098;
wire x_55099;
wire x_55100;
wire x_55101;
wire x_55102;
wire x_55103;
wire x_55104;
wire x_55105;
wire x_55106;
wire x_55107;
wire x_55108;
wire x_55109;
wire x_55110;
wire x_55111;
wire x_55112;
wire x_55113;
wire x_55114;
wire x_55115;
wire x_55116;
wire x_55117;
wire x_55118;
wire x_55119;
wire x_55120;
wire x_55121;
wire x_55122;
wire x_55123;
wire x_55124;
wire x_55125;
wire x_55126;
wire x_55127;
wire x_55128;
wire x_55129;
wire x_55130;
wire x_55131;
wire x_55132;
wire x_55133;
wire x_55134;
wire x_55135;
wire x_55136;
wire x_55137;
wire x_55138;
wire x_55139;
wire x_55140;
wire x_55141;
wire x_55142;
wire x_55143;
wire x_55144;
wire x_55145;
wire x_55146;
wire x_55147;
wire x_55148;
wire x_55149;
wire x_55150;
wire x_55151;
wire x_55152;
wire x_55153;
wire x_55154;
wire x_55155;
wire x_55156;
wire x_55157;
wire x_55158;
wire x_55159;
wire x_55160;
wire x_55161;
wire x_55162;
wire x_55163;
wire x_55164;
wire x_55165;
wire x_55166;
wire x_55167;
wire x_55168;
wire x_55169;
wire x_55170;
wire x_55171;
wire x_55172;
wire x_55173;
wire x_55174;
wire x_55175;
wire x_55176;
wire x_55177;
wire x_55178;
wire x_55179;
wire x_55180;
wire x_55181;
wire x_55182;
wire x_55183;
wire x_55184;
wire x_55185;
wire x_55186;
wire x_55187;
wire x_55188;
wire x_55189;
wire x_55190;
wire x_55191;
wire x_55192;
wire x_55193;
wire x_55194;
wire x_55195;
wire x_55196;
wire x_55197;
wire x_55198;
wire x_55199;
wire x_55200;
wire x_55201;
wire x_55202;
wire x_55203;
wire x_55204;
wire x_55205;
wire x_55206;
wire x_55207;
wire x_55208;
wire x_55209;
wire x_55210;
wire x_55211;
wire x_55212;
wire x_55213;
wire x_55214;
wire x_55215;
wire x_55216;
wire x_55217;
wire x_55218;
wire x_55219;
wire x_55220;
wire x_55221;
wire x_55222;
wire x_55223;
wire x_55224;
wire x_55225;
wire x_55226;
wire x_55227;
wire x_55228;
wire x_55229;
wire x_55230;
wire x_55231;
wire x_55232;
wire x_55233;
wire x_55234;
wire x_55235;
wire x_55236;
wire x_55237;
wire x_55238;
wire x_55239;
wire x_55240;
wire x_55241;
wire x_55242;
wire x_55243;
wire x_55244;
wire x_55245;
wire x_55246;
wire x_55247;
wire x_55248;
wire x_55249;
wire x_55250;
wire x_55251;
wire x_55252;
wire x_55253;
wire x_55254;
wire x_55255;
wire x_55256;
wire x_55257;
wire x_55258;
wire x_55259;
wire x_55260;
wire x_55261;
wire x_55262;
wire x_55263;
wire x_55264;
wire x_55265;
wire x_55266;
wire x_55267;
wire x_55268;
wire x_55269;
wire x_55270;
wire x_55271;
wire x_55272;
wire x_55273;
wire x_55274;
wire x_55275;
wire x_55276;
wire x_55277;
wire x_55278;
wire x_55279;
wire x_55280;
wire x_55281;
wire x_55282;
wire x_55283;
wire x_55284;
wire x_55285;
wire x_55286;
wire x_55287;
wire x_55288;
wire x_55289;
wire x_55290;
wire x_55291;
wire x_55292;
wire x_55293;
wire x_55294;
wire x_55295;
wire x_55296;
wire x_55297;
wire x_55298;
wire x_55299;
wire x_55300;
wire x_55301;
wire x_55302;
wire x_55303;
wire x_55304;
wire x_55305;
wire x_55306;
wire x_55307;
wire x_55308;
wire x_55309;
wire x_55310;
wire x_55311;
wire x_55312;
wire x_55313;
wire x_55314;
wire x_55315;
wire x_55316;
wire x_55317;
wire x_55318;
wire x_55319;
wire x_55320;
wire x_55321;
wire x_55322;
wire x_55323;
wire x_55324;
wire x_55325;
wire x_55326;
wire x_55327;
wire x_55328;
wire x_55329;
wire x_55330;
wire x_55331;
wire x_55332;
wire x_55333;
wire x_55334;
wire x_55335;
wire x_55336;
wire x_55337;
wire x_55338;
wire x_55339;
wire x_55340;
wire x_55341;
wire x_55342;
wire x_55343;
wire x_55344;
wire x_55345;
wire x_55346;
wire x_55347;
wire x_55348;
wire x_55349;
wire x_55350;
wire x_55351;
wire x_55352;
wire x_55353;
wire x_55354;
wire x_55355;
wire x_55356;
wire x_55357;
wire x_55358;
wire x_55359;
wire x_55360;
wire x_55361;
wire x_55362;
wire x_55363;
wire x_55364;
wire x_55365;
wire x_55366;
wire x_55367;
wire x_55368;
wire x_55369;
wire x_55370;
wire x_55371;
wire x_55372;
wire x_55373;
wire x_55374;
wire x_55375;
wire x_55376;
wire x_55377;
wire x_55378;
wire x_55379;
wire x_55380;
wire x_55381;
wire x_55382;
wire x_55383;
wire x_55384;
wire x_55385;
wire x_55386;
wire x_55387;
wire x_55388;
wire x_55389;
wire x_55390;
wire x_55391;
wire x_55392;
wire x_55393;
wire x_55394;
wire x_55395;
wire x_55396;
wire x_55397;
wire x_55398;
wire x_55399;
wire x_55400;
wire x_55401;
wire x_55402;
wire x_55403;
wire x_55404;
wire x_55405;
wire x_55406;
wire x_55407;
wire x_55408;
wire x_55409;
wire x_55410;
wire x_55411;
wire x_55412;
wire x_55413;
wire x_55414;
wire x_55415;
wire x_55416;
wire x_55417;
wire x_55418;
wire x_55419;
wire x_55420;
wire x_55421;
wire x_55422;
wire x_55423;
wire x_55424;
wire x_55425;
wire x_55426;
wire x_55427;
wire x_55428;
wire x_55429;
wire x_55430;
wire x_55431;
wire x_55432;
wire x_55433;
wire x_55434;
wire x_55435;
wire x_55436;
wire x_55437;
wire x_55438;
wire x_55439;
wire x_55440;
wire x_55441;
wire x_55442;
wire x_55443;
wire x_55444;
wire x_55445;
wire x_55446;
wire x_55447;
wire x_55448;
wire x_55449;
wire x_55450;
wire x_55451;
wire x_55452;
wire x_55453;
wire x_55454;
wire x_55455;
wire x_55456;
wire x_55457;
wire x_55458;
wire x_55459;
wire x_55460;
wire x_55461;
wire x_55462;
wire x_55463;
wire x_55464;
wire x_55465;
wire x_55466;
wire x_55467;
wire x_55468;
wire x_55469;
wire x_55470;
wire x_55471;
wire x_55472;
wire x_55473;
wire x_55474;
wire x_55475;
wire x_55476;
wire x_55477;
wire x_55478;
wire x_55479;
wire x_55480;
wire x_55481;
wire x_55482;
wire x_55483;
wire x_55484;
wire x_55485;
wire x_55486;
wire x_55487;
wire x_55488;
wire x_55489;
wire x_55490;
wire x_55491;
wire x_55492;
wire x_55493;
wire x_55494;
wire x_55495;
wire x_55496;
wire x_55497;
wire x_55498;
wire x_55499;
wire x_55500;
wire x_55501;
wire x_55502;
wire x_55503;
wire x_55504;
wire x_55505;
wire x_55506;
wire x_55507;
wire x_55508;
wire x_55509;
wire x_55510;
wire x_55511;
wire x_55512;
wire x_55513;
wire x_55514;
wire x_55515;
wire x_55516;
wire x_55517;
wire x_55518;
wire x_55519;
wire x_55520;
wire x_55521;
wire x_55522;
wire x_55523;
wire x_55524;
wire x_55525;
wire x_55526;
wire x_55527;
wire x_55528;
wire x_55529;
wire x_55530;
wire x_55531;
wire x_55532;
wire x_55533;
wire x_55534;
wire x_55535;
wire x_55536;
wire x_55537;
wire x_55538;
wire x_55539;
wire x_55540;
wire x_55541;
wire x_55542;
wire x_55543;
wire x_55544;
wire x_55545;
wire x_55546;
wire x_55547;
wire x_55548;
wire x_55549;
wire x_55550;
wire x_55551;
wire x_55552;
wire x_55553;
wire x_55554;
wire x_55555;
wire x_55556;
wire x_55557;
wire x_55558;
wire x_55559;
wire x_55560;
wire x_55561;
wire x_55562;
wire x_55563;
wire x_55564;
wire x_55565;
wire x_55566;
wire x_55567;
wire x_55568;
wire x_55569;
wire x_55570;
wire x_55571;
wire x_55572;
wire x_55573;
wire x_55574;
wire x_55575;
wire x_55576;
wire x_55577;
wire x_55578;
wire x_55579;
wire x_55580;
wire x_55581;
wire x_55582;
wire x_55583;
wire x_55584;
wire x_55585;
wire x_55586;
wire x_55587;
wire x_55588;
wire x_55589;
wire x_55590;
wire x_55591;
wire x_55592;
wire x_55593;
wire x_55594;
wire x_55595;
wire x_55596;
wire x_55597;
wire x_55598;
wire x_55599;
wire x_55600;
wire x_55601;
wire x_55602;
wire x_55603;
wire x_55604;
wire x_55605;
wire x_55606;
wire x_55607;
wire x_55608;
wire x_55609;
wire x_55610;
wire x_55611;
wire x_55612;
wire x_55613;
wire x_55614;
wire x_55615;
wire x_55616;
wire x_55617;
wire x_55618;
wire x_55619;
wire x_55620;
wire x_55621;
wire x_55622;
wire x_55623;
wire x_55624;
wire x_55625;
wire x_55626;
wire x_55627;
wire x_55628;
wire x_55629;
wire x_55630;
wire x_55631;
wire x_55632;
wire x_55633;
wire x_55634;
wire x_55635;
wire x_55636;
wire x_55637;
wire x_55638;
wire x_55639;
wire x_55640;
wire x_55641;
wire x_55642;
wire x_55643;
wire x_55644;
wire x_55645;
wire x_55646;
wire x_55647;
wire x_55648;
wire x_55649;
wire x_55650;
wire x_55651;
wire x_55652;
wire x_55653;
wire x_55654;
wire x_55655;
wire x_55656;
wire x_55657;
wire x_55658;
wire x_55659;
wire x_55660;
wire x_55661;
wire x_55662;
wire x_55663;
wire x_55664;
wire x_55665;
wire x_55666;
wire x_55667;
wire x_55668;
wire x_55669;
wire x_55670;
wire x_55671;
wire x_55672;
wire x_55673;
wire x_55674;
wire x_55675;
wire x_55676;
wire x_55677;
wire x_55678;
wire x_55679;
wire x_55680;
wire x_55681;
wire x_55682;
wire x_55683;
wire x_55684;
wire x_55685;
wire x_55686;
wire x_55687;
wire x_55688;
wire x_55689;
wire x_55690;
wire x_55691;
wire x_55692;
wire x_55693;
wire x_55694;
wire x_55695;
wire x_55696;
wire x_55697;
wire x_55698;
wire x_55699;
wire x_55700;
wire x_55701;
wire x_55702;
wire x_55703;
wire x_55704;
wire x_55705;
wire x_55706;
wire x_55707;
wire x_55708;
wire x_55709;
wire x_55710;
wire x_55711;
wire x_55712;
wire x_55713;
wire x_55714;
wire x_55715;
wire x_55716;
wire x_55717;
wire x_55718;
wire x_55719;
wire x_55720;
wire x_55721;
wire x_55722;
wire x_55723;
wire x_55724;
wire x_55725;
wire x_55726;
wire x_55727;
wire x_55728;
wire x_55729;
wire x_55730;
wire x_55731;
wire x_55732;
wire x_55733;
wire x_55734;
wire x_55735;
wire x_55736;
wire x_55737;
wire x_55738;
wire x_55739;
wire x_55740;
wire x_55741;
wire x_55742;
wire x_55743;
wire x_55744;
wire x_55745;
wire x_55746;
wire x_55747;
wire x_55748;
wire x_55749;
wire x_55750;
wire x_55751;
wire x_55752;
wire x_55753;
wire x_55754;
wire x_55755;
wire x_55756;
wire x_55757;
wire x_55758;
wire x_55759;
wire x_55760;
wire x_55761;
wire x_55762;
wire x_55763;
wire x_55764;
wire x_55765;
wire x_55766;
wire x_55767;
wire x_55768;
wire x_55769;
wire x_55770;
wire x_55771;
wire x_55772;
wire x_55773;
wire x_55774;
wire x_55775;
wire x_55776;
wire x_55777;
wire x_55778;
wire x_55779;
wire x_55780;
wire x_55781;
wire x_55782;
wire x_55783;
wire x_55784;
wire x_55785;
wire x_55786;
wire x_55787;
wire x_55788;
wire x_55789;
wire x_55790;
wire x_55791;
wire x_55792;
wire x_55793;
wire x_55794;
wire x_55795;
wire x_55796;
wire x_55797;
wire x_55798;
wire x_55799;
wire x_55800;
wire x_55801;
wire x_55802;
wire x_55803;
wire x_55804;
wire x_55805;
wire x_55806;
wire x_55807;
wire x_55808;
wire x_55809;
wire x_55810;
wire x_55811;
wire x_55812;
wire x_55813;
wire x_55814;
wire x_55815;
wire x_55816;
wire x_55817;
wire x_55818;
wire x_55819;
wire x_55820;
wire x_55821;
wire x_55822;
wire x_55823;
wire x_55824;
wire x_55825;
wire x_55826;
wire x_55827;
wire x_55828;
wire x_55829;
wire x_55830;
wire x_55831;
wire x_55832;
wire x_55833;
wire x_55834;
wire x_55835;
wire x_55836;
wire x_55837;
wire x_55838;
wire x_55839;
wire x_55840;
wire x_55841;
wire x_55842;
wire x_55843;
wire x_55844;
wire x_55845;
wire x_55846;
wire x_55847;
wire x_55848;
wire x_55849;
wire x_55850;
wire x_55851;
wire x_55852;
wire x_55853;
wire x_55854;
wire x_55855;
wire x_55856;
wire x_55857;
wire x_55858;
wire x_55859;
wire x_55860;
wire x_55861;
wire x_55862;
wire x_55863;
wire x_55864;
wire x_55865;
wire x_55866;
wire x_55867;
wire x_55868;
wire x_55869;
wire x_55870;
wire x_55871;
wire x_55872;
wire x_55873;
wire x_55874;
wire x_55875;
wire x_55876;
wire x_55877;
wire x_55878;
wire x_55879;
wire x_55880;
wire x_55881;
wire x_55882;
wire x_55883;
wire x_55884;
wire x_55885;
wire x_55886;
wire x_55887;
wire x_55888;
wire x_55889;
wire x_55890;
wire x_55891;
wire x_55892;
wire x_55893;
wire x_55894;
wire x_55895;
wire x_55896;
wire x_55897;
wire x_55898;
wire x_55899;
wire x_55900;
wire x_55901;
wire x_55902;
wire x_55903;
wire x_55904;
wire x_55905;
wire x_55906;
wire x_55907;
wire x_55908;
wire x_55909;
wire x_55910;
wire x_55911;
wire x_55912;
wire x_55913;
wire x_55914;
wire x_55915;
wire x_55916;
wire x_55917;
wire x_55918;
wire x_55919;
wire x_55920;
wire x_55921;
wire x_55922;
wire x_55923;
wire x_55924;
wire x_55925;
wire x_55926;
wire x_55927;
wire x_55928;
wire x_55929;
wire x_55930;
wire x_55931;
wire x_55932;
wire x_55933;
wire x_55934;
wire x_55935;
wire x_55936;
wire x_55937;
wire x_55938;
wire x_55939;
wire x_55940;
wire x_55941;
wire x_55942;
wire x_55943;
wire x_55944;
wire x_55945;
wire x_55946;
wire x_55947;
wire x_55948;
wire x_55949;
wire x_55950;
wire x_55951;
wire x_55952;
wire x_55953;
wire x_55954;
wire x_55955;
wire x_55956;
wire x_55957;
wire x_55958;
wire x_55959;
wire x_55960;
wire x_55961;
wire x_55962;
wire x_55963;
wire x_55964;
wire x_55965;
wire x_55966;
wire x_55967;
wire x_55968;
wire x_55969;
wire x_55970;
wire x_55971;
wire x_55972;
wire x_55973;
wire x_55974;
wire x_55975;
wire x_55976;
wire x_55977;
wire x_55978;
wire x_55979;
wire x_55980;
wire x_55981;
wire x_55982;
wire x_55983;
wire x_55984;
wire x_55985;
wire x_55986;
wire x_55987;
wire x_55988;
wire x_55989;
wire x_55990;
wire x_55991;
wire x_55992;
wire x_55993;
wire x_55994;
wire x_55995;
wire x_55996;
wire x_55997;
wire x_55998;
wire x_55999;
wire x_56000;
wire x_56001;
wire x_56002;
wire x_56003;
wire x_56004;
wire x_56005;
wire x_56006;
wire x_56007;
wire x_56008;
wire x_56009;
wire x_56010;
wire x_56011;
wire x_56012;
wire x_56013;
wire x_56014;
wire x_56015;
wire x_56016;
wire x_56017;
wire x_56018;
wire x_56019;
wire x_56020;
wire x_56021;
wire x_56022;
wire x_56023;
wire x_56024;
wire x_56025;
wire x_56026;
wire x_56027;
wire x_56028;
wire x_56029;
wire x_56030;
wire x_56031;
wire x_56032;
wire x_56033;
wire x_56034;
wire x_56035;
wire x_56036;
wire x_56037;
wire x_56038;
wire x_56039;
wire x_56040;
wire x_56041;
wire x_56042;
wire x_56043;
wire x_56044;
wire x_56045;
wire x_56046;
wire x_56047;
wire x_56048;
wire x_56049;
wire x_56050;
wire x_56051;
wire x_56052;
wire x_56053;
wire x_56054;
wire x_56055;
wire x_56056;
wire x_56057;
wire x_56058;
wire x_56059;
wire x_56060;
wire x_56061;
wire x_56062;
wire x_56063;
wire x_56064;
wire x_56065;
wire x_56066;
wire x_56067;
wire x_56068;
wire x_56069;
wire x_56070;
wire x_56071;
wire x_56072;
wire x_56073;
wire x_56074;
wire x_56075;
wire x_56076;
wire x_56077;
wire x_56078;
wire x_56079;
wire x_56080;
wire x_56081;
wire x_56082;
wire x_56083;
wire x_56084;
wire x_56085;
wire x_56086;
wire x_56087;
wire x_56088;
wire x_56089;
wire x_56090;
wire x_56091;
wire x_56092;
wire x_56093;
wire x_56094;
wire x_56095;
wire x_56096;
wire x_56097;
wire x_56098;
wire x_56099;
wire x_56100;
wire x_56101;
wire x_56102;
wire x_56103;
wire x_56104;
wire x_56105;
wire x_56106;
wire x_56107;
wire x_56108;
wire x_56109;
wire x_56110;
wire x_56111;
wire x_56112;
wire x_56113;
wire x_56114;
wire x_56115;
wire x_56116;
wire x_56117;
wire x_56118;
wire x_56119;
wire x_56120;
wire x_56121;
wire x_56122;
wire x_56123;
wire x_56124;
wire x_56125;
wire x_56126;
wire x_56127;
wire x_56128;
wire x_56129;
wire x_56130;
wire x_56131;
wire x_56132;
wire x_56133;
wire x_56134;
wire x_56135;
wire x_56136;
wire x_56137;
wire x_56138;
wire x_56139;
wire x_56140;
wire x_56141;
wire x_56142;
wire x_56143;
wire x_56144;
wire x_56145;
wire x_56146;
wire x_56147;
wire x_56148;
wire x_56149;
wire x_56150;
wire x_56151;
wire x_56152;
wire x_56153;
wire x_56154;
wire x_56155;
wire x_56156;
wire x_56157;
wire x_56158;
wire x_56159;
wire x_56160;
wire x_56161;
wire x_56162;
wire x_56163;
wire x_56164;
wire x_56165;
wire x_56166;
wire x_56167;
wire x_56168;
wire x_56169;
wire x_56170;
wire x_56171;
wire x_56172;
wire x_56173;
wire x_56174;
wire x_56175;
wire x_56176;
wire x_56177;
wire x_56178;
wire x_56179;
wire x_56180;
wire x_56181;
wire x_56182;
wire x_56183;
wire x_56184;
wire x_56185;
wire x_56186;
wire x_56187;
wire x_56188;
wire x_56189;
wire x_56190;
wire x_56191;
wire x_56192;
wire x_56193;
wire x_56194;
wire x_56195;
wire x_56196;
wire x_56197;
wire x_56198;
wire x_56199;
wire x_56200;
wire x_56201;
wire x_56202;
wire x_56203;
wire x_56204;
wire x_56205;
wire x_56206;
wire x_56207;
wire x_56208;
wire x_56209;
wire x_56210;
wire x_56211;
wire x_56212;
wire x_56213;
wire x_56214;
wire x_56215;
wire x_56216;
wire x_56217;
wire x_56218;
wire x_56219;
wire x_56220;
wire x_56221;
wire x_56222;
wire x_56223;
wire x_56224;
wire x_56225;
wire x_56226;
wire x_56227;
wire x_56228;
wire x_56229;
wire x_56230;
wire x_56231;
wire x_56232;
wire x_56233;
wire x_56234;
wire x_56235;
wire x_56236;
wire x_56237;
wire x_56238;
wire x_56239;
wire x_56240;
wire x_56241;
wire x_56242;
wire x_56243;
wire x_56244;
wire x_56245;
wire x_56246;
wire x_56247;
wire x_56248;
wire x_56249;
wire x_56250;
wire x_56251;
wire x_56252;
wire x_56253;
wire x_56254;
wire x_56255;
wire x_56256;
wire x_56257;
wire x_56258;
wire x_56259;
wire x_56260;
wire x_56261;
wire x_56262;
wire x_56263;
wire x_56264;
wire x_56265;
wire x_56266;
wire x_56267;
wire x_56268;
wire x_56269;
wire x_56270;
wire x_56271;
wire x_56272;
wire x_56273;
wire x_56274;
wire x_56275;
wire x_56276;
wire x_56277;
wire x_56278;
wire x_56279;
wire x_56280;
wire x_56281;
wire x_56282;
wire x_56283;
wire x_56284;
wire x_56285;
wire x_56286;
wire x_56287;
wire x_56288;
wire x_56289;
wire x_56290;
wire x_56291;
wire x_56292;
wire x_56293;
wire x_56294;
wire x_56295;
wire x_56296;
wire x_56297;
wire x_56298;
wire x_56299;
wire x_56300;
wire x_56301;
wire x_56302;
wire x_56303;
wire x_56304;
wire x_56305;
wire x_56306;
wire x_56307;
wire x_56308;
wire x_56309;
wire x_56310;
wire x_56311;
wire x_56312;
wire x_56313;
wire x_56314;
wire x_56315;
wire x_56316;
wire x_56317;
wire x_56318;
wire x_56319;
wire x_56320;
wire x_56321;
wire x_56322;
wire x_56323;
wire x_56324;
wire x_56325;
wire x_56326;
wire x_56327;
wire x_56328;
wire x_56329;
wire x_56330;
wire x_56331;
wire x_56332;
wire x_56333;
wire x_56334;
wire x_56335;
wire x_56336;
wire x_56337;
wire x_56338;
wire x_56339;
wire x_56340;
wire x_56341;
wire x_56342;
wire x_56343;
wire x_56344;
wire x_56345;
wire x_56346;
wire x_56347;
wire x_56348;
wire x_56349;
wire x_56350;
wire x_56351;
wire x_56352;
wire x_56353;
wire x_56354;
wire x_56355;
wire x_56356;
wire x_56357;
wire x_56358;
wire x_56359;
wire x_56360;
wire x_56361;
wire x_56362;
wire x_56363;
wire x_56364;
wire x_56365;
wire x_56366;
wire x_56367;
wire x_56368;
wire x_56369;
wire x_56370;
wire x_56371;
wire x_56372;
wire x_56373;
wire x_56374;
wire x_56375;
wire x_56376;
wire x_56377;
wire x_56378;
wire x_56379;
wire x_56380;
wire x_56381;
wire x_56382;
wire x_56383;
wire x_56384;
wire x_56385;
wire x_56386;
wire x_56387;
wire x_56388;
wire x_56389;
wire x_56390;
wire x_56391;
wire x_56392;
wire x_56393;
wire x_56394;
wire x_56395;
wire x_56396;
wire x_56397;
wire x_56398;
wire x_56399;
wire x_56400;
wire x_56401;
wire x_56402;
wire x_56403;
wire x_56404;
wire x_56405;
wire x_56406;
wire x_56407;
wire x_56408;
wire x_56409;
wire x_56410;
wire x_56411;
wire x_56412;
wire x_56413;
wire x_56414;
wire x_56415;
wire x_56416;
wire x_56417;
wire x_56418;
wire x_56419;
wire x_56420;
wire x_56421;
wire x_56422;
wire x_56423;
wire x_56424;
wire x_56425;
wire x_56426;
wire x_56427;
wire x_56428;
wire x_56429;
wire x_56430;
wire x_56431;
wire x_56432;
wire x_56433;
wire x_56434;
wire x_56435;
wire x_56436;
wire x_56437;
wire x_56438;
wire x_56439;
wire x_56440;
wire x_56441;
wire x_56442;
wire x_56443;
wire x_56444;
wire x_56445;
wire x_56446;
wire x_56447;
wire x_56448;
wire x_56449;
wire x_56450;
wire x_56451;
wire x_56452;
wire x_56453;
wire x_56454;
wire x_56455;
wire x_56456;
wire x_56457;
wire x_56458;
wire x_56459;
wire x_56460;
wire x_56461;
wire x_56462;
wire x_56463;
wire x_56464;
wire x_56465;
wire x_56466;
wire x_56467;
wire x_56468;
wire x_56469;
wire x_56470;
wire x_56471;
wire x_56472;
wire x_56473;
wire x_56474;
wire x_56475;
wire x_56476;
wire x_56477;
wire x_56478;
wire x_56479;
wire x_56480;
wire x_56481;
wire x_56482;
wire x_56483;
wire x_56484;
wire x_56485;
wire x_56486;
wire x_56487;
wire x_56488;
wire x_56489;
wire x_56490;
wire x_56491;
wire x_56492;
wire x_56493;
wire x_56494;
wire x_56495;
wire x_56496;
wire x_56497;
wire x_56498;
wire x_56499;
wire x_56500;
wire x_56501;
wire x_56502;
wire x_56503;
wire x_56504;
wire x_56505;
wire x_56506;
wire x_56507;
wire x_56508;
wire x_56509;
wire x_56510;
wire x_56511;
wire x_56512;
wire x_56513;
wire x_56514;
wire x_56515;
wire x_56516;
wire x_56517;
wire x_56518;
wire x_56519;
wire x_56520;
wire x_56521;
wire x_56522;
wire x_56523;
wire x_56524;
wire x_56525;
wire x_56526;
wire x_56527;
wire x_56528;
wire x_56529;
wire x_56530;
wire x_56531;
wire x_56532;
wire x_56533;
wire x_56534;
wire x_56535;
wire x_56536;
wire x_56537;
wire x_56538;
wire x_56539;
wire x_56540;
wire x_56541;
wire x_56542;
wire x_56543;
wire x_56544;
wire x_56545;
wire x_56546;
wire x_56547;
wire x_56548;
wire x_56549;
wire x_56550;
wire x_56551;
wire x_56552;
wire x_56553;
wire x_56554;
wire x_56555;
wire x_56556;
wire x_56557;
wire x_56558;
wire x_56559;
wire x_56560;
wire x_56561;
wire x_56562;
wire x_56563;
wire x_56564;
wire x_56565;
wire x_56566;
wire x_56567;
wire x_56568;
wire x_56569;
wire x_56570;
wire x_56571;
wire x_56572;
wire x_56573;
wire x_56574;
wire x_56575;
wire x_56576;
wire x_56577;
wire x_56578;
wire x_56579;
wire x_56580;
wire x_56581;
wire x_56582;
wire x_56583;
wire x_56584;
wire x_56585;
wire x_56586;
wire x_56587;
wire x_56588;
wire x_56589;
wire x_56590;
wire x_56591;
wire x_56592;
wire x_56593;
wire x_56594;
wire x_56595;
wire x_56596;
wire x_56597;
wire x_56598;
wire x_56599;
wire x_56600;
wire x_56601;
wire x_56602;
wire x_56603;
wire x_56604;
wire x_56605;
wire x_56606;
wire x_56607;
wire x_56608;
wire x_56609;
wire x_56610;
wire x_56611;
wire x_56612;
wire x_56613;
wire x_56614;
wire x_56615;
wire x_56616;
wire x_56617;
wire x_56618;
wire x_56619;
wire x_56620;
wire x_56621;
wire x_56622;
wire x_56623;
wire x_56624;
wire x_56625;
wire x_56626;
wire x_56627;
wire x_56628;
wire x_56629;
wire x_56630;
wire x_56631;
wire x_56632;
wire x_56633;
wire x_56634;
wire x_56635;
wire x_56636;
wire x_56637;
wire x_56638;
wire x_56639;
wire x_56640;
wire x_56641;
wire x_56642;
wire x_56643;
wire x_56644;
wire x_56645;
wire x_56646;
wire x_56647;
wire x_56648;
wire x_56649;
wire x_56650;
wire x_56651;
wire x_56652;
wire x_56653;
wire x_56654;
wire x_56655;
wire x_56656;
wire x_56657;
wire x_56658;
wire x_56659;
wire x_56660;
wire x_56661;
wire x_56662;
wire x_56663;
wire x_56664;
wire x_56665;
wire x_56666;
wire x_56667;
wire x_56668;
wire x_56669;
wire x_56670;
wire x_56671;
wire x_56672;
wire x_56673;
wire x_56674;
wire x_56675;
wire x_56676;
wire x_56677;
wire x_56678;
wire x_56679;
wire x_56680;
wire x_56681;
wire x_56682;
wire x_56683;
wire x_56684;
wire x_56685;
wire x_56686;
wire x_56687;
wire x_56688;
wire x_56689;
wire x_56690;
wire x_56691;
wire x_56692;
wire x_56693;
wire x_56694;
wire x_56695;
wire x_56696;
wire x_56697;
wire x_56698;
wire x_56699;
wire x_56700;
wire x_56701;
wire x_56702;
wire x_56703;
wire x_56704;
wire x_56705;
wire x_56706;
wire x_56707;
wire x_56708;
wire x_56709;
wire x_56710;
wire x_56711;
wire x_56712;
wire x_56713;
wire x_56714;
wire x_56715;
wire x_56716;
wire x_56717;
wire x_56718;
wire x_56719;
wire x_56720;
wire x_56721;
wire x_56722;
wire x_56723;
wire x_56724;
wire x_56725;
wire x_56726;
wire x_56727;
wire x_56728;
wire x_56729;
wire x_56730;
wire x_56731;
wire x_56732;
wire x_56733;
wire x_56734;
wire x_56735;
wire x_56736;
wire x_56737;
wire x_56738;
wire x_56739;
wire x_56740;
wire x_56741;
wire x_56742;
wire x_56743;
wire x_56744;
wire x_56745;
wire x_56746;
wire x_56747;
wire x_56748;
wire x_56749;
wire x_56750;
wire x_56751;
wire x_56752;
wire x_56753;
wire x_56754;
wire x_56755;
wire x_56756;
wire x_56757;
wire x_56758;
wire x_56759;
wire x_56760;
wire x_56761;
wire x_56762;
wire x_56763;
wire x_56764;
wire x_56765;
wire x_56766;
wire x_56767;
wire x_56768;
wire x_56769;
wire x_56770;
wire x_56771;
wire x_56772;
wire x_56773;
wire x_56774;
wire x_56775;
wire x_56776;
wire x_56777;
wire x_56778;
wire x_56779;
wire x_56780;
wire x_56781;
wire x_56782;
wire x_56783;
wire x_56784;
wire x_56785;
wire x_56786;
wire x_56787;
wire x_56788;
wire x_56789;
wire x_56790;
wire x_56791;
wire x_56792;
wire x_56793;
wire x_56794;
wire x_56795;
wire x_56796;
wire x_56797;
wire x_56798;
wire x_56799;
wire x_56800;
wire x_56801;
wire x_56802;
wire x_56803;
wire x_56804;
wire x_56805;
wire x_56806;
wire x_56807;
wire x_56808;
wire x_56809;
wire x_56810;
wire x_56811;
wire x_56812;
wire x_56813;
wire x_56814;
wire x_56815;
wire x_56816;
wire x_56817;
wire x_56818;
wire x_56819;
wire x_56820;
wire x_56821;
wire x_56822;
wire x_56823;
wire x_56824;
wire x_56825;
wire x_56826;
wire x_56827;
wire x_56828;
wire x_56829;
wire x_56830;
wire x_56831;
wire x_56832;
wire x_56833;
wire x_56834;
wire x_56835;
wire x_56836;
wire x_56837;
wire x_56838;
wire x_56839;
wire x_56840;
wire x_56841;
wire x_56842;
wire x_56843;
wire x_56844;
wire x_56845;
wire x_56846;
wire x_56847;
wire x_56848;
wire x_56849;
wire x_56850;
wire x_56851;
wire x_56852;
wire x_56853;
wire x_56854;
wire x_56855;
wire x_56856;
wire x_56857;
wire x_56858;
wire x_56859;
wire x_56860;
wire x_56861;
wire x_56862;
wire x_56863;
wire x_56864;
wire x_56865;
wire x_56866;
wire x_56867;
wire x_56868;
wire x_56869;
wire x_56870;
wire x_56871;
wire x_56872;
wire x_56873;
wire x_56874;
wire x_56875;
wire x_56876;
wire x_56877;
wire x_56878;
wire x_56879;
wire x_56880;
wire x_56881;
wire x_56882;
wire x_56883;
wire x_56884;
wire x_56885;
wire x_56886;
wire x_56887;
wire x_56888;
wire x_56889;
wire x_56890;
wire x_56891;
wire x_56892;
wire x_56893;
wire x_56894;
wire x_56895;
wire x_56896;
wire x_56897;
wire x_56898;
wire x_56899;
wire x_56900;
wire x_56901;
wire x_56902;
wire x_56903;
wire x_56904;
wire x_56905;
wire x_56906;
wire x_56907;
wire x_56908;
wire x_56909;
wire x_56910;
wire x_56911;
wire x_56912;
wire x_56913;
wire x_56914;
wire x_56915;
wire x_56916;
wire x_56917;
wire x_56918;
wire x_56919;
wire x_56920;
wire x_56921;
wire x_56922;
wire x_56923;
wire x_56924;
wire x_56925;
wire x_56926;
wire x_56927;
wire x_56928;
wire x_56929;
wire x_56930;
wire x_56931;
wire x_56932;
wire x_56933;
wire x_56934;
wire x_56935;
wire x_56936;
wire x_56937;
wire x_56938;
wire x_56939;
wire x_56940;
wire x_56941;
wire x_56942;
wire x_56943;
wire x_56944;
wire x_56945;
wire x_56946;
wire x_56947;
wire x_56948;
wire x_56949;
wire x_56950;
wire x_56951;
wire x_56952;
wire x_56953;
wire x_56954;
wire x_56955;
wire x_56956;
wire x_56957;
wire x_56958;
wire x_56959;
wire x_56960;
wire x_56961;
wire x_56962;
wire x_56963;
wire x_56964;
wire x_56965;
wire x_56966;
wire x_56967;
wire x_56968;
wire x_56969;
wire x_56970;
wire x_56971;
wire x_56972;
wire x_56973;
wire x_56974;
wire x_56975;
wire x_56976;
wire x_56977;
wire x_56978;
wire x_56979;
wire x_56980;
wire x_56981;
wire x_56982;
wire x_56983;
wire x_56984;
wire x_56985;
wire x_56986;
wire x_56987;
wire x_56988;
wire x_56989;
wire x_56990;
wire x_56991;
wire x_56992;
wire x_56993;
wire x_56994;
wire x_56995;
wire x_56996;
wire x_56997;
wire x_56998;
wire x_56999;
wire x_57000;
wire x_57001;
wire x_57002;
wire x_57003;
wire x_57004;
wire x_57005;
wire x_57006;
wire x_57007;
wire x_57008;
wire x_57009;
wire x_57010;
wire x_57011;
wire x_57012;
wire x_57013;
wire x_57014;
wire x_57015;
wire x_57016;
wire x_57017;
wire x_57018;
wire x_57019;
wire x_57020;
wire x_57021;
wire x_57022;
wire x_57023;
wire x_57024;
wire x_57025;
wire x_57026;
wire x_57027;
wire x_57028;
wire x_57029;
wire x_57030;
wire x_57031;
wire x_57032;
wire x_57033;
wire x_57034;
wire x_57035;
wire x_57036;
wire x_57037;
wire x_57038;
wire x_57039;
wire x_57040;
wire x_57041;
wire x_57042;
wire x_57043;
wire x_57044;
wire x_57045;
wire x_57046;
wire x_57047;
wire x_57048;
wire x_57049;
wire x_57050;
wire x_57051;
wire x_57052;
wire x_57053;
wire x_57054;
wire x_57055;
wire x_57056;
wire x_57057;
wire x_57058;
wire x_57059;
wire x_57060;
wire x_57061;
wire x_57062;
wire x_57063;
wire x_57064;
wire x_57065;
wire x_57066;
wire x_57067;
wire x_57068;
wire x_57069;
wire x_57070;
wire x_57071;
wire x_57072;
wire x_57073;
wire x_57074;
wire x_57075;
wire x_57076;
wire x_57077;
wire x_57078;
wire x_57079;
wire x_57080;
wire x_57081;
wire x_57082;
wire x_57083;
wire x_57084;
wire x_57085;
wire x_57086;
wire x_57087;
wire x_57088;
wire x_57089;
wire x_57090;
wire x_57091;
wire x_57092;
wire x_57093;
wire x_57094;
wire x_57095;
wire x_57096;
wire x_57097;
wire x_57098;
wire x_57099;
wire x_57100;
wire x_57101;
wire x_57102;
wire x_57103;
wire x_57104;
wire x_57105;
wire x_57106;
wire x_57107;
wire x_57108;
wire x_57109;
wire x_57110;
wire x_57111;
wire x_57112;
wire x_57113;
wire x_57114;
wire x_57115;
wire x_57116;
wire x_57117;
wire x_57118;
wire x_57119;
wire x_57120;
wire x_57121;
wire x_57122;
wire x_57123;
wire x_57124;
wire x_57125;
wire x_57126;
wire x_57127;
wire x_57128;
wire x_57129;
wire x_57130;
wire x_57131;
wire x_57132;
wire x_57133;
wire x_57134;
wire x_57135;
wire x_57136;
wire x_57137;
wire x_57138;
wire x_57139;
wire x_57140;
wire x_57141;
wire x_57142;
wire x_57143;
wire x_57144;
wire x_57145;
wire x_57146;
wire x_57147;
wire x_57148;
wire x_57149;
wire x_57150;
wire x_57151;
wire x_57152;
wire x_57153;
wire x_57154;
wire x_57155;
wire x_57156;
wire x_57157;
wire x_57158;
wire x_57159;
wire x_57160;
wire x_57161;
wire x_57162;
wire x_57163;
wire x_57164;
wire x_57165;
wire x_57166;
wire x_57167;
wire x_57168;
wire x_57169;
wire x_57170;
wire x_57171;
wire x_57172;
wire x_57173;
wire x_57174;
wire x_57175;
wire x_57176;
wire x_57177;
wire x_57178;
wire x_57179;
wire x_57180;
wire x_57181;
wire x_57182;
wire x_57183;
wire x_57184;
wire x_57185;
wire x_57186;
wire x_57187;
wire x_57188;
wire x_57189;
wire x_57190;
wire x_57191;
wire x_57192;
wire x_57193;
wire x_57194;
wire x_57195;
wire x_57196;
wire x_57197;
wire x_57198;
wire x_57199;
wire x_57200;
wire x_57201;
wire x_57202;
wire x_57203;
wire x_57204;
wire x_57205;
wire x_57206;
wire x_57207;
wire x_57208;
wire x_57209;
wire x_57210;
wire x_57211;
wire x_57212;
wire x_57213;
wire x_57214;
wire x_57215;
wire x_57216;
wire x_57217;
wire x_57218;
wire x_57219;
wire x_57220;
wire x_57221;
wire x_57222;
wire x_57223;
wire x_57224;
wire x_57225;
wire x_57226;
wire x_57227;
wire x_57228;
wire x_57229;
wire x_57230;
wire x_57231;
wire x_57232;
wire x_57233;
wire x_57234;
wire x_57235;
wire x_57236;
wire x_57237;
wire x_57238;
wire x_57239;
wire x_57240;
wire x_57241;
wire x_57242;
wire x_57243;
wire x_57244;
wire x_57245;
wire x_57246;
wire x_57247;
wire x_57248;
wire x_57249;
wire x_57250;
wire x_57251;
wire x_57252;
wire x_57253;
wire x_57254;
wire x_57255;
wire x_57256;
wire x_57257;
wire x_57258;
wire x_57259;
wire x_57260;
wire x_57261;
wire x_57262;
wire x_57263;
wire x_57264;
wire x_57265;
wire x_57266;
wire x_57267;
wire x_57268;
wire x_57269;
wire x_57270;
wire x_57271;
wire x_57272;
wire x_57273;
wire x_57274;
wire x_57275;
wire x_57276;
wire x_57277;
wire x_57278;
wire x_57279;
wire x_57280;
wire x_57281;
wire x_57282;
wire x_57283;
wire x_57284;
wire x_57285;
wire x_57286;
wire x_57287;
wire x_57288;
wire x_57289;
wire x_57290;
wire x_57291;
wire x_57292;
wire x_57293;
wire x_57294;
wire x_57295;
wire x_57296;
wire x_57297;
wire x_57298;
wire x_57299;
wire x_57300;
wire x_57301;
wire x_57302;
wire x_57303;
wire x_57304;
wire x_57305;
wire x_57306;
wire x_57307;
wire x_57308;
wire x_57309;
wire x_57310;
wire x_57311;
wire x_57312;
wire x_57313;
wire x_57314;
wire x_57315;
wire x_57316;
wire x_57317;
wire x_57318;
wire x_57319;
wire x_57320;
wire x_57321;
wire x_57322;
wire x_57323;
wire x_57324;
wire x_57325;
wire x_57326;
wire x_57327;
wire x_57328;
wire x_57329;
wire x_57330;
wire x_57331;
wire x_57332;
wire x_57333;
wire x_57334;
wire x_57335;
wire x_57336;
wire x_57337;
wire x_57338;
wire x_57339;
wire x_57340;
wire x_57341;
wire x_57342;
wire x_57343;
wire x_57344;
wire x_57345;
wire x_57346;
wire x_57347;
wire x_57348;
wire x_57349;
wire x_57350;
wire x_57351;
wire x_57352;
wire x_57353;
wire x_57354;
wire x_57355;
wire x_57356;
wire x_57357;
wire x_57358;
wire x_57359;
wire x_57360;
wire x_57361;
wire x_57362;
wire x_57363;
wire x_57364;
wire x_57365;
wire x_57366;
wire x_57367;
wire x_57368;
wire x_57369;
wire x_57370;
wire x_57371;
wire x_57372;
wire x_57373;
wire x_57374;
wire x_57375;
wire x_57376;
wire x_57377;
wire x_57378;
wire x_57379;
wire x_57380;
wire x_57381;
wire x_57382;
wire x_57383;
wire x_57384;
wire x_57385;
wire x_57386;
wire x_57387;
wire x_57388;
wire x_57389;
wire x_57390;
wire x_57391;
wire x_57392;
wire x_57393;
wire x_57394;
wire x_57395;
wire x_57396;
wire x_57397;
wire x_57398;
wire x_57399;
wire x_57400;
wire x_57401;
wire x_57402;
wire x_57403;
wire x_57404;
wire x_57405;
wire x_57406;
wire x_57407;
wire x_57408;
wire x_57409;
wire x_57410;
wire x_57411;
wire x_57412;
wire x_57413;
wire x_57414;
wire x_57415;
wire x_57416;
wire x_57417;
wire x_57418;
wire x_57419;
wire x_57420;
wire x_57421;
wire x_57422;
wire x_57423;
wire x_57424;
wire x_57425;
wire x_57426;
wire x_57427;
wire x_57428;
wire x_57429;
wire x_57430;
wire x_57431;
wire x_57432;
wire x_57433;
wire x_57434;
wire x_57435;
wire x_57436;
wire x_57437;
wire x_57438;
wire x_57439;
wire x_57440;
wire x_57441;
wire x_57442;
wire x_57443;
wire x_57444;
wire x_57445;
wire x_57446;
wire x_57447;
wire x_57448;
wire x_57449;
wire x_57450;
wire x_57451;
wire x_57452;
wire x_57453;
wire x_57454;
wire x_57455;
wire x_57456;
wire x_57457;
wire x_57458;
wire x_57459;
wire x_57460;
wire x_57461;
wire x_57462;
wire x_57463;
wire x_57464;
wire x_57465;
wire x_57466;
wire x_57467;
wire x_57468;
wire x_57469;
wire x_57470;
wire x_57471;
wire x_57472;
wire x_57473;
wire x_57474;
wire x_57475;
wire x_57476;
wire x_57477;
wire x_57478;
wire x_57479;
wire x_57480;
wire x_57481;
wire x_57482;
wire x_57483;
wire x_57484;
wire x_57485;
wire x_57486;
wire x_57487;
wire x_57488;
wire x_57489;
wire x_57490;
wire x_57491;
wire x_57492;
wire x_57493;
wire x_57494;
wire x_57495;
wire x_57496;
wire x_57497;
wire x_57498;
wire x_57499;
wire x_57500;
wire x_57501;
wire x_57502;
wire x_57503;
wire x_57504;
wire x_57505;
wire x_57506;
wire x_57507;
wire x_57508;
wire x_57509;
wire x_57510;
wire x_57511;
wire x_57512;
wire x_57513;
wire x_57514;
wire x_57515;
wire x_57516;
wire x_57517;
wire x_57518;
wire x_57519;
wire x_57520;
wire x_57521;
wire x_57522;
wire x_57523;
wire x_57524;
wire x_57525;
wire x_57526;
wire x_57527;
wire x_57528;
wire x_57529;
wire x_57530;
wire x_57531;
wire x_57532;
wire x_57533;
wire x_57534;
wire x_57535;
wire x_57536;
wire x_57537;
wire x_57538;
wire x_57539;
wire x_57540;
wire x_57541;
wire x_57542;
wire x_57543;
wire x_57544;
wire x_57545;
wire x_57546;
wire x_57547;
wire x_57548;
wire x_57549;
wire x_57550;
wire x_57551;
wire x_57552;
wire x_57553;
wire x_57554;
wire x_57555;
wire x_57556;
wire x_57557;
wire x_57558;
wire x_57559;
wire x_57560;
wire x_57561;
wire x_57562;
wire x_57563;
wire x_57564;
wire x_57565;
wire x_57566;
wire x_57567;
wire x_57568;
wire x_57569;
wire x_57570;
wire x_57571;
wire x_57572;
wire x_57573;
wire x_57574;
wire x_57575;
wire x_57576;
wire x_57577;
wire x_57578;
wire x_57579;
wire x_57580;
wire x_57581;
wire x_57582;
wire x_57583;
wire x_57584;
wire x_57585;
wire x_57586;
wire x_57587;
wire x_57588;
wire x_57589;
wire x_57590;
wire x_57591;
wire x_57592;
wire x_57593;
wire x_57594;
wire x_57595;
wire x_57596;
wire x_57597;
wire x_57598;
wire x_57599;
wire x_57600;
wire x_57601;
wire x_57602;
wire x_57603;
wire x_57604;
wire x_57605;
wire x_57606;
wire x_57607;
wire x_57608;
wire x_57609;
wire x_57610;
wire x_57611;
wire x_57612;
wire x_57613;
wire x_57614;
wire x_57615;
wire x_57616;
wire x_57617;
wire x_57618;
wire x_57619;
wire x_57620;
wire x_57621;
wire x_57622;
wire x_57623;
wire x_57624;
wire x_57625;
wire x_57626;
wire x_57627;
wire x_57628;
wire x_57629;
wire x_57630;
wire x_57631;
wire x_57632;
wire x_57633;
wire x_57634;
wire x_57635;
wire x_57636;
wire x_57637;
wire x_57638;
wire x_57639;
wire x_57640;
wire x_57641;
wire x_57642;
wire x_57643;
wire x_57644;
wire x_57645;
wire x_57646;
wire x_57647;
wire x_57648;
wire x_57649;
wire x_57650;
wire x_57651;
wire x_57652;
wire x_57653;
wire x_57654;
wire x_57655;
wire x_57656;
wire x_57657;
wire x_57658;
wire x_57659;
wire x_57660;
wire x_57661;
wire x_57662;
wire x_57663;
wire x_57664;
wire x_57665;
wire x_57666;
wire x_57667;
wire x_57668;
wire x_57669;
wire x_57670;
wire x_57671;
wire x_57672;
wire x_57673;
wire x_57674;
wire x_57675;
wire x_57676;
wire x_57677;
wire x_57678;
wire x_57679;
wire x_57680;
wire x_57681;
wire x_57682;
wire x_57683;
wire x_57684;
wire x_57685;
wire x_57686;
wire x_57687;
wire x_57688;
wire x_57689;
wire x_57690;
wire x_57691;
wire x_57692;
wire x_57693;
wire x_57694;
wire x_57695;
wire x_57696;
wire x_57697;
wire x_57698;
wire x_57699;
wire x_57700;
wire x_57701;
wire x_57702;
wire x_57703;
wire x_57704;
wire x_57705;
wire x_57706;
wire x_57707;
wire x_57708;
wire x_57709;
wire x_57710;
wire x_57711;
wire x_57712;
wire x_57713;
wire x_57714;
wire x_57715;
wire x_57716;
wire x_57717;
wire x_57718;
wire x_57719;
wire x_57720;
wire x_57721;
wire x_57722;
wire x_57723;
wire x_57724;
wire x_57725;
wire x_57726;
wire x_57727;
wire x_57728;
wire x_57729;
wire x_57730;
wire x_57731;
wire x_57732;
wire x_57733;
wire x_57734;
wire x_57735;
wire x_57736;
wire x_57737;
wire x_57738;
wire x_57739;
wire x_57740;
wire x_57741;
wire x_57742;
wire x_57743;
wire x_57744;
wire x_57745;
wire x_57746;
wire x_57747;
wire x_57748;
wire x_57749;
wire x_57750;
wire x_57751;
wire x_57752;
wire x_57753;
wire x_57754;
wire x_57755;
wire x_57756;
wire x_57757;
wire x_57758;
wire x_57759;
wire x_57760;
wire x_57761;
wire x_57762;
wire x_57763;
wire x_57764;
wire x_57765;
wire x_57766;
wire x_57767;
wire x_57768;
wire x_57769;
wire x_57770;
wire x_57771;
wire x_57772;
wire x_57773;
wire x_57774;
wire x_57775;
wire x_57776;
wire x_57777;
wire x_57778;
wire x_57779;
wire x_57780;
wire x_57781;
wire x_57782;
wire x_57783;
wire x_57784;
wire x_57785;
wire x_57786;
wire x_57787;
wire x_57788;
wire x_57789;
wire x_57790;
wire x_57791;
wire x_57792;
wire x_57793;
wire x_57794;
wire x_57795;
wire x_57796;
wire x_57797;
wire x_57798;
wire x_57799;
wire x_57800;
wire x_57801;
wire x_57802;
wire x_57803;
wire x_57804;
wire x_57805;
wire x_57806;
wire x_57807;
wire x_57808;
wire x_57809;
wire x_57810;
wire x_57811;
wire x_57812;
wire x_57813;
wire x_57814;
wire x_57815;
wire x_57816;
wire x_57817;
wire x_57818;
wire x_57819;
wire x_57820;
wire x_57821;
wire x_57822;
wire x_57823;
wire x_57824;
wire x_57825;
wire x_57826;
wire x_57827;
wire x_57828;
wire x_57829;
wire x_57830;
wire x_57831;
wire x_57832;
wire x_57833;
wire x_57834;
wire x_57835;
wire x_57836;
wire x_57837;
wire x_57838;
wire x_57839;
wire x_57840;
wire x_57841;
wire x_57842;
wire x_57843;
wire x_57844;
wire x_57845;
wire x_57846;
wire x_57847;
wire x_57848;
wire x_57849;
wire x_57850;
wire x_57851;
wire x_57852;
wire x_57853;
wire x_57854;
wire x_57855;
wire x_57856;
wire x_57857;
wire x_57858;
wire x_57859;
wire x_57860;
wire x_57861;
wire x_57862;
wire x_57863;
wire x_57864;
wire x_57865;
wire x_57866;
wire x_57867;
wire x_57868;
wire x_57869;
wire x_57870;
wire x_57871;
wire x_57872;
wire x_57873;
wire x_57874;
wire x_57875;
wire x_57876;
wire x_57877;
wire x_57878;
wire x_57879;
wire x_57880;
wire x_57881;
wire x_57882;
wire x_57883;
wire x_57884;
wire x_57885;
wire x_57886;
wire x_57887;
wire x_57888;
wire x_57889;
wire x_57890;
wire x_57891;
wire x_57892;
wire x_57893;
wire x_57894;
wire x_57895;
wire x_57896;
wire x_57897;
wire x_57898;
wire x_57899;
wire x_57900;
wire x_57901;
wire x_57902;
wire x_57903;
wire x_57904;
wire x_57905;
wire x_57906;
wire x_57907;
wire x_57908;
wire x_57909;
wire x_57910;
wire x_57911;
wire x_57912;
wire x_57913;
wire x_57914;
wire x_57915;
wire x_57916;
wire x_57917;
wire x_57918;
wire x_57919;
wire x_57920;
wire x_57921;
wire x_57922;
wire x_57923;
wire x_57924;
wire x_57925;
wire x_57926;
wire x_57927;
wire x_57928;
wire x_57929;
wire x_57930;
wire x_57931;
wire x_57932;
wire x_57933;
wire x_57934;
wire x_57935;
wire x_57936;
wire x_57937;
wire x_57938;
wire x_57939;
wire x_57940;
wire x_57941;
wire x_57942;
wire x_57943;
wire x_57944;
wire x_57945;
wire x_57946;
wire x_57947;
wire x_57948;
wire x_57949;
wire x_57950;
wire x_57951;
wire x_57952;
wire x_57953;
wire x_57954;
wire x_57955;
wire x_57956;
wire x_57957;
wire x_57958;
wire x_57959;
wire x_57960;
wire x_57961;
wire x_57962;
wire x_57963;
wire x_57964;
wire x_57965;
wire x_57966;
wire x_57967;
wire x_57968;
wire x_57969;
wire x_57970;
wire x_57971;
wire x_57972;
wire x_57973;
wire x_57974;
wire x_57975;
wire x_57976;
wire x_57977;
wire x_57978;
wire x_57979;
wire x_57980;
wire x_57981;
wire x_57982;
wire x_57983;
wire x_57984;
wire x_57985;
wire x_57986;
wire x_57987;
wire x_57988;
wire x_57989;
wire x_57990;
wire x_57991;
wire x_57992;
wire x_57993;
wire x_57994;
wire x_57995;
wire x_57996;
wire x_57997;
wire x_57998;
wire x_57999;
wire x_58000;
wire x_58001;
wire x_58002;
wire x_58003;
wire x_58004;
wire x_58005;
wire x_58006;
wire x_58007;
wire x_58008;
wire x_58009;
wire x_58010;
wire x_58011;
wire x_58012;
wire x_58013;
wire x_58014;
wire x_58015;
wire x_58016;
wire x_58017;
wire x_58018;
wire x_58019;
wire x_58020;
wire x_58021;
wire x_58022;
wire x_58023;
wire x_58024;
wire x_58025;
wire x_58026;
wire x_58027;
wire x_58028;
wire x_58029;
wire x_58030;
wire x_58031;
wire x_58032;
wire x_58033;
wire x_58034;
wire x_58035;
wire x_58036;
wire x_58037;
wire x_58038;
wire x_58039;
wire x_58040;
wire x_58041;
wire x_58042;
wire x_58043;
wire x_58044;
wire x_58045;
wire x_58046;
wire x_58047;
wire x_58048;
wire x_58049;
wire x_58050;
wire x_58051;
wire x_58052;
wire x_58053;
wire x_58054;
wire x_58055;
wire x_58056;
wire x_58057;
wire x_58058;
wire x_58059;
wire x_58060;
wire x_58061;
wire x_58062;
wire x_58063;
wire x_58064;
wire x_58065;
wire x_58066;
wire x_58067;
wire x_58068;
wire x_58069;
wire x_58070;
wire x_58071;
wire x_58072;
wire x_58073;
wire x_58074;
wire x_58075;
wire x_58076;
wire x_58077;
wire x_58078;
wire x_58079;
wire x_58080;
wire x_58081;
wire x_58082;
wire x_58083;
wire x_58084;
wire x_58085;
wire x_58086;
wire x_58087;
wire x_58088;
wire x_58089;
wire x_58090;
wire x_58091;
wire x_58092;
wire x_58093;
wire x_58094;
wire x_58095;
wire x_58096;
wire x_58097;
wire x_58098;
wire x_58099;
wire x_58100;
wire x_58101;
wire x_58102;
wire x_58103;
wire x_58104;
wire x_58105;
wire x_58106;
wire x_58107;
wire x_58108;
wire x_58109;
wire x_58110;
wire x_58111;
wire x_58112;
wire x_58113;
wire x_58114;
wire x_58115;
wire x_58116;
wire x_58117;
wire x_58118;
wire x_58119;
wire x_58120;
wire x_58121;
wire x_58122;
wire x_58123;
wire x_58124;
wire x_58125;
wire x_58126;
wire x_58127;
wire x_58128;
wire x_58129;
wire x_58130;
wire x_58131;
wire x_58132;
wire x_58133;
wire x_58134;
wire x_58135;
wire x_58136;
wire x_58137;
wire x_58138;
wire x_58139;
wire x_58140;
wire x_58141;
wire x_58142;
wire x_58143;
wire x_58144;
wire x_58145;
wire x_58146;
wire x_58147;
wire x_58148;
wire x_58149;
wire x_58150;
wire x_58151;
wire x_58152;
wire x_58153;
wire x_58154;
wire x_58155;
wire x_58156;
wire x_58157;
wire x_58158;
wire x_58159;
wire x_58160;
wire x_58161;
wire x_58162;
wire x_58163;
wire x_58164;
wire x_58165;
wire x_58166;
wire x_58167;
wire x_58168;
wire x_58169;
wire x_58170;
wire x_58171;
wire x_58172;
wire x_58173;
wire x_58174;
wire x_58175;
wire x_58176;
wire x_58177;
wire x_58178;
wire x_58179;
wire x_58180;
wire x_58181;
wire x_58182;
wire x_58183;
wire x_58184;
wire x_58185;
wire x_58186;
wire x_58187;
wire x_58188;
wire x_58189;
wire x_58190;
wire x_58191;
wire x_58192;
wire x_58193;
wire x_58194;
wire x_58195;
wire x_58196;
wire x_58197;
wire x_58198;
wire x_58199;
wire x_58200;
wire x_58201;
wire x_58202;
wire x_58203;
wire x_58204;
wire x_58205;
wire x_58206;
wire x_58207;
wire x_58208;
wire x_58209;
wire x_58210;
wire x_58211;
wire x_58212;
wire x_58213;
wire x_58214;
wire x_58215;
wire x_58216;
wire x_58217;
wire x_58218;
wire x_58219;
wire x_58220;
wire x_58221;
wire x_58222;
wire x_58223;
wire x_58224;
wire x_58225;
wire x_58226;
wire x_58227;
wire x_58228;
wire x_58229;
wire x_58230;
wire x_58231;
wire x_58232;
wire x_58233;
wire x_58234;
wire x_58235;
wire x_58236;
wire x_58237;
wire x_58238;
wire x_58239;
wire x_58240;
wire x_58241;
wire x_58242;
wire x_58243;
wire x_58244;
wire x_58245;
wire x_58246;
wire x_58247;
wire x_58248;
wire x_58249;
wire x_58250;
wire x_58251;
wire x_58252;
wire x_58253;
wire x_58254;
wire x_58255;
wire x_58256;
wire x_58257;
wire x_58258;
wire x_58259;
wire x_58260;
wire x_58261;
wire x_58262;
wire x_58263;
wire x_58264;
wire x_58265;
wire x_58266;
wire x_58267;
wire x_58268;
wire x_58269;
wire x_58270;
wire x_58271;
wire x_58272;
wire x_58273;
wire x_58274;
wire x_58275;
wire x_58276;
wire x_58277;
wire x_58278;
wire x_58279;
wire x_58280;
wire x_58281;
wire x_58282;
wire x_58283;
wire x_58284;
wire x_58285;
wire x_58286;
wire x_58287;
wire x_58288;
wire x_58289;
wire x_58290;
wire x_58291;
wire x_58292;
wire x_58293;
wire x_58294;
wire x_58295;
wire x_58296;
wire x_58297;
wire x_58298;
wire x_58299;
wire x_58300;
wire x_58301;
wire x_58302;
wire x_58303;
wire x_58304;
wire x_58305;
wire x_58306;
wire x_58307;
wire x_58308;
wire x_58309;
wire x_58310;
wire x_58311;
wire x_58312;
wire x_58313;
wire x_58314;
wire x_58315;
wire x_58316;
wire x_58317;
wire x_58318;
wire x_58319;
wire x_58320;
wire x_58321;
wire x_58322;
wire x_58323;
wire x_58324;
wire x_58325;
wire x_58326;
wire x_58327;
wire x_58328;
wire x_58329;
wire x_58330;
wire x_58331;
wire x_58332;
wire x_58333;
wire x_58334;
wire x_58335;
wire x_58336;
wire x_58337;
wire x_58338;
wire x_58339;
wire x_58340;
wire x_58341;
wire x_58342;
wire x_58343;
wire x_58344;
wire x_58345;
wire x_58346;
wire x_58347;
wire x_58348;
wire x_58349;
wire x_58350;
wire x_58351;
wire x_58352;
wire x_58353;
wire x_58354;
wire x_58355;
wire x_58356;
wire x_58357;
wire x_58358;
wire x_58359;
wire x_58360;
wire x_58361;
wire x_58362;
wire x_58363;
wire x_58364;
wire x_58365;
wire x_58366;
wire x_58367;
wire x_58368;
wire x_58369;
wire x_58370;
wire x_58371;
wire x_58372;
wire x_58373;
wire x_58374;
wire x_58375;
wire x_58376;
wire x_58377;
wire x_58378;
wire x_58379;
wire x_58380;
wire x_58381;
wire x_58382;
wire x_58383;
wire x_58384;
wire x_58385;
wire x_58386;
wire x_58387;
wire x_58388;
wire x_58389;
wire x_58390;
wire x_58391;
wire x_58392;
wire x_58393;
wire x_58394;
wire x_58395;
wire x_58396;
wire x_58397;
wire x_58398;
wire x_58399;
wire x_58400;
wire x_58401;
wire x_58402;
wire x_58403;
wire x_58404;
wire x_58405;
wire x_58406;
wire x_58407;
wire x_58408;
wire x_58409;
wire x_58410;
wire x_58411;
wire x_58412;
wire x_58413;
wire x_58414;
wire x_58415;
wire x_58416;
wire x_58417;
wire x_58418;
wire x_58419;
wire x_58420;
wire x_58421;
wire x_58422;
wire x_58423;
wire x_58424;
wire x_58425;
wire x_58426;
wire x_58427;
wire x_58428;
wire x_58429;
wire x_58430;
wire x_58431;
wire x_58432;
wire x_58433;
wire x_58434;
wire x_58435;
wire x_58436;
wire x_58437;
wire x_58438;
wire x_58439;
wire x_58440;
wire x_58441;
wire x_58442;
wire x_58443;
wire x_58444;
wire x_58445;
wire x_58446;
wire x_58447;
wire x_58448;
wire x_58449;
wire x_58450;
wire x_58451;
wire x_58452;
wire x_58453;
wire x_58454;
wire x_58455;
wire x_58456;
wire x_58457;
wire x_58458;
wire x_58459;
wire x_58460;
wire x_58461;
wire x_58462;
wire x_58463;
wire x_58464;
wire x_58465;
wire x_58466;
wire x_58467;
wire x_58468;
wire x_58469;
wire x_58470;
wire x_58471;
wire x_58472;
wire x_58473;
wire x_58474;
wire x_58475;
wire x_58476;
wire x_58477;
wire x_58478;
wire x_58479;
wire x_58480;
wire x_58481;
wire x_58482;
wire x_58483;
wire x_58484;
wire x_58485;
wire x_58486;
wire x_58487;
wire x_58488;
wire x_58489;
wire x_58490;
wire x_58491;
wire x_58492;
wire x_58493;
wire x_58494;
wire x_58495;
wire x_58496;
wire x_58497;
wire x_58498;
wire x_58499;
wire x_58500;
wire x_58501;
wire x_58502;
wire x_58503;
wire x_58504;
wire x_58505;
wire x_58506;
wire x_58507;
wire x_58508;
wire x_58509;
wire x_58510;
wire x_58511;
wire x_58512;
wire x_58513;
wire x_58514;
wire x_58515;
wire x_58516;
wire x_58517;
wire x_58518;
wire x_58519;
wire x_58520;
wire x_58521;
wire x_58522;
wire x_58523;
wire x_58524;
wire x_58525;
wire x_58526;
wire x_58527;
wire x_58528;
wire x_58529;
wire x_58530;
wire x_58531;
wire x_58532;
wire x_58533;
wire x_58534;
wire x_58535;
wire x_58536;
wire x_58537;
wire x_58538;
wire x_58539;
wire x_58540;
wire x_58541;
wire x_58542;
wire x_58543;
wire x_58544;
wire x_58545;
wire x_58546;
wire x_58547;
wire x_58548;
wire x_58549;
wire x_58550;
wire x_58551;
wire x_58552;
wire x_58553;
wire x_58554;
wire x_58555;
wire x_58556;
wire x_58557;
wire x_58558;
wire x_58559;
wire x_58560;
wire x_58561;
wire x_58562;
wire x_58563;
wire x_58564;
wire x_58565;
wire x_58566;
wire x_58567;
wire x_58568;
wire x_58569;
wire x_58570;
wire x_58571;
wire x_58572;
wire x_58573;
wire x_58574;
wire x_58575;
wire x_58576;
wire x_58577;
wire x_58578;
wire x_58579;
wire x_58580;
wire x_58581;
wire x_58582;
wire x_58583;
wire x_58584;
wire x_58585;
wire x_58586;
wire x_58587;
wire x_58588;
wire x_58589;
wire x_58590;
wire x_58591;
wire x_58592;
wire x_58593;
wire x_58594;
wire x_58595;
wire x_58596;
wire x_58597;
wire x_58598;
wire x_58599;
wire x_58600;
wire x_58601;
wire x_58602;
wire x_58603;
wire x_58604;
wire x_58605;
wire x_58606;
wire x_58607;
wire x_58608;
wire x_58609;
wire x_58610;
wire x_58611;
wire x_58612;
wire x_58613;
wire x_58614;
wire x_58615;
wire x_58616;
wire x_58617;
wire x_58618;
wire x_58619;
wire x_58620;
wire x_58621;
wire x_58622;
wire x_58623;
wire x_58624;
wire x_58625;
wire x_58626;
wire x_58627;
wire x_58628;
wire x_58629;
wire x_58630;
wire x_58631;
wire x_58632;
wire x_58633;
wire x_58634;
wire x_58635;
wire x_58636;
wire x_58637;
wire x_58638;
wire x_58639;
wire x_58640;
wire x_58641;
wire x_58642;
wire x_58643;
wire x_58644;
wire x_58645;
wire x_58646;
wire x_58647;
wire x_58648;
wire x_58649;
wire x_58650;
wire x_58651;
wire x_58652;
wire x_58653;
wire x_58654;
wire x_58655;
wire x_58656;
wire x_58657;
wire x_58658;
wire x_58659;
wire x_58660;
wire x_58661;
wire x_58662;
wire x_58663;
wire x_58664;
wire x_58665;
wire x_58666;
wire x_58667;
wire x_58668;
wire x_58669;
wire x_58670;
wire x_58671;
wire x_58672;
wire x_58673;
wire x_58674;
wire x_58675;
wire x_58676;
wire x_58677;
wire x_58678;
wire x_58679;
wire x_58680;
wire x_58681;
wire x_58682;
wire x_58683;
wire x_58684;
wire x_58685;
wire x_58686;
wire x_58687;
wire x_58688;
wire x_58689;
wire x_58690;
wire x_58691;
wire x_58692;
wire x_58693;
wire x_58694;
wire x_58695;
wire x_58696;
wire x_58697;
wire x_58698;
wire x_58699;
wire x_58700;
wire x_58701;
wire x_58702;
wire x_58703;
wire x_58704;
wire x_58705;
wire x_58706;
wire x_58707;
wire x_58708;
wire x_58709;
wire x_58710;
wire x_58711;
wire x_58712;
wire x_58713;
wire x_58714;
wire x_58715;
wire x_58716;
wire x_58717;
wire x_58718;
wire x_58719;
wire x_58720;
wire x_58721;
wire x_58722;
wire x_58723;
wire x_58724;
wire x_58725;
wire x_58726;
wire x_58727;
wire x_58728;
wire x_58729;
wire x_58730;
wire x_58731;
wire x_58732;
wire x_58733;
wire x_58734;
wire x_58735;
wire x_58736;
wire x_58737;
wire x_58738;
wire x_58739;
wire x_58740;
wire x_58741;
wire x_58742;
wire x_58743;
wire x_58744;
wire x_58745;
wire x_58746;
wire x_58747;
wire x_58748;
wire x_58749;
wire x_58750;
wire x_58751;
wire x_58752;
wire x_58753;
wire x_58754;
wire x_58755;
wire x_58756;
wire x_58757;
wire x_58758;
wire x_58759;
wire x_58760;
wire x_58761;
wire x_58762;
wire x_58763;
wire x_58764;
wire x_58765;
wire x_58766;
wire x_58767;
wire x_58768;
wire x_58769;
wire x_58770;
wire x_58771;
wire x_58772;
wire x_58773;
wire x_58774;
wire x_58775;
wire x_58776;
wire x_58777;
wire x_58778;
wire x_58779;
wire x_58780;
wire x_58781;
wire x_58782;
wire x_58783;
wire x_58784;
wire x_58785;
wire x_58786;
wire x_58787;
wire x_58788;
wire x_58789;
wire x_58790;
wire x_58791;
wire x_58792;
wire x_58793;
wire x_58794;
wire x_58795;
wire x_58796;
wire x_58797;
wire x_58798;
wire x_58799;
wire x_58800;
wire x_58801;
wire x_58802;
wire x_58803;
wire x_58804;
wire x_58805;
wire x_58806;
wire x_58807;
wire x_58808;
wire x_58809;
wire x_58810;
wire x_58811;
wire x_58812;
wire x_58813;
wire x_58814;
wire x_58815;
wire x_58816;
wire x_58817;
wire x_58818;
wire x_58819;
wire x_58820;
wire x_58821;
wire x_58822;
wire x_58823;
wire x_58824;
wire x_58825;
wire x_58826;
wire x_58827;
wire x_58828;
wire x_58829;
wire x_58830;
wire x_58831;
wire x_58832;
wire x_58833;
wire x_58834;
wire x_58835;
wire x_58836;
wire x_58837;
wire x_58838;
wire x_58839;
wire x_58840;
wire x_58841;
wire x_58842;
wire x_58843;
wire x_58844;
wire x_58845;
wire x_58846;
wire x_58847;
wire x_58848;
wire x_58849;
wire x_58850;
wire x_58851;
wire x_58852;
wire x_58853;
wire x_58854;
wire x_58855;
wire x_58856;
wire x_58857;
wire x_58858;
wire x_58859;
wire x_58860;
wire x_58861;
wire x_58862;
wire x_58863;
wire x_58864;
wire x_58865;
wire x_58866;
wire x_58867;
wire x_58868;
wire x_58869;
wire x_58870;
wire x_58871;
wire x_58872;
wire x_58873;
wire x_58874;
wire x_58875;
wire x_58876;
wire x_58877;
wire x_58878;
wire x_58879;
wire x_58880;
wire x_58881;
wire x_58882;
wire x_58883;
wire x_58884;
wire x_58885;
wire x_58886;
wire x_58887;
wire x_58888;
wire x_58889;
wire x_58890;
wire x_58891;
wire x_58892;
wire x_58893;
wire x_58894;
wire x_58895;
wire x_58896;
wire x_58897;
wire x_58898;
wire x_58899;
wire x_58900;
wire x_58901;
wire x_58902;
wire x_58903;
wire x_58904;
wire x_58905;
wire x_58906;
wire x_58907;
wire x_58908;
wire x_58909;
wire x_58910;
wire x_58911;
wire x_58912;
wire x_58913;
wire x_58914;
wire x_58915;
wire x_58916;
wire x_58917;
wire x_58918;
wire x_58919;
wire x_58920;
wire x_58921;
wire x_58922;
wire x_58923;
wire x_58924;
wire x_58925;
wire x_58926;
wire x_58927;
wire x_58928;
wire x_58929;
wire x_58930;
wire x_58931;
wire x_58932;
wire x_58933;
wire x_58934;
wire x_58935;
wire x_58936;
wire x_58937;
wire x_58938;
wire x_58939;
wire x_58940;
wire x_58941;
wire x_58942;
wire x_58943;
wire x_58944;
wire x_58945;
wire x_58946;
wire x_58947;
wire x_58948;
wire x_58949;
wire x_58950;
wire x_58951;
wire x_58952;
wire x_58953;
wire x_58954;
wire x_58955;
wire x_58956;
wire x_58957;
wire x_58958;
wire x_58959;
wire x_58960;
wire x_58961;
wire x_58962;
wire x_58963;
wire x_58964;
wire x_58965;
wire x_58966;
wire x_58967;
wire x_58968;
wire x_58969;
wire x_58970;
wire x_58971;
wire x_58972;
wire x_58973;
wire x_58974;
wire x_58975;
wire x_58976;
wire x_58977;
wire x_58978;
wire x_58979;
wire x_58980;
wire x_58981;
wire x_58982;
wire x_58983;
wire x_58984;
wire x_58985;
wire x_58986;
wire x_58987;
wire x_58988;
wire x_58989;
wire x_58990;
wire x_58991;
wire x_58992;
wire x_58993;
wire x_58994;
wire x_58995;
wire x_58996;
wire x_58997;
wire x_58998;
wire x_58999;
wire x_59000;
wire x_59001;
wire x_59002;
wire x_59003;
wire x_59004;
wire x_59005;
wire x_59006;
wire x_59007;
wire x_59008;
wire x_59009;
wire x_59010;
wire x_59011;
wire x_59012;
wire x_59013;
wire x_59014;
wire x_59015;
wire x_59016;
wire x_59017;
wire x_59018;
wire x_59019;
wire x_59020;
wire x_59021;
wire x_59022;
wire x_59023;
wire x_59024;
wire x_59025;
wire x_59026;
wire x_59027;
wire x_59028;
wire x_59029;
wire x_59030;
wire x_59031;
wire x_59032;
wire x_59033;
wire x_59034;
wire x_59035;
wire x_59036;
wire x_59037;
wire x_59038;
wire x_59039;
wire x_59040;
wire x_59041;
wire x_59042;
wire x_59043;
wire x_59044;
wire x_59045;
wire x_59046;
wire x_59047;
wire x_59048;
wire x_59049;
wire x_59050;
wire x_59051;
wire x_59052;
wire x_59053;
wire x_59054;
wire x_59055;
wire x_59056;
wire x_59057;
wire x_59058;
wire x_59059;
wire x_59060;
wire x_59061;
wire x_59062;
wire x_59063;
wire x_59064;
wire x_59065;
wire x_59066;
wire x_59067;
wire x_59068;
wire x_59069;
wire x_59070;
wire x_59071;
wire x_59072;
wire x_59073;
wire x_59074;
wire x_59075;
wire x_59076;
wire x_59077;
wire x_59078;
wire x_59079;
wire x_59080;
wire x_59081;
wire x_59082;
wire x_59083;
wire x_59084;
wire x_59085;
wire x_59086;
wire x_59087;
wire x_59088;
wire x_59089;
wire x_59090;
wire x_59091;
wire x_59092;
wire x_59093;
wire x_59094;
wire x_59095;
wire x_59096;
wire x_59097;
wire x_59098;
wire x_59099;
wire x_59100;
wire x_59101;
wire x_59102;
wire x_59103;
wire x_59104;
wire x_59105;
wire x_59106;
wire x_59107;
wire x_59108;
wire x_59109;
wire x_59110;
wire x_59111;
wire x_59112;
wire x_59113;
wire x_59114;
wire x_59115;
wire x_59116;
wire x_59117;
wire x_59118;
wire x_59119;
wire x_59120;
wire x_59121;
wire x_59122;
wire x_59123;
wire x_59124;
wire x_59125;
wire x_59126;
wire x_59127;
wire x_59128;
wire x_59129;
wire x_59130;
wire x_59131;
wire x_59132;
wire x_59133;
wire x_59134;
wire x_59135;
wire x_59136;
wire x_59137;
wire x_59138;
wire x_59139;
wire x_59140;
wire x_59141;
wire x_59142;
wire x_59143;
wire x_59144;
wire x_59145;
wire x_59146;
wire x_59147;
wire x_59148;
wire x_59149;
wire x_59150;
wire x_59151;
wire x_59152;
wire x_59153;
wire x_59154;
wire x_59155;
wire x_59156;
wire x_59157;
wire x_59158;
wire x_59159;
wire x_59160;
wire x_59161;
wire x_59162;
wire x_59163;
wire x_59164;
wire x_59165;
wire x_59166;
wire x_59167;
wire x_59168;
wire x_59169;
wire x_59170;
wire x_59171;
wire x_59172;
wire x_59173;
wire x_59174;
wire x_59175;
wire x_59176;
wire x_59177;
wire x_59178;
wire x_59179;
wire x_59180;
wire x_59181;
wire x_59182;
wire x_59183;
wire x_59184;
wire x_59185;
wire x_59186;
wire x_59187;
wire x_59188;
wire x_59189;
wire x_59190;
wire x_59191;
wire x_59192;
wire x_59193;
wire x_59194;
wire x_59195;
wire x_59196;
wire x_59197;
wire x_59198;
wire x_59199;
wire x_59200;
wire x_59201;
wire x_59202;
wire x_59203;
wire x_59204;
wire x_59205;
wire x_59206;
wire x_59207;
wire x_59208;
wire x_59209;
wire x_59210;
wire x_59211;
wire x_59212;
wire x_59213;
wire x_59214;
wire x_59215;
wire x_59216;
wire x_59217;
wire x_59218;
wire x_59219;
wire x_59220;
wire x_59221;
wire x_59222;
wire x_59223;
wire x_59224;
wire x_59225;
wire x_59226;
wire x_59227;
wire x_59228;
wire x_59229;
wire x_59230;
wire x_59231;
wire x_59232;
wire x_59233;
wire x_59234;
wire x_59235;
wire x_59236;
wire x_59237;
wire x_59238;
wire x_59239;
wire x_59240;
wire x_59241;
wire x_59242;
wire x_59243;
wire x_59244;
wire x_59245;
wire x_59246;
wire x_59247;
wire x_59248;
wire x_59249;
wire x_59250;
wire x_59251;
wire x_59252;
wire x_59253;
wire x_59254;
wire x_59255;
wire x_59256;
wire x_59257;
wire x_59258;
wire x_59259;
wire x_59260;
wire x_59261;
wire x_59262;
wire x_59263;
wire x_59264;
wire x_59265;
wire x_59266;
wire x_59267;
wire x_59268;
wire x_59269;
wire x_59270;
wire x_59271;
wire x_59272;
wire x_59273;
wire x_59274;
wire x_59275;
wire x_59276;
wire x_59277;
wire x_59278;
wire x_59279;
wire x_59280;
wire x_59281;
wire x_59282;
wire x_59283;
wire x_59284;
wire x_59285;
wire x_59286;
wire x_59287;
wire x_59288;
wire x_59289;
wire x_59290;
wire x_59291;
wire x_59292;
wire x_59293;
wire x_59294;
wire x_59295;
wire x_59296;
wire x_59297;
wire x_59298;
wire x_59299;
wire x_59300;
wire x_59301;
wire x_59302;
wire x_59303;
wire x_59304;
wire x_59305;
wire x_59306;
wire x_59307;
wire x_59308;
wire x_59309;
wire x_59310;
wire x_59311;
wire x_59312;
wire x_59313;
wire x_59314;
wire x_59315;
wire x_59316;
wire x_59317;
wire x_59318;
wire x_59319;
wire x_59320;
wire x_59321;
wire x_59322;
wire x_59323;
wire x_59324;
wire x_59325;
wire x_59326;
wire x_59327;
wire x_59328;
wire x_59329;
wire x_59330;
wire x_59331;
wire x_59332;
wire x_59333;
wire x_59334;
wire x_59335;
wire x_59336;
wire x_59337;
wire x_59338;
wire x_59339;
wire x_59340;
wire x_59341;
wire x_59342;
wire x_59343;
wire x_59344;
wire x_59345;
wire x_59346;
wire x_59347;
wire x_59348;
wire x_59349;
wire x_59350;
wire x_59351;
wire x_59352;
wire x_59353;
wire x_59354;
wire x_59355;
wire x_59356;
wire x_59357;
wire x_59358;
wire x_59359;
wire x_59360;
wire x_59361;
wire x_59362;
wire x_59363;
wire x_59364;
wire x_59365;
wire x_59366;
wire x_59367;
wire x_59368;
wire x_59369;
wire x_59370;
wire x_59371;
wire x_59372;
wire x_59373;
wire x_59374;
wire x_59375;
wire x_59376;
wire x_59377;
wire x_59378;
wire x_59379;
wire x_59380;
wire x_59381;
wire x_59382;
wire x_59383;
wire x_59384;
wire x_59385;
wire x_59386;
wire x_59387;
wire x_59388;
wire x_59389;
wire x_59390;
wire x_59391;
wire x_59392;
wire x_59393;
wire x_59394;
wire x_59395;
wire x_59396;
wire x_59397;
wire x_59398;
wire x_59399;
wire x_59400;
wire x_59401;
wire x_59402;
wire x_59403;
wire x_59404;
wire x_59405;
wire x_59406;
wire x_59407;
wire x_59408;
wire x_59409;
wire x_59410;
wire x_59411;
wire x_59412;
wire x_59413;
wire x_59414;
wire x_59415;
wire x_59416;
wire x_59417;
wire x_59418;
wire x_59419;
wire x_59420;
wire x_59421;
wire x_59422;
wire x_59423;
wire x_59424;
wire x_59425;
wire x_59426;
wire x_59427;
wire x_59428;
wire x_59429;
wire x_59430;
wire x_59431;
wire x_59432;
wire x_59433;
wire x_59434;
wire x_59435;
wire x_59436;
wire x_59437;
wire x_59438;
wire x_59439;
wire x_59440;
wire x_59441;
wire x_59442;
wire x_59443;
wire x_59444;
wire x_59445;
wire x_59446;
wire x_59447;
wire x_59448;
wire x_59449;
wire x_59450;
wire x_59451;
wire x_59452;
wire x_59453;
wire x_59454;
wire x_59455;
wire x_59456;
wire x_59457;
wire x_59458;
wire x_59459;
wire x_59460;
wire x_59461;
wire x_59462;
wire x_59463;
wire x_59464;
wire x_59465;
wire x_59466;
wire x_59467;
wire x_59468;
wire x_59469;
wire x_59470;
wire x_59471;
wire x_59472;
wire x_59473;
wire x_59474;
wire x_59475;
wire x_59476;
wire x_59477;
wire x_59478;
wire x_59479;
wire x_59480;
wire x_59481;
wire x_59482;
wire x_59483;
wire x_59484;
wire x_59485;
wire x_59486;
wire x_59487;
wire x_59488;
wire x_59489;
wire x_59490;
wire x_59491;
wire x_59492;
wire x_59493;
wire x_59494;
wire x_59495;
wire x_59496;
wire x_59497;
wire x_59498;
wire x_59499;
wire x_59500;
wire x_59501;
wire x_59502;
wire x_59503;
wire x_59504;
wire x_59505;
wire x_59506;
wire x_59507;
wire x_59508;
wire x_59509;
wire x_59510;
wire x_59511;
wire x_59512;
wire x_59513;
wire x_59514;
wire x_59515;
wire x_59516;
wire x_59517;
wire x_59518;
wire x_59519;
wire x_59520;
wire x_59521;
wire x_59522;
wire x_59523;
wire x_59524;
wire x_59525;
wire x_59526;
wire x_59527;
wire x_59528;
wire x_59529;
wire x_59530;
wire x_59531;
wire x_59532;
wire x_59533;
wire x_59534;
wire x_59535;
wire x_59536;
wire x_59537;
wire x_59538;
wire x_59539;
wire x_59540;
wire x_59541;
wire x_59542;
wire x_59543;
wire x_59544;
wire x_59545;
wire x_59546;
wire x_59547;
wire x_59548;
wire x_59549;
wire x_59550;
wire x_59551;
wire x_59552;
wire x_59553;
wire x_59554;
wire x_59555;
wire x_59556;
wire x_59557;
wire x_59558;
wire x_59559;
wire x_59560;
wire x_59561;
wire x_59562;
wire x_59563;
wire x_59564;
wire x_59565;
wire x_59566;
wire x_59567;
wire x_59568;
wire x_59569;
wire x_59570;
wire x_59571;
wire x_59572;
wire x_59573;
wire x_59574;
wire x_59575;
wire x_59576;
wire x_59577;
wire x_59578;
wire x_59579;
wire x_59580;
wire x_59581;
wire x_59582;
wire x_59583;
wire x_59584;
wire x_59585;
wire x_59586;
wire x_59587;
wire x_59588;
wire x_59589;
wire x_59590;
wire x_59591;
wire x_59592;
wire x_59593;
wire x_59594;
wire x_59595;
wire x_59596;
wire x_59597;
wire x_59598;
wire x_59599;
wire x_59600;
wire x_59601;
wire x_59602;
wire x_59603;
wire x_59604;
wire x_59605;
wire x_59606;
wire x_59607;
wire x_59608;
wire x_59609;
wire x_59610;
wire x_59611;
wire x_59612;
wire x_59613;
wire x_59614;
wire x_59615;
wire x_59616;
wire x_59617;
wire x_59618;
wire x_59619;
wire x_59620;
wire x_59621;
wire x_59622;
wire x_59623;
wire x_59624;
wire x_59625;
wire x_59626;
wire x_59627;
wire x_59628;
wire x_59629;
wire x_59630;
wire x_59631;
wire x_59632;
wire x_59633;
wire x_59634;
wire x_59635;
wire x_59636;
wire x_59637;
wire x_59638;
wire x_59639;
wire x_59640;
wire x_59641;
wire x_59642;
wire x_59643;
wire x_59644;
wire x_59645;
wire x_59646;
wire x_59647;
wire x_59648;
wire x_59649;
wire x_59650;
wire x_59651;
wire x_59652;
wire x_59653;
wire x_59654;
wire x_59655;
wire x_59656;
wire x_59657;
wire x_59658;
wire x_59659;
wire x_59660;
wire x_59661;
wire x_59662;
wire x_59663;
wire x_59664;
wire x_59665;
wire x_59666;
wire x_59667;
wire x_59668;
wire x_59669;
wire x_59670;
wire x_59671;
wire x_59672;
wire x_59673;
wire x_59674;
wire x_59675;
wire x_59676;
wire x_59677;
wire x_59678;
wire x_59679;
wire x_59680;
wire x_59681;
wire x_59682;
wire x_59683;
wire x_59684;
wire x_59685;
wire x_59686;
wire x_59687;
wire x_59688;
wire x_59689;
wire x_59690;
wire x_59691;
wire x_59692;
wire x_59693;
wire x_59694;
wire x_59695;
wire x_59696;
wire x_59697;
wire x_59698;
wire x_59699;
wire x_59700;
wire x_59701;
wire x_59702;
wire x_59703;
wire x_59704;
wire x_59705;
wire x_59706;
wire x_59707;
wire x_59708;
wire x_59709;
wire x_59710;
wire x_59711;
wire x_59712;
wire x_59713;
wire x_59714;
wire x_59715;
wire x_59716;
wire x_59717;
wire x_59718;
wire x_59719;
wire x_59720;
wire x_59721;
wire x_59722;
wire x_59723;
wire x_59724;
wire x_59725;
wire x_59726;
wire x_59727;
wire x_59728;
wire x_59729;
wire x_59730;
wire x_59731;
wire x_59732;
wire x_59733;
wire x_59734;
wire x_59735;
wire x_59736;
wire x_59737;
wire x_59738;
wire x_59739;
wire x_59740;
wire x_59741;
wire x_59742;
wire x_59743;
wire x_59744;
wire x_59745;
wire x_59746;
wire x_59747;
wire x_59748;
wire x_59749;
wire x_59750;
wire x_59751;
wire x_59752;
wire x_59753;
wire x_59754;
wire x_59755;
wire x_59756;
wire x_59757;
wire x_59758;
wire x_59759;
wire x_59760;
wire x_59761;
wire x_59762;
wire x_59763;
wire x_59764;
wire x_59765;
wire x_59766;
wire x_59767;
wire x_59768;
wire x_59769;
wire x_59770;
wire x_59771;
wire x_59772;
wire x_59773;
wire x_59774;
wire x_59775;
wire x_59776;
wire x_59777;
wire x_59778;
wire x_59779;
wire x_59780;
wire x_59781;
wire x_59782;
wire x_59783;
wire x_59784;
wire x_59785;
wire x_59786;
wire x_59787;
wire x_59788;
wire x_59789;
wire x_59790;
wire x_59791;
wire x_59792;
wire x_59793;
wire x_59794;
wire x_59795;
wire x_59796;
wire x_59797;
wire x_59798;
wire x_59799;
wire x_59800;
wire x_59801;
wire x_59802;
wire x_59803;
wire x_59804;
wire x_59805;
wire x_59806;
wire x_59807;
wire x_59808;
wire x_59809;
wire x_59810;
wire x_59811;
wire x_59812;
wire x_59813;
wire x_59814;
wire x_59815;
wire x_59816;
wire x_59817;
wire x_59818;
wire x_59819;
wire x_59820;
wire x_59821;
wire x_59822;
wire x_59823;
wire x_59824;
wire x_59825;
wire x_59826;
wire x_59827;
wire x_59828;
wire x_59829;
wire x_59830;
wire x_59831;
wire x_59832;
wire x_59833;
wire x_59834;
wire x_59835;
wire x_59836;
wire x_59837;
wire x_59838;
wire x_59839;
wire x_59840;
wire x_59841;
wire x_59842;
wire x_59843;
wire x_59844;
wire x_59845;
wire x_59846;
wire x_59847;
wire x_59848;
wire x_59849;
wire x_59850;
wire x_59851;
wire x_59852;
wire x_59853;
wire x_59854;
wire x_59855;
wire x_59856;
wire x_59857;
wire x_59858;
wire x_59859;
wire x_59860;
wire x_59861;
wire x_59862;
wire x_59863;
wire x_59864;
wire x_59865;
wire x_59866;
wire x_59867;
wire x_59868;
wire x_59869;
wire x_59870;
wire x_59871;
wire x_59872;
wire x_59873;
wire x_59874;
wire x_59875;
wire x_59876;
wire x_59877;
wire x_59878;
wire x_59879;
wire x_59880;
wire x_59881;
wire x_59882;
wire x_59883;
wire x_59884;
wire x_59885;
wire x_59886;
wire x_59887;
wire x_59888;
wire x_59889;
wire x_59890;
wire x_59891;
wire x_59892;
wire x_59893;
wire x_59894;
wire x_59895;
wire x_59896;
wire x_59897;
wire x_59898;
wire x_59899;
wire x_59900;
wire x_59901;
wire x_59902;
wire x_59903;
wire x_59904;
wire x_59905;
wire x_59906;
wire x_59907;
wire x_59908;
wire x_59909;
wire x_59910;
wire x_59911;
wire x_59912;
wire x_59913;
wire x_59914;
wire x_59915;
wire x_59916;
wire x_59917;
wire x_59918;
wire x_59919;
wire x_59920;
wire x_59921;
wire x_59922;
wire x_59923;
wire x_59924;
wire x_59925;
wire x_59926;
wire x_59927;
wire x_59928;
wire x_59929;
wire x_59930;
wire x_59931;
wire x_59932;
wire x_59933;
wire x_59934;
wire x_59935;
wire x_59936;
wire x_59937;
wire x_59938;
wire x_59939;
wire x_59940;
wire x_59941;
wire x_59942;
wire x_59943;
wire x_59944;
wire x_59945;
wire x_59946;
wire x_59947;
wire x_59948;
wire x_59949;
wire x_59950;
wire x_59951;
wire x_59952;
wire x_59953;
wire x_59954;
wire x_59955;
wire x_59956;
wire x_59957;
wire x_59958;
wire x_59959;
wire x_59960;
wire x_59961;
wire x_59962;
wire x_59963;
wire x_59964;
wire x_59965;
wire x_59966;
wire x_59967;
wire x_59968;
wire x_59969;
wire x_59970;
wire x_59971;
wire x_59972;
wire x_59973;
wire x_59974;
wire x_59975;
wire x_59976;
wire x_59977;
wire x_59978;
wire x_59979;
wire x_59980;
wire x_59981;
wire x_59982;
wire x_59983;
wire x_59984;
wire x_59985;
wire x_59986;
wire x_59987;
wire x_59988;
wire x_59989;
wire x_59990;
wire x_59991;
wire x_59992;
wire x_59993;
wire x_59994;
wire x_59995;
wire x_59996;
wire x_59997;
wire x_59998;
wire x_59999;
wire x_60000;
wire x_60001;
wire x_60002;
wire x_60003;
wire x_60004;
wire x_60005;
wire x_60006;
wire x_60007;
wire x_60008;
wire x_60009;
wire x_60010;
wire x_60011;
wire x_60012;
wire x_60013;
wire x_60014;
wire x_60015;
wire x_60016;
wire x_60017;
wire x_60018;
wire x_60019;
wire x_60020;
wire x_60021;
wire x_60022;
wire x_60023;
wire x_60024;
wire x_60025;
wire x_60026;
wire x_60027;
wire x_60028;
wire x_60029;
wire x_60030;
wire x_60031;
wire x_60032;
wire x_60033;
wire x_60034;
wire x_60035;
wire x_60036;
wire x_60037;
wire x_60038;
wire x_60039;
wire x_60040;
wire x_60041;
wire x_60042;
wire x_60043;
wire x_60044;
wire x_60045;
wire x_60046;
wire x_60047;
wire x_60048;
wire x_60049;
wire x_60050;
wire x_60051;
wire x_60052;
wire x_60053;
wire x_60054;
wire x_60055;
wire x_60056;
wire x_60057;
wire x_60058;
wire x_60059;
wire x_60060;
wire x_60061;
wire x_60062;
wire x_60063;
wire x_60064;
wire x_60065;
wire x_60066;
wire x_60067;
wire x_60068;
wire x_60069;
wire x_60070;
wire x_60071;
wire x_60072;
wire x_60073;
wire x_60074;
wire x_60075;
wire x_60076;
wire x_60077;
wire x_60078;
wire x_60079;
wire x_60080;
wire x_60081;
wire x_60082;
wire x_60083;
wire x_60084;
wire x_60085;
wire x_60086;
wire x_60087;
wire x_60088;
wire x_60089;
wire x_60090;
wire x_60091;
wire x_60092;
wire x_60093;
wire x_60094;
wire x_60095;
wire x_60096;
wire x_60097;
wire x_60098;
wire x_60099;
wire x_60100;
wire x_60101;
wire x_60102;
wire x_60103;
wire x_60104;
wire x_60105;
wire x_60106;
wire x_60107;
wire x_60108;
wire x_60109;
wire x_60110;
wire x_60111;
wire x_60112;
wire x_60113;
wire x_60114;
wire x_60115;
wire x_60116;
wire x_60117;
wire x_60118;
wire x_60119;
wire x_60120;
wire x_60121;
wire x_60122;
wire x_60123;
wire x_60124;
wire x_60125;
wire x_60126;
wire x_60127;
wire x_60128;
wire x_60129;
wire x_60130;
wire x_60131;
wire x_60132;
wire x_60133;
wire x_60134;
wire x_60135;
wire x_60136;
wire x_60137;
wire x_60138;
wire x_60139;
wire x_60140;
wire x_60141;
wire x_60142;
wire x_60143;
wire x_60144;
wire x_60145;
wire x_60146;
wire x_60147;
wire x_60148;
wire x_60149;
wire x_60150;
wire x_60151;
wire x_60152;
wire x_60153;
wire x_60154;
wire x_60155;
wire x_60156;
wire x_60157;
wire x_60158;
wire x_60159;
wire x_60160;
wire x_60161;
wire x_60162;
wire x_60163;
wire x_60164;
wire x_60165;
wire x_60166;
wire x_60167;
wire x_60168;
wire x_60169;
wire x_60170;
wire x_60171;
wire x_60172;
wire x_60173;
wire x_60174;
wire x_60175;
wire x_60176;
wire x_60177;
wire x_60178;
wire x_60179;
wire x_60180;
wire x_60181;
wire x_60182;
wire x_60183;
wire x_60184;
wire x_60185;
wire x_60186;
wire x_60187;
wire x_60188;
wire x_60189;
wire x_60190;
wire x_60191;
wire x_60192;
wire x_60193;
wire x_60194;
wire x_60195;
wire x_60196;
wire x_60197;
wire x_60198;
wire x_60199;
wire x_60200;
wire x_60201;
wire x_60202;
wire x_60203;
wire x_60204;
wire x_60205;
wire x_60206;
wire x_60207;
wire x_60208;
wire x_60209;
wire x_60210;
wire x_60211;
wire x_60212;
wire x_60213;
wire x_60214;
wire x_60215;
wire x_60216;
wire x_60217;
wire x_60218;
wire x_60219;
wire x_60220;
wire x_60221;
wire x_60222;
wire x_60223;
wire x_60224;
wire x_60225;
wire x_60226;
wire x_60227;
wire x_60228;
wire x_60229;
wire x_60230;
wire x_60231;
wire x_60232;
wire x_60233;
wire x_60234;
wire x_60235;
wire x_60236;
wire x_60237;
wire x_60238;
wire x_60239;
wire x_60240;
wire x_60241;
wire x_60242;
wire x_60243;
wire x_60244;
wire x_60245;
wire x_60246;
wire x_60247;
wire x_60248;
wire x_60249;
wire x_60250;
wire x_60251;
wire x_60252;
wire x_60253;
wire x_60254;
wire x_60255;
wire x_60256;
wire x_60257;
wire x_60258;
wire x_60259;
wire x_60260;
wire x_60261;
wire x_60262;
wire x_60263;
wire x_60264;
wire x_60265;
wire x_60266;
wire x_60267;
wire x_60268;
wire x_60269;
wire x_60270;
wire x_60271;
wire x_60272;
wire x_60273;
wire x_60274;
wire x_60275;
wire x_60276;
wire x_60277;
wire x_60278;
wire x_60279;
wire x_60280;
wire x_60281;
wire x_60282;
wire x_60283;
wire x_60284;
wire x_60285;
wire x_60286;
wire x_60287;
wire x_60288;
wire x_60289;
wire x_60290;
wire x_60291;
wire x_60292;
wire x_60293;
wire x_60294;
wire x_60295;
wire x_60296;
wire x_60297;
wire x_60298;
wire x_60299;
wire x_60300;
wire x_60301;
wire x_60302;
wire x_60303;
wire x_60304;
wire x_60305;
wire x_60306;
wire x_60307;
wire x_60308;
wire x_60309;
wire x_60310;
wire x_60311;
wire x_60312;
wire x_60313;
wire x_60314;
wire x_60315;
wire x_60316;
wire x_60317;
wire x_60318;
wire x_60319;
wire x_60320;
wire x_60321;
wire x_60322;
wire x_60323;
wire x_60324;
wire x_60325;
wire x_60326;
wire x_60327;
wire x_60328;
wire x_60329;
wire x_60330;
wire x_60331;
wire x_60332;
wire x_60333;
wire x_60334;
wire x_60335;
wire x_60336;
wire x_60337;
wire x_60338;
wire x_60339;
wire x_60340;
wire x_60341;
wire x_60342;
wire x_60343;
wire x_60344;
wire x_60345;
wire x_60346;
wire x_60347;
wire x_60348;
wire x_60349;
wire x_60350;
wire x_60351;
wire x_60352;
wire x_60353;
wire x_60354;
wire x_60355;
wire x_60356;
wire x_60357;
wire x_60358;
wire x_60359;
wire x_60360;
wire x_60361;
wire x_60362;
wire x_60363;
wire x_60364;
wire x_60365;
wire x_60366;
wire x_60367;
wire x_60368;
wire x_60369;
wire x_60370;
wire x_60371;
wire x_60372;
wire x_60373;
wire x_60374;
wire x_60375;
wire x_60376;
wire x_60377;
wire x_60378;
wire x_60379;
wire x_60380;
wire x_60381;
wire x_60382;
wire x_60383;
wire x_60384;
wire x_60385;
wire x_60386;
wire x_60387;
wire x_60388;
wire x_60389;
wire x_60390;
wire x_60391;
wire x_60392;
wire x_60393;
wire x_60394;
wire x_60395;
wire x_60396;
wire x_60397;
wire x_60398;
wire x_60399;
wire x_60400;
wire x_60401;
wire x_60402;
wire x_60403;
wire x_60404;
wire x_60405;
wire x_60406;
wire x_60407;
wire x_60408;
wire x_60409;
wire x_60410;
wire x_60411;
wire x_60412;
wire x_60413;
wire x_60414;
wire x_60415;
wire x_60416;
wire x_60417;
wire x_60418;
wire x_60419;
wire x_60420;
wire x_60421;
wire x_60422;
wire x_60423;
wire x_60424;
wire x_60425;
wire x_60426;
wire x_60427;
wire x_60428;
wire x_60429;
wire x_60430;
wire x_60431;
wire x_60432;
wire x_60433;
wire x_60434;
wire x_60435;
wire x_60436;
wire x_60437;
wire x_60438;
wire x_60439;
wire x_60440;
wire x_60441;
wire x_60442;
wire x_60443;
wire x_60444;
wire x_60445;
wire x_60446;
wire x_60447;
wire x_60448;
wire x_60449;
wire x_60450;
wire x_60451;
wire x_60452;
wire x_60453;
wire x_60454;
wire x_60455;
wire x_60456;
wire x_60457;
wire x_60458;
wire x_60459;
wire x_60460;
wire x_60461;
wire x_60462;
wire x_60463;
wire x_60464;
wire x_60465;
wire x_60466;
wire x_60467;
wire x_60468;
wire x_60469;
wire x_60470;
wire x_60471;
wire x_60472;
wire x_60473;
wire x_60474;
wire x_60475;
wire x_60476;
wire x_60477;
wire x_60478;
wire x_60479;
wire x_60480;
wire x_60481;
wire x_60482;
wire x_60483;
wire x_60484;
wire x_60485;
wire x_60486;
wire x_60487;
wire x_60488;
wire x_60489;
wire x_60490;
wire x_60491;
wire x_60492;
wire x_60493;
wire x_60494;
wire x_60495;
wire x_60496;
wire x_60497;
wire x_60498;
wire x_60499;
wire x_60500;
wire x_60501;
wire x_60502;
wire x_60503;
wire x_60504;
wire x_60505;
wire x_60506;
wire x_60507;
wire x_60508;
wire x_60509;
wire x_60510;
wire x_60511;
wire x_60512;
wire x_60513;
wire x_60514;
wire x_60515;
wire x_60516;
wire x_60517;
wire x_60518;
wire x_60519;
wire x_60520;
wire x_60521;
wire x_60522;
wire x_60523;
wire x_60524;
wire x_60525;
wire x_60526;
wire x_60527;
wire x_60528;
wire x_60529;
wire x_60530;
wire x_60531;
wire x_60532;
wire x_60533;
wire x_60534;
wire x_60535;
wire x_60536;
wire x_60537;
wire x_60538;
wire x_60539;
wire x_60540;
wire x_60541;
wire x_60542;
wire x_60543;
wire x_60544;
wire x_60545;
wire x_60546;
wire x_60547;
wire x_60548;
wire x_60549;
wire x_60550;
wire x_60551;
wire x_60552;
wire x_60553;
wire x_60554;
wire x_60555;
wire x_60556;
wire x_60557;
wire x_60558;
wire x_60559;
wire x_60560;
wire x_60561;
wire x_60562;
wire x_60563;
wire x_60564;
wire x_60565;
wire x_60566;
wire x_60567;
wire x_60568;
wire x_60569;
wire x_60570;
wire x_60571;
wire x_60572;
wire x_60573;
wire x_60574;
wire x_60575;
wire x_60576;
wire x_60577;
wire x_60578;
wire x_60579;
wire x_60580;
wire x_60581;
wire x_60582;
wire x_60583;
wire x_60584;
wire x_60585;
wire x_60586;
wire x_60587;
wire x_60588;
wire x_60589;
wire x_60590;
wire x_60591;
wire x_60592;
wire x_60593;
wire x_60594;
wire x_60595;
wire x_60596;
wire x_60597;
wire x_60598;
wire x_60599;
wire x_60600;
wire x_60601;
wire x_60602;
wire x_60603;
wire x_60604;
wire x_60605;
wire x_60606;
wire x_60607;
wire x_60608;
wire x_60609;
wire x_60610;
wire x_60611;
wire x_60612;
wire x_60613;
wire x_60614;
wire x_60615;
wire x_60616;
wire x_60617;
wire x_60618;
wire x_60619;
wire x_60620;
wire x_60621;
wire x_60622;
wire x_60623;
wire x_60624;
wire x_60625;
wire x_60626;
wire x_60627;
wire x_60628;
wire x_60629;
wire x_60630;
wire x_60631;
wire x_60632;
wire x_60633;
wire x_60634;
wire x_60635;
wire x_60636;
wire x_60637;
wire x_60638;
wire x_60639;
wire x_60640;
wire x_60641;
wire x_60642;
wire x_60643;
wire x_60644;
wire x_60645;
wire x_60646;
wire x_60647;
wire x_60648;
wire x_60649;
wire x_60650;
wire x_60651;
wire x_60652;
wire x_60653;
wire x_60654;
wire x_60655;
wire x_60656;
wire x_60657;
wire x_60658;
wire x_60659;
wire x_60660;
wire x_60661;
wire x_60662;
wire x_60663;
wire x_60664;
wire x_60665;
wire x_60666;
wire x_60667;
wire x_60668;
wire x_60669;
wire x_60670;
wire x_60671;
wire x_60672;
wire x_60673;
wire x_60674;
wire x_60675;
wire x_60676;
wire x_60677;
wire x_60678;
wire x_60679;
wire x_60680;
wire x_60681;
wire x_60682;
wire x_60683;
wire x_60684;
wire x_60685;
wire x_60686;
wire x_60687;
wire x_60688;
wire x_60689;
wire x_60690;
wire x_60691;
wire x_60692;
wire x_60693;
wire x_60694;
wire x_60695;
wire x_60696;
wire x_60697;
wire x_60698;
wire x_60699;
wire x_60700;
wire x_60701;
wire x_60702;
wire x_60703;
wire x_60704;
wire x_60705;
wire x_60706;
wire x_60707;
wire x_60708;
wire x_60709;
wire x_60710;
wire x_60711;
wire x_60712;
wire x_60713;
wire x_60714;
wire x_60715;
wire x_60716;
wire x_60717;
wire x_60718;
wire x_60719;
wire x_60720;
wire x_60721;
wire x_60722;
wire x_60723;
wire x_60724;
wire x_60725;
wire x_60726;
wire x_60727;
wire x_60728;
wire x_60729;
wire x_60730;
wire x_60731;
wire x_60732;
wire x_60733;
wire x_60734;
wire x_60735;
wire x_60736;
wire x_60737;
wire x_60738;
wire x_60739;
wire x_60740;
wire x_60741;
wire x_60742;
wire x_60743;
wire x_60744;
wire x_60745;
wire x_60746;
wire x_60747;
wire x_60748;
wire x_60749;
wire x_60750;
wire x_60751;
wire x_60752;
wire x_60753;
wire x_60754;
wire x_60755;
wire x_60756;
wire x_60757;
wire x_60758;
wire x_60759;
wire x_60760;
wire x_60761;
wire x_60762;
wire x_60763;
wire x_60764;
wire x_60765;
wire x_60766;
wire x_60767;
wire x_60768;
wire x_60769;
wire x_60770;
wire x_60771;
wire x_60772;
wire x_60773;
wire x_60774;
wire x_60775;
wire x_60776;
wire x_60777;
wire x_60778;
wire x_60779;
wire x_60780;
wire x_60781;
wire x_60782;
wire x_60783;
wire x_60784;
wire x_60785;
wire x_60786;
wire x_60787;
wire x_60788;
wire x_60789;
wire x_60790;
wire x_60791;
wire x_60792;
wire x_60793;
wire x_60794;
wire x_60795;
wire x_60796;
wire x_60797;
wire x_60798;
wire x_60799;
wire x_60800;
wire x_60801;
wire x_60802;
wire x_60803;
wire x_60804;
wire x_60805;
wire x_60806;
wire x_60807;
wire x_60808;
wire x_60809;
wire x_60810;
wire x_60811;
wire x_60812;
wire x_60813;
wire x_60814;
wire x_60815;
wire x_60816;
wire x_60817;
wire x_60818;
wire x_60819;
wire x_60820;
wire x_60821;
wire x_60822;
wire x_60823;
wire x_60824;
wire x_60825;
wire x_60826;
wire x_60827;
wire x_60828;
wire x_60829;
wire x_60830;
wire x_60831;
wire x_60832;
wire x_60833;
wire x_60834;
wire x_60835;
wire x_60836;
wire x_60837;
wire x_60838;
wire x_60839;
wire x_60840;
wire x_60841;
wire x_60842;
wire x_60843;
wire x_60844;
wire x_60845;
wire x_60846;
wire x_60847;
wire x_60848;
wire x_60849;
wire x_60850;
wire x_60851;
wire x_60852;
wire x_60853;
wire x_60854;
wire x_60855;
wire x_60856;
wire x_60857;
wire x_60858;
wire x_60859;
wire x_60860;
wire x_60861;
wire x_60862;
wire x_60863;
wire x_60864;
wire x_60865;
wire x_60866;
wire x_60867;
wire x_60868;
wire x_60869;
wire x_60870;
wire x_60871;
wire x_60872;
wire x_60873;
wire x_60874;
wire x_60875;
wire x_60876;
wire x_60877;
wire x_60878;
wire x_60879;
wire x_60880;
wire x_60881;
wire x_60882;
wire x_60883;
wire x_60884;
wire x_60885;
wire x_60886;
wire x_60887;
wire x_60888;
wire x_60889;
wire x_60890;
wire x_60891;
wire x_60892;
wire x_60893;
wire x_60894;
wire x_60895;
wire x_60896;
wire x_60897;
wire x_60898;
wire x_60899;
wire x_60900;
wire x_60901;
wire x_60902;
wire x_60903;
wire x_60904;
wire x_60905;
wire x_60906;
wire x_60907;
wire x_60908;
wire x_60909;
wire x_60910;
wire x_60911;
wire x_60912;
wire x_60913;
wire x_60914;
wire x_60915;
wire x_60916;
wire x_60917;
wire x_60918;
wire x_60919;
wire x_60920;
wire x_60921;
wire x_60922;
wire x_60923;
wire x_60924;
wire x_60925;
wire x_60926;
wire x_60927;
wire x_60928;
wire x_60929;
wire x_60930;
wire x_60931;
wire x_60932;
wire x_60933;
wire x_60934;
wire x_60935;
wire x_60936;
wire x_60937;
wire x_60938;
wire x_60939;
wire x_60940;
wire x_60941;
wire x_60942;
wire x_60943;
wire x_60944;
wire x_60945;
wire x_60946;
wire x_60947;
wire x_60948;
wire x_60949;
wire x_60950;
wire x_60951;
wire x_60952;
wire x_60953;
wire x_60954;
wire x_60955;
wire x_60956;
wire x_60957;
wire x_60958;
wire x_60959;
wire x_60960;
wire x_60961;
wire x_60962;
wire x_60963;
wire x_60964;
wire x_60965;
wire x_60966;
wire x_60967;
wire x_60968;
wire x_60969;
wire x_60970;
wire x_60971;
wire x_60972;
wire x_60973;
wire x_60974;
wire x_60975;
wire x_60976;
wire x_60977;
wire x_60978;
wire x_60979;
wire x_60980;
wire x_60981;
wire x_60982;
wire x_60983;
wire x_60984;
wire x_60985;
wire x_60986;
wire x_60987;
wire x_60988;
wire x_60989;
wire x_60990;
wire x_60991;
wire x_60992;
wire x_60993;
wire x_60994;
wire x_60995;
wire x_60996;
wire x_60997;
wire x_60998;
wire x_60999;
wire x_61000;
wire x_61001;
wire x_61002;
wire x_61003;
wire x_61004;
wire x_61005;
wire x_61006;
wire x_61007;
wire x_61008;
wire x_61009;
wire x_61010;
wire x_61011;
wire x_61012;
wire x_61013;
wire x_61014;
wire x_61015;
wire x_61016;
wire x_61017;
wire x_61018;
wire x_61019;
wire x_61020;
wire x_61021;
wire x_61022;
wire x_61023;
wire x_61024;
wire x_61025;
wire x_61026;
wire x_61027;
wire x_61028;
wire x_61029;
wire x_61030;
wire x_61031;
wire x_61032;
wire x_61033;
wire x_61034;
wire x_61035;
wire x_61036;
wire x_61037;
wire x_61038;
wire x_61039;
wire x_61040;
wire x_61041;
wire x_61042;
wire x_61043;
wire x_61044;
wire x_61045;
wire x_61046;
wire x_61047;
wire x_61048;
wire x_61049;
wire x_61050;
wire x_61051;
wire x_61052;
wire x_61053;
wire x_61054;
wire x_61055;
wire x_61056;
wire x_61057;
wire x_61058;
wire x_61059;
wire x_61060;
wire x_61061;
wire x_61062;
wire x_61063;
wire x_61064;
wire x_61065;
wire x_61066;
wire x_61067;
wire x_61068;
wire x_61069;
wire x_61070;
wire x_61071;
wire x_61072;
wire x_61073;
wire x_61074;
wire x_61075;
wire x_61076;
wire x_61077;
wire x_61078;
wire x_61079;
wire x_61080;
wire x_61081;
wire x_61082;
wire x_61083;
wire x_61084;
wire x_61085;
wire x_61086;
wire x_61087;
wire x_61088;
wire x_61089;
wire x_61090;
wire x_61091;
wire x_61092;
wire x_61093;
wire x_61094;
wire x_61095;
wire x_61096;
wire x_61097;
wire x_61098;
wire x_61099;
wire x_61100;
wire x_61101;
wire x_61102;
wire x_61103;
wire x_61104;
wire x_61105;
wire x_61106;
wire x_61107;
wire x_61108;
wire x_61109;
wire x_61110;
wire x_61111;
wire x_61112;
wire x_61113;
wire x_61114;
wire x_61115;
wire x_61116;
wire x_61117;
wire x_61118;
wire x_61119;
wire x_61120;
wire x_61121;
wire x_61122;
wire x_61123;
wire x_61124;
wire x_61125;
wire x_61126;
wire x_61127;
wire x_61128;
wire x_61129;
wire x_61130;
wire x_61131;
wire x_61132;
wire x_61133;
wire x_61134;
wire x_61135;
wire x_61136;
wire x_61137;
wire x_61138;
wire x_61139;
wire x_61140;
wire x_61141;
wire x_61142;
wire x_61143;
wire x_61144;
wire x_61145;
wire x_61146;
wire x_61147;
wire x_61148;
wire x_61149;
wire x_61150;
wire x_61151;
wire x_61152;
wire x_61153;
wire x_61154;
wire x_61155;
wire x_61156;
wire x_61157;
wire x_61158;
wire x_61159;
wire x_61160;
wire x_61161;
wire x_61162;
wire x_61163;
wire x_61164;
wire x_61165;
wire x_61166;
wire x_61167;
wire x_61168;
wire x_61169;
wire x_61170;
wire x_61171;
wire x_61172;
wire x_61173;
wire x_61174;
wire x_61175;
wire x_61176;
wire x_61177;
wire x_61178;
wire x_61179;
wire x_61180;
wire x_61181;
wire x_61182;
wire x_61183;
wire x_61184;
wire x_61185;
wire x_61186;
wire x_61187;
wire x_61188;
wire x_61189;
wire x_61190;
wire x_61191;
wire x_61192;
wire x_61193;
wire x_61194;
wire x_61195;
wire x_61196;
wire x_61197;
wire x_61198;
wire x_61199;
wire x_61200;
wire x_61201;
wire x_61202;
wire x_61203;
wire x_61204;
wire x_61205;
wire x_61206;
wire x_61207;
wire x_61208;
wire x_61209;
wire x_61210;
wire x_61211;
wire x_61212;
wire x_61213;
wire x_61214;
wire x_61215;
wire x_61216;
wire x_61217;
wire x_61218;
wire x_61219;
wire x_61220;
wire x_61221;
wire x_61222;
wire x_61223;
wire x_61224;
wire x_61225;
wire x_61226;
wire x_61227;
wire x_61228;
wire x_61229;
wire x_61230;
wire x_61231;
wire x_61232;
wire x_61233;
wire x_61234;
wire x_61235;
wire x_61236;
wire x_61237;
wire x_61238;
wire x_61239;
wire x_61240;
wire x_61241;
wire x_61242;
wire x_61243;
wire x_61244;
wire x_61245;
wire x_61246;
wire x_61247;
wire x_61248;
wire x_61249;
wire x_61250;
wire x_61251;
wire x_61252;
wire x_61253;
wire x_61254;
wire x_61255;
wire x_61256;
wire x_61257;
wire x_61258;
wire x_61259;
wire x_61260;
wire x_61261;
wire x_61262;
wire x_61263;
wire x_61264;
wire x_61265;
wire x_61266;
wire x_61267;
wire x_61268;
wire x_61269;
wire x_61270;
wire x_61271;
wire x_61272;
wire x_61273;
wire x_61274;
wire x_61275;
wire x_61276;
wire x_61277;
wire x_61278;
wire x_61279;
wire x_61280;
wire x_61281;
wire x_61282;
wire x_61283;
wire x_61284;
wire x_61285;
wire x_61286;
wire x_61287;
wire x_61288;
wire x_61289;
wire x_61290;
wire x_61291;
wire x_61292;
wire x_61293;
wire x_61294;
wire x_61295;
wire x_61296;
wire x_61297;
wire x_61298;
wire x_61299;
wire x_61300;
wire x_61301;
wire x_61302;
wire x_61303;
wire x_61304;
wire x_61305;
wire x_61306;
wire x_61307;
wire x_61308;
wire x_61309;
wire x_61310;
wire x_61311;
wire x_61312;
wire x_61313;
wire x_61314;
wire x_61315;
wire x_61316;
wire x_61317;
wire x_61318;
wire x_61319;
wire x_61320;
wire x_61321;
wire x_61322;
wire x_61323;
wire x_61324;
wire x_61325;
wire x_61326;
wire x_61327;
wire x_61328;
wire x_61329;
wire x_61330;
wire x_61331;
wire x_61332;
wire x_61333;
wire x_61334;
wire x_61335;
wire x_61336;
wire x_61337;
wire x_61338;
wire x_61339;
wire x_61340;
wire x_61341;
wire x_61342;
wire x_61343;
wire x_61344;
wire x_61345;
wire x_61346;
wire x_61347;
wire x_61348;
wire x_61349;
wire x_61350;
wire x_61351;
wire x_61352;
wire x_61353;
wire x_61354;
wire x_61355;
wire x_61356;
wire x_61357;
wire x_61358;
wire x_61359;
wire x_61360;
wire x_61361;
wire x_61362;
wire x_61363;
wire x_61364;
wire x_61365;
wire x_61366;
wire x_61367;
wire x_61368;
wire x_61369;
wire x_61370;
wire x_61371;
wire x_61372;
wire x_61373;
wire x_61374;
wire x_61375;
wire x_61376;
wire x_61377;
wire x_61378;
wire x_61379;
wire x_61380;
wire x_61381;
wire x_61382;
wire x_61383;
wire x_61384;
wire x_61385;
wire x_61386;
wire x_61387;
wire x_61388;
wire x_61389;
wire x_61390;
wire x_61391;
wire x_61392;
wire x_61393;
wire x_61394;
wire x_61395;
wire x_61396;
wire x_61397;
wire x_61398;
wire x_61399;
wire x_61400;
wire x_61401;
wire x_61402;
wire x_61403;
wire x_61404;
wire x_61405;
wire x_61406;
wire x_61407;
wire x_61408;
wire x_61409;
wire x_61410;
wire x_61411;
wire x_61412;
wire x_61413;
wire x_61414;
wire x_61415;
wire x_61416;
wire x_61417;
wire x_61418;
wire x_61419;
wire x_61420;
wire x_61421;
wire x_61422;
wire x_61423;
wire x_61424;
wire x_61425;
wire x_61426;
wire x_61427;
wire x_61428;
wire x_61429;
wire x_61430;
wire x_61431;
wire x_61432;
wire x_61433;
wire x_61434;
wire x_61435;
wire x_61436;
wire x_61437;
wire x_61438;
wire x_61439;
wire x_61440;
wire x_61441;
wire x_61442;
wire x_61443;
wire x_61444;
wire x_61445;
wire x_61446;
wire x_61447;
wire x_61448;
wire x_61449;
wire x_61450;
wire x_61451;
wire x_61452;
wire x_61453;
wire x_61454;
wire x_61455;
wire x_61456;
wire x_61457;
wire x_61458;
wire x_61459;
wire x_61460;
wire x_61461;
wire x_61462;
wire x_61463;
wire x_61464;
wire x_61465;
wire x_61466;
wire x_61467;
wire x_61468;
wire x_61469;
wire x_61470;
wire x_61471;
wire x_61472;
wire x_61473;
wire x_61474;
wire x_61475;
wire x_61476;
wire x_61477;
wire x_61478;
wire x_61479;
wire x_61480;
wire x_61481;
wire x_61482;
wire x_61483;
wire x_61484;
wire x_61485;
wire x_61486;
wire x_61487;
wire x_61488;
wire x_61489;
wire x_61490;
wire x_61491;
wire x_61492;
wire x_61493;
wire x_61494;
wire x_61495;
wire x_61496;
wire x_61497;
wire x_61498;
wire x_61499;
wire x_61500;
wire x_61501;
wire x_61502;
wire x_61503;
wire x_61504;
wire x_61505;
wire x_61506;
wire x_61507;
wire x_61508;
wire x_61509;
wire x_61510;
wire x_61511;
wire x_61512;
wire x_61513;
wire x_61514;
wire x_61515;
wire x_61516;
wire x_61517;
wire x_61518;
wire x_61519;
wire x_61520;
wire x_61521;
wire x_61522;
wire x_61523;
wire x_61524;
wire x_61525;
wire x_61526;
wire x_61527;
wire x_61528;
wire x_61529;
wire x_61530;
wire x_61531;
wire x_61532;
wire x_61533;
wire x_61534;
wire x_61535;
wire x_61536;
wire x_61537;
wire x_61538;
wire x_61539;
wire x_61540;
wire x_61541;
wire x_61542;
wire x_61543;
wire x_61544;
wire x_61545;
wire x_61546;
wire x_61547;
wire x_61548;
wire x_61549;
wire x_61550;
wire x_61551;
wire x_61552;
wire x_61553;
wire x_61554;
wire x_61555;
wire x_61556;
wire x_61557;
wire x_61558;
wire x_61559;
wire x_61560;
wire x_61561;
wire x_61562;
wire x_61563;
wire x_61564;
wire x_61565;
wire x_61566;
wire x_61567;
wire x_61568;
wire x_61569;
wire x_61570;
wire x_61571;
wire x_61572;
wire x_61573;
wire x_61574;
wire x_61575;
wire x_61576;
wire x_61577;
wire x_61578;
wire x_61579;
wire x_61580;
wire x_61581;
wire x_61582;
wire x_61583;
wire x_61584;
wire x_61585;
wire x_61586;
wire x_61587;
wire x_61588;
wire x_61589;
wire x_61590;
wire x_61591;
wire x_61592;
wire x_61593;
wire x_61594;
wire x_61595;
wire x_61596;
wire x_61597;
wire x_61598;
wire x_61599;
wire x_61600;
wire x_61601;
wire x_61602;
wire x_61603;
wire x_61604;
wire x_61605;
wire x_61606;
wire x_61607;
wire x_61608;
wire x_61609;
wire x_61610;
wire x_61611;
wire x_61612;
wire x_61613;
wire x_61614;
wire x_61615;
wire x_61616;
wire x_61617;
wire x_61618;
wire x_61619;
wire x_61620;
wire x_61621;
wire x_61622;
wire x_61623;
wire x_61624;
wire x_61625;
wire x_61626;
wire x_61627;
wire x_61628;
wire x_61629;
wire x_61630;
wire x_61631;
wire x_61632;
wire x_61633;
wire x_61634;
wire x_61635;
wire x_61636;
wire x_61637;
wire x_61638;
wire x_61639;
wire x_61640;
wire x_61641;
wire x_61642;
wire x_61643;
wire x_61644;
wire x_61645;
wire x_61646;
wire x_61647;
wire x_61648;
wire x_61649;
wire x_61650;
wire x_61651;
wire x_61652;
wire x_61653;
wire x_61654;
wire x_61655;
wire x_61656;
wire x_61657;
wire x_61658;
wire x_61659;
wire x_61660;
wire x_61661;
wire x_61662;
wire x_61663;
wire x_61664;
wire x_61665;
wire x_61666;
wire x_61667;
wire x_61668;
wire x_61669;
wire x_61670;
wire x_61671;
wire x_61672;
wire x_61673;
wire x_61674;
wire x_61675;
wire x_61676;
wire x_61677;
wire x_61678;
wire x_61679;
wire x_61680;
wire x_61681;
wire x_61682;
wire x_61683;
wire x_61684;
wire x_61685;
wire x_61686;
wire x_61687;
wire x_61688;
wire x_61689;
wire x_61690;
wire x_61691;
wire x_61692;
wire x_61693;
wire x_61694;
wire x_61695;
wire x_61696;
wire x_61697;
wire x_61698;
wire x_61699;
wire x_61700;
wire x_61701;
wire x_61702;
wire x_61703;
wire x_61704;
wire x_61705;
wire x_61706;
wire x_61707;
wire x_61708;
wire x_61709;
wire x_61710;
wire x_61711;
wire x_61712;
wire x_61713;
wire x_61714;
wire x_61715;
wire x_61716;
wire x_61717;
wire x_61718;
wire x_61719;
wire x_61720;
wire x_61721;
wire x_61722;
wire x_61723;
wire x_61724;
wire x_61725;
wire x_61726;
wire x_61727;
wire x_61728;
wire x_61729;
wire x_61730;
wire x_61731;
wire x_61732;
wire x_61733;
wire x_61734;
wire x_61735;
wire x_61736;
wire x_61737;
wire x_61738;
wire x_61739;
wire x_61740;
wire x_61741;
wire x_61742;
wire x_61743;
wire x_61744;
wire x_61745;
wire x_61746;
wire x_61747;
wire x_61748;
wire x_61749;
wire x_61750;
wire x_61751;
wire x_61752;
wire x_61753;
wire x_61754;
wire x_61755;
wire x_61756;
wire x_61757;
wire x_61758;
wire x_61759;
wire x_61760;
wire x_61761;
wire x_61762;
wire x_61763;
wire x_61764;
wire x_61765;
wire x_61766;
wire x_61767;
wire x_61768;
wire x_61769;
wire x_61770;
wire x_61771;
wire x_61772;
wire x_61773;
wire x_61774;
wire x_61775;
wire x_61776;
wire x_61777;
wire x_61778;
wire x_61779;
wire x_61780;
wire x_61781;
wire x_61782;
wire x_61783;
wire x_61784;
wire x_61785;
wire x_61786;
wire x_61787;
wire x_61788;
wire x_61789;
wire x_61790;
wire x_61791;
wire x_61792;
wire x_61793;
wire x_61794;
wire x_61795;
wire x_61796;
wire x_61797;
wire x_61798;
wire x_61799;
wire x_61800;
wire x_61801;
wire x_61802;
wire x_61803;
wire x_61804;
wire x_61805;
wire x_61806;
wire x_61807;
wire x_61808;
wire x_61809;
wire x_61810;
wire x_61811;
wire x_61812;
wire x_61813;
wire x_61814;
wire x_61815;
wire x_61816;
wire x_61817;
wire x_61818;
wire x_61819;
wire x_61820;
wire x_61821;
wire x_61822;
wire x_61823;
wire x_61824;
wire x_61825;
wire x_61826;
wire x_61827;
wire x_61828;
wire x_61829;
wire x_61830;
wire x_61831;
wire x_61832;
wire x_61833;
wire x_61834;
wire x_61835;
wire x_61836;
wire x_61837;
wire x_61838;
wire x_61839;
wire x_61840;
wire x_61841;
wire x_61842;
wire x_61843;
wire x_61844;
wire x_61845;
wire x_61846;
wire x_61847;
wire x_61848;
wire x_61849;
wire x_61850;
wire x_61851;
wire x_61852;
wire x_61853;
wire x_61854;
wire x_61855;
wire x_61856;
wire x_61857;
wire x_61858;
wire x_61859;
wire x_61860;
wire x_61861;
wire x_61862;
wire x_61863;
wire x_61864;
wire x_61865;
wire x_61866;
wire x_61867;
wire x_61868;
wire x_61869;
wire x_61870;
wire x_61871;
wire x_61872;
wire x_61873;
wire x_61874;
wire x_61875;
wire x_61876;
wire x_61877;
wire x_61878;
wire x_61879;
wire x_61880;
wire x_61881;
wire x_61882;
wire x_61883;
wire x_61884;
wire x_61885;
wire x_61886;
wire x_61887;
wire x_61888;
wire x_61889;
wire x_61890;
wire x_61891;
wire x_61892;
wire x_61893;
wire x_61894;
wire x_61895;
wire x_61896;
wire x_61897;
wire x_61898;
wire x_61899;
wire x_61900;
wire x_61901;
wire x_61902;
wire x_61903;
wire x_61904;
wire x_61905;
wire x_61906;
wire x_61907;
wire x_61908;
wire x_61909;
wire x_61910;
wire x_61911;
wire x_61912;
wire x_61913;
wire x_61914;
wire x_61915;
wire x_61916;
wire x_61917;
wire x_61918;
wire x_61919;
wire x_61920;
wire x_61921;
wire x_61922;
wire x_61923;
wire x_61924;
wire x_61925;
wire x_61926;
wire x_61927;
wire x_61928;
wire x_61929;
wire x_61930;
wire x_61931;
wire x_61932;
wire x_61933;
wire x_61934;
wire x_61935;
wire x_61936;
wire x_61937;
wire x_61938;
wire x_61939;
wire x_61940;
wire x_61941;
wire x_61942;
wire x_61943;
wire x_61944;
wire x_61945;
wire x_61946;
wire x_61947;
wire x_61948;
wire x_61949;
wire x_61950;
wire x_61951;
wire x_61952;
wire x_61953;
wire x_61954;
wire x_61955;
wire x_61956;
wire x_61957;
wire x_61958;
wire x_61959;
wire x_61960;
wire x_61961;
wire x_61962;
wire x_61963;
wire x_61964;
wire x_61965;
wire x_61966;
wire x_61967;
wire x_61968;
wire x_61969;
wire x_61970;
wire x_61971;
wire x_61972;
wire x_61973;
wire x_61974;
wire x_61975;
wire x_61976;
wire x_61977;
wire x_61978;
wire x_61979;
wire x_61980;
wire x_61981;
wire x_61982;
wire x_61983;
wire x_61984;
wire x_61985;
wire x_61986;
wire x_61987;
wire x_61988;
wire x_61989;
wire x_61990;
wire x_61991;
wire x_61992;
wire x_61993;
wire x_61994;
wire x_61995;
wire x_61996;
wire x_61997;
wire x_61998;
wire x_61999;
wire x_62000;
wire x_62001;
wire x_62002;
wire x_62003;
wire x_62004;
wire x_62005;
wire x_62006;
wire x_62007;
wire x_62008;
wire x_62009;
wire x_62010;
wire x_62011;
wire x_62012;
wire x_62013;
wire x_62014;
wire x_62015;
wire x_62016;
wire x_62017;
wire x_62018;
wire x_62019;
wire x_62020;
wire x_62021;
wire x_62022;
wire x_62023;
wire x_62024;
wire x_62025;
wire x_62026;
wire x_62027;
wire x_62028;
wire x_62029;
wire x_62030;
wire x_62031;
wire x_62032;
wire x_62033;
wire x_62034;
wire x_62035;
wire x_62036;
wire x_62037;
wire x_62038;
wire x_62039;
wire x_62040;
wire x_62041;
wire x_62042;
wire x_62043;
wire x_62044;
wire x_62045;
wire x_62046;
wire x_62047;
wire x_62048;
wire x_62049;
wire x_62050;
wire x_62051;
wire x_62052;
wire x_62053;
wire x_62054;
wire x_62055;
wire x_62056;
wire x_62057;
wire x_62058;
wire x_62059;
wire x_62060;
wire x_62061;
wire x_62062;
wire x_62063;
wire x_62064;
wire x_62065;
wire x_62066;
wire x_62067;
wire x_62068;
wire x_62069;
wire x_62070;
wire x_62071;
wire x_62072;
wire x_62073;
wire x_62074;
wire x_62075;
wire x_62076;
wire x_62077;
wire x_62078;
wire x_62079;
wire x_62080;
wire x_62081;
wire x_62082;
wire x_62083;
wire x_62084;
wire x_62085;
wire x_62086;
wire x_62087;
wire x_62088;
wire x_62089;
wire x_62090;
wire x_62091;
wire x_62092;
wire x_62093;
wire x_62094;
wire x_62095;
wire x_62096;
wire x_62097;
wire x_62098;
wire x_62099;
wire x_62100;
wire x_62101;
wire x_62102;
wire x_62103;
wire x_62104;
wire x_62105;
wire x_62106;
wire x_62107;
wire x_62108;
wire x_62109;
wire x_62110;
wire x_62111;
wire x_62112;
wire x_62113;
wire x_62114;
wire x_62115;
wire x_62116;
wire x_62117;
wire x_62118;
wire x_62119;
wire x_62120;
wire x_62121;
wire x_62122;
wire x_62123;
wire x_62124;
wire x_62125;
wire x_62126;
wire x_62127;
wire x_62128;
wire x_62129;
wire x_62130;
wire x_62131;
wire x_62132;
wire x_62133;
wire x_62134;
wire x_62135;
wire x_62136;
wire x_62137;
wire x_62138;
wire x_62139;
wire x_62140;
wire x_62141;
wire x_62142;
wire x_62143;
wire x_62144;
wire x_62145;
wire x_62146;
wire x_62147;
wire x_62148;
wire x_62149;
wire x_62150;
wire x_62151;
wire x_62152;
wire x_62153;
wire x_62154;
wire x_62155;
wire x_62156;
wire x_62157;
wire x_62158;
wire x_62159;
wire x_62160;
wire x_62161;
wire x_62162;
wire x_62163;
wire x_62164;
wire x_62165;
wire x_62166;
wire x_62167;
wire x_62168;
wire x_62169;
wire x_62170;
wire x_62171;
wire x_62172;
wire x_62173;
wire x_62174;
wire x_62175;
wire x_62176;
wire x_62177;
wire x_62178;
wire x_62179;
wire x_62180;
wire x_62181;
wire x_62182;
wire x_62183;
wire x_62184;
wire x_62185;
wire x_62186;
wire x_62187;
wire x_62188;
wire x_62189;
wire x_62190;
wire x_62191;
wire x_62192;
wire x_62193;
wire x_62194;
wire x_62195;
wire x_62196;
wire x_62197;
wire x_62198;
wire x_62199;
wire x_62200;
wire x_62201;
wire x_62202;
wire x_62203;
wire x_62204;
wire x_62205;
wire x_62206;
wire x_62207;
wire x_62208;
wire x_62209;
wire x_62210;
wire x_62211;
wire x_62212;
wire x_62213;
wire x_62214;
wire x_62215;
wire x_62216;
wire x_62217;
wire x_62218;
wire x_62219;
wire x_62220;
wire x_62221;
wire x_62222;
wire x_62223;
wire x_62224;
wire x_62225;
wire x_62226;
wire x_62227;
wire x_62228;
wire x_62229;
wire x_62230;
wire x_62231;
wire x_62232;
wire x_62233;
wire x_62234;
wire x_62235;
wire x_62236;
wire x_62237;
wire x_62238;
wire x_62239;
wire x_62240;
wire x_62241;
wire x_62242;
wire x_62243;
wire x_62244;
wire x_62245;
wire x_62246;
wire x_62247;
wire x_62248;
wire x_62249;
wire x_62250;
wire x_62251;
wire x_62252;
wire x_62253;
wire x_62254;
wire x_62255;
wire x_62256;
wire x_62257;
wire x_62258;
wire x_62259;
wire x_62260;
wire x_62261;
wire x_62262;
wire x_62263;
wire x_62264;
wire x_62265;
wire x_62266;
wire x_62267;
wire x_62268;
wire x_62269;
wire x_62270;
wire x_62271;
wire x_62272;
wire x_62273;
wire x_62274;
wire x_62275;
wire x_62276;
wire x_62277;
wire x_62278;
wire x_62279;
wire x_62280;
wire x_62281;
wire x_62282;
wire x_62283;
wire x_62284;
wire x_62285;
wire x_62286;
wire x_62287;
wire x_62288;
wire x_62289;
wire x_62290;
wire x_62291;
wire x_62292;
wire x_62293;
wire x_62294;
wire x_62295;
wire x_62296;
wire x_62297;
wire x_62298;
wire x_62299;
wire x_62300;
wire x_62301;
wire x_62302;
wire x_62303;
wire x_62304;
wire x_62305;
wire x_62306;
wire x_62307;
wire x_62308;
wire x_62309;
wire x_62310;
wire x_62311;
wire x_62312;
wire x_62313;
wire x_62314;
wire x_62315;
wire x_62316;
wire x_62317;
wire x_62318;
wire x_62319;
wire x_62320;
wire x_62321;
wire x_62322;
wire x_62323;
wire x_62324;
wire x_62325;
wire x_62326;
wire x_62327;
wire x_62328;
wire x_62329;
wire x_62330;
wire x_62331;
wire x_62332;
wire x_62333;
wire x_62334;
wire x_62335;
wire x_62336;
wire x_62337;
wire x_62338;
wire x_62339;
wire x_62340;
wire x_62341;
wire x_62342;
wire x_62343;
wire x_62344;
wire x_62345;
wire x_62346;
wire x_62347;
wire x_62348;
wire x_62349;
wire x_62350;
wire x_62351;
wire x_62352;
wire x_62353;
wire x_62354;
wire x_62355;
wire x_62356;
wire x_62357;
wire x_62358;
wire x_62359;
wire x_62360;
wire x_62361;
wire x_62362;
wire x_62363;
wire x_62364;
wire x_62365;
wire x_62366;
wire x_62367;
wire x_62368;
wire x_62369;
wire x_62370;
wire x_62371;
wire x_62372;
wire x_62373;
wire x_62374;
wire x_62375;
wire x_62376;
wire x_62377;
wire x_62378;
wire x_62379;
wire x_62380;
wire x_62381;
wire x_62382;
wire x_62383;
wire x_62384;
wire x_62385;
wire x_62386;
wire x_62387;
wire x_62388;
wire x_62389;
wire x_62390;
wire x_62391;
wire x_62392;
wire x_62393;
wire x_62394;
wire x_62395;
wire x_62396;
wire x_62397;
wire x_62398;
wire x_62399;
wire x_62400;
wire x_62401;
wire x_62402;
wire x_62403;
wire x_62404;
wire x_62405;
wire x_62406;
wire x_62407;
wire x_62408;
wire x_62409;
wire x_62410;
wire x_62411;
wire x_62412;
wire x_62413;
wire x_62414;
wire x_62415;
wire x_62416;
wire x_62417;
wire x_62418;
wire x_62419;
wire x_62420;
wire x_62421;
wire x_62422;
wire x_62423;
wire x_62424;
wire x_62425;
wire x_62426;
wire x_62427;
wire x_62428;
wire x_62429;
wire x_62430;
wire x_62431;
wire x_62432;
wire x_62433;
wire x_62434;
wire x_62435;
wire x_62436;
wire x_62437;
wire x_62438;
wire x_62439;
wire x_62440;
wire x_62441;
wire x_62442;
wire x_62443;
wire x_62444;
wire x_62445;
wire x_62446;
wire x_62447;
wire x_62448;
wire x_62449;
wire x_62450;
wire x_62451;
wire x_62452;
wire x_62453;
wire x_62454;
wire x_62455;
wire x_62456;
wire x_62457;
wire x_62458;
wire x_62459;
wire x_62460;
wire x_62461;
wire x_62462;
wire x_62463;
wire x_62464;
wire x_62465;
wire x_62466;
wire x_62467;
wire x_62468;
wire x_62469;
wire x_62470;
wire x_62471;
wire x_62472;
wire x_62473;
wire x_62474;
wire x_62475;
wire x_62476;
wire x_62477;
wire x_62478;
wire x_62479;
wire x_62480;
wire x_62481;
wire x_62482;
wire x_62483;
wire x_62484;
wire x_62485;
wire x_62486;
wire x_62487;
wire x_62488;
wire x_62489;
wire x_62490;
wire x_62491;
wire x_62492;
wire x_62493;
wire x_62494;
wire x_62495;
wire x_62496;
wire x_62497;
wire x_62498;
wire x_62499;
wire x_62500;
wire x_62501;
wire x_62502;
wire x_62503;
wire x_62504;
wire x_62505;
wire x_62506;
wire x_62507;
wire x_62508;
wire x_62509;
wire x_62510;
wire x_62511;
wire x_62512;
wire x_62513;
wire x_62514;
wire x_62515;
wire x_62516;
wire x_62517;
wire x_62518;
wire x_62519;
wire x_62520;
wire x_62521;
wire x_62522;
wire x_62523;
wire x_62524;
wire x_62525;
wire x_62526;
wire x_62527;
wire x_62528;
wire x_62529;
wire x_62530;
wire x_62531;
wire x_62532;
wire x_62533;
wire x_62534;
wire x_62535;
wire x_62536;
wire x_62537;
wire x_62538;
wire x_62539;
wire x_62540;
wire x_62541;
wire x_62542;
wire x_62543;
wire x_62544;
wire x_62545;
wire x_62546;
wire x_62547;
wire x_62548;
wire x_62549;
wire x_62550;
wire x_62551;
wire x_62552;
wire x_62553;
wire x_62554;
wire x_62555;
wire x_62556;
wire x_62557;
wire x_62558;
wire x_62559;
wire x_62560;
wire x_62561;
wire x_62562;
wire x_62563;
wire x_62564;
wire x_62565;
wire x_62566;
wire x_62567;
wire x_62568;
wire x_62569;
wire x_62570;
wire x_62571;
wire x_62572;
wire x_62573;
wire x_62574;
wire x_62575;
wire x_62576;
wire x_62577;
wire x_62578;
wire x_62579;
wire x_62580;
wire x_62581;
wire x_62582;
wire x_62583;
wire x_62584;
wire x_62585;
wire x_62586;
wire x_62587;
wire x_62588;
wire x_62589;
wire x_62590;
wire x_62591;
wire x_62592;
wire x_62593;
assign v_4589 = 0;
assign x_1 = ~v_725 | ~v_724 | ~v_723 | ~v_722 | ~v_4588 | ~v_4584 | ~v_4580 | ~v_4576 | ~v_4572 | ~v_4568 | ~v_4564 | ~v_4560 | ~v_4556 | ~v_4552 | ~v_4548 | ~v_4544 | ~v_4540 | ~v_4536 | ~v_4532 | ~v_4528 | ~v_4512 | ~v_4508 | ~v_4504 | ~v_4500 | ~v_4496 | ~v_4492 | ~v_4488 | ~v_4484 | ~v_4480 | ~v_4476 | ~v_4472 | ~v_4468 | ~v_4464 | ~v_4460 | ~v_4456 | ~v_4452 | ~v_4436 | ~v_4432 | ~v_4428 | ~v_4424 | ~v_4420 | ~v_4416 | ~v_4412 | ~v_4408 | ~v_4404 | ~v_4400 | ~v_4396 | ~v_4392 | ~v_4388 | ~v_4384 | ~v_4380 | ~v_4376 | ~v_4360 | ~v_4356 | ~v_4352 | ~v_4348 | ~v_4344 | ~v_4340 | ~v_4336 | ~v_4332 | ~v_4328 | ~v_4324 | ~v_4320 | ~v_4316 | ~v_4312 | ~v_4308 | ~v_4304 | ~v_4300 | ~v_4284 | ~v_4123 | ~v_3962 | ~v_3801 | ~v_3640 | ~v_3275 | ~v_2910 | ~v_2749 | ~v_2588 | ~v_2217 | ~v_1850 | ~v_1269;
assign x_2 = v_4588 | ~v_4585;
assign x_3 = v_4588 | ~v_4586;
assign x_4 = v_4588 | ~v_4587;
assign x_5 = v_98 | v_103 | v_101 | v_97 | v_96 | v_100 | v_95 | v_94 | v_99 | v_93 | v_92 | v_102 | ~v_719 | ~v_718 | ~v_483 | ~v_717 | ~v_3021 | ~v_299 | ~v_2957 | ~v_3020 | ~v_2956 | ~v_2955 | ~v_482 | ~v_716 | ~v_3019 | ~v_298 | ~v_2954 | ~v_3018 | ~v_2953 | ~v_2952 | ~v_3386 | ~v_3320 | ~v_3385 | ~v_3319 | ~v_3318 | ~v_3384 | ~v_3317 | ~v_3383 | ~v_3316 | ~v_3315 | ~v_4526 | ~v_4525 | ~v_4524 | ~v_4523 | v_4587;
assign x_6 = v_54 | v_53 | v_56 | v_55 | v_61 | v_52 | v_50 | v_51 | v_60 | v_59 | v_58 | v_57 | ~v_714 | ~v_713 | ~v_3016 | ~v_3381 | ~v_3305 | ~v_3015 | ~v_266 | ~v_2942 | ~v_3380 | ~v_468 | ~v_712 | ~v_2941 | ~v_2940 | ~v_467 | ~v_711 | ~v_3014 | ~v_265 | ~v_2939 | ~v_3013 | ~v_2938 | ~v_2937 | ~v_3304 | ~v_3303 | ~v_3379 | ~v_3302 | ~v_3378 | ~v_3301 | ~v_3300 | ~v_4521 | ~v_4520 | ~v_4519 | ~v_4518 | v_4586;
assign x_7 = v_13 | v_9 | v_7 | v_18 | v_17 | v_16 | v_8 | v_15 | v_14 | v_12 | v_11 | v_10 | ~v_453 | ~v_709 | ~v_4516 | ~v_2927 | ~v_452 | ~v_708 | ~v_4515 | ~v_2926 | ~v_707 | ~v_706 | ~v_3292 | ~v_3011 | ~v_233 | ~v_2925 | ~v_3010 | ~v_2924 | ~v_3009 | ~v_232 | ~v_2923 | ~v_3008 | ~v_2922 | ~v_3376 | ~v_3289 | ~v_3375 | ~v_3288 | ~v_3374 | ~v_3287 | ~v_3373 | ~v_3286 | ~v_3285 | ~v_4514 | ~v_4513 | v_4585;
assign x_8 = v_4584 | ~v_4581;
assign x_9 = v_4584 | ~v_4582;
assign x_10 = v_4584 | ~v_4583;
assign x_11 = v_101 | v_97 | v_96 | v_100 | v_99 | v_92 | v_102 | v_172 | v_171 | v_170 | v_169 | v_147 | ~v_483 | ~v_3021 | ~v_3020 | ~v_2955 | ~v_482 | ~v_3019 | ~v_3018 | ~v_2952 | ~v_593 | ~v_592 | ~v_545 | ~v_3041 | ~v_3040 | ~v_591 | ~v_590 | ~v_544 | ~v_3039 | ~v_3038 | ~v_3386 | ~v_3385 | ~v_3318 | ~v_3384 | ~v_3383 | ~v_3315 | ~v_3406 | ~v_3405 | ~v_3404 | ~v_3403 | ~v_4526 | ~v_4525 | ~v_4524 | ~v_4523 | v_4583;
assign x_12 = v_54 | v_55 | v_50 | v_60 | v_59 | v_58 | v_57 | ~v_3016 | v_142 | v_168 | v_167 | v_166 | v_165 | ~v_3381 | ~v_3015 | ~v_3380 | ~v_468 | ~v_2940 | ~v_467 | ~v_3014 | ~v_3013 | ~v_2937 | ~v_588 | ~v_587 | ~v_530 | ~v_3036 | ~v_3035 | ~v_586 | ~v_585 | ~v_529 | ~v_3034 | ~v_3033 | ~v_3303 | ~v_3379 | ~v_3378 | ~v_3300 | ~v_3401 | ~v_3400 | ~v_3399 | ~v_3398 | ~v_4521 | ~v_4520 | ~v_4519 | ~v_4518 | v_4582;
assign x_13 = v_7 | v_17 | v_16 | v_15 | v_14 | v_12 | v_11 | ~v_453 | ~v_4516 | ~v_2927 | ~v_452 | ~v_4515 | ~v_2926 | v_134 | v_164 | v_163 | v_162 | v_161 | ~v_3011 | ~v_3010 | ~v_3009 | ~v_3008 | ~v_583 | ~v_582 | ~v_515 | ~v_3031 | ~v_3030 | ~v_581 | ~v_580 | ~v_514 | ~v_3029 | ~v_3028 | ~v_3376 | ~v_3375 | ~v_3288 | ~v_3374 | ~v_3373 | ~v_3285 | ~v_3396 | ~v_3395 | ~v_3394 | ~v_3393 | ~v_4514 | ~v_4513 | v_4581;
assign x_14 = v_4580 | ~v_4577;
assign x_15 = v_4580 | ~v_4578;
assign x_16 = v_4580 | ~v_4579;
assign x_17 = v_103 | v_101 | v_100 | v_95 | v_92 | v_102 | v_171 | v_170 | v_169 | v_150 | v_149 | v_148 | ~v_2955 | ~v_2952 | ~v_545 | ~v_3041 | ~v_3040 | ~v_544 | ~v_3039 | ~v_3038 | ~v_561 | ~v_560 | ~v_559 | ~v_558 | ~v_387 | ~v_2989 | ~v_2988 | ~v_386 | ~v_2987 | ~v_2986 | ~v_3318 | ~v_3315 | ~v_3406 | ~v_3405 | ~v_3404 | ~v_3403 | ~v_3354 | ~v_3353 | ~v_3352 | ~v_3351 | ~v_4526 | ~v_4525 | ~v_4524 | ~v_4523 | v_4579;
assign x_18 = v_53 | v_61 | v_50 | v_60 | v_59 | v_58 | v_144 | v_145 | v_143 | v_167 | v_166 | v_165 | ~v_2940 | ~v_2937 | ~v_530 | ~v_3036 | ~v_3035 | ~v_529 | ~v_3034 | ~v_3033 | ~v_556 | ~v_555 | ~v_554 | ~v_553 | ~v_372 | ~v_2984 | ~v_2983 | ~v_371 | ~v_2982 | ~v_2981 | ~v_3303 | ~v_3300 | ~v_3401 | ~v_3400 | ~v_3399 | ~v_3398 | ~v_3349 | ~v_3348 | ~v_3347 | ~v_3346 | ~v_4521 | ~v_4520 | ~v_4519 | ~v_4518 | v_4578;
assign x_19 = v_7 | v_18 | v_17 | v_16 | v_15 | v_10 | ~v_4516 | ~v_2927 | ~v_4515 | ~v_2926 | v_136 | v_135 | v_137 | v_163 | v_162 | v_161 | ~v_515 | ~v_3031 | ~v_3030 | ~v_514 | ~v_3029 | ~v_3028 | ~v_551 | ~v_550 | ~v_549 | ~v_548 | ~v_357 | ~v_2979 | ~v_2978 | ~v_356 | ~v_2977 | ~v_2976 | ~v_3288 | ~v_3285 | ~v_3396 | ~v_3395 | ~v_3394 | ~v_3393 | ~v_3344 | ~v_3343 | ~v_3342 | ~v_3341 | ~v_4514 | ~v_4513 | v_4577;
assign x_20 = v_4576 | ~v_4573;
assign x_21 = v_4576 | ~v_4574;
assign x_22 = v_4576 | ~v_4575;
assign x_23 = v_98 | v_103 | v_101 | v_100 | v_94 | v_93 | v_92 | v_151 | v_150 | v_149 | v_148 | v_147 | ~v_299 | ~v_2957 | ~v_2956 | ~v_2955 | ~v_298 | ~v_2954 | ~v_2953 | ~v_2952 | ~v_387 | ~v_2989 | ~v_2988 | ~v_386 | ~v_2987 | ~v_2986 | ~v_499 | ~v_498 | ~v_497 | ~v_496 | ~v_3320 | ~v_3319 | ~v_3318 | ~v_3317 | ~v_3316 | ~v_3315 | ~v_3354 | ~v_3353 | ~v_3352 | ~v_3351 | ~v_4526 | ~v_4525 | ~v_4524 | ~v_4523 | v_4575;
assign x_24 = v_56 | v_61 | v_52 | v_50 | v_51 | v_59 | v_58 | v_144 | v_145 | v_143 | v_142 | v_146 | ~v_3305 | ~v_266 | ~v_2942 | ~v_2941 | ~v_2940 | ~v_265 | ~v_2939 | ~v_2938 | ~v_2937 | ~v_372 | ~v_2984 | ~v_2983 | ~v_371 | ~v_2982 | ~v_2981 | ~v_494 | ~v_493 | ~v_492 | ~v_491 | ~v_3304 | ~v_3303 | ~v_3302 | ~v_3301 | ~v_3300 | ~v_3349 | ~v_3348 | ~v_3347 | ~v_3346 | ~v_4521 | ~v_4520 | ~v_4519 | ~v_4518 | v_4574;
assign x_25 = v_13 | v_9 | v_7 | v_18 | v_16 | v_8 | v_15 | ~v_4516 | ~v_2927 | ~v_4515 | ~v_2926 | v_136 | v_135 | v_134 | ~v_3292 | v_137 | v_138 | ~v_233 | ~v_2925 | ~v_2924 | ~v_232 | ~v_2923 | ~v_2922 | ~v_357 | ~v_2979 | ~v_2978 | ~v_356 | ~v_2977 | ~v_2976 | ~v_489 | ~v_488 | ~v_487 | ~v_486 | ~v_3289 | ~v_3288 | ~v_3287 | ~v_3286 | ~v_3285 | ~v_3344 | ~v_3343 | ~v_3342 | ~v_3341 | ~v_4514 | ~v_4513 | v_4573;
assign x_26 = v_4572 | ~v_4569;
assign x_27 = v_4572 | ~v_4570;
assign x_28 = v_4572 | ~v_4571;
assign x_29 = v_103 | v_101 | v_97 | v_96 | v_100 | v_99 | v_92 | v_102 | v_171 | v_170 | v_169 | v_147 | ~v_703 | ~v_702 | ~v_483 | ~v_3021 | ~v_3020 | ~v_2955 | ~v_482 | ~v_3019 | ~v_3018 | ~v_2952 | ~v_701 | ~v_653 | ~v_2973 | ~v_2972 | ~v_700 | ~v_652 | ~v_2971 | ~v_2970 | ~v_3386 | ~v_3385 | ~v_3318 | ~v_3384 | ~v_3383 | ~v_3315 | ~v_3338 | ~v_3337 | ~v_3336 | ~v_3335 | ~v_4526 | ~v_4525 | ~v_4524 | ~v_4523 | v_4571;
assign x_30 = v_54 | v_55 | v_61 | v_50 | v_60 | v_59 | v_58 | v_57 | ~v_3016 | v_142 | v_167 | v_166 | v_165 | ~v_698 | ~v_697 | ~v_3381 | ~v_3015 | ~v_3380 | ~v_468 | ~v_2940 | ~v_467 | ~v_3014 | ~v_3013 | ~v_2937 | ~v_696 | ~v_638 | ~v_2968 | ~v_2967 | ~v_695 | ~v_637 | ~v_2966 | ~v_2965 | ~v_3303 | ~v_3379 | ~v_3378 | ~v_3300 | ~v_3333 | ~v_3332 | ~v_3331 | ~v_3330 | ~v_4521 | ~v_4520 | ~v_4519 | ~v_4518 | v_4570;
assign x_31 = v_7 | v_18 | v_17 | v_16 | v_15 | v_14 | v_12 | v_11 | ~v_453 | ~v_4516 | ~v_2927 | ~v_452 | ~v_4515 | ~v_2926 | v_134 | v_163 | v_162 | v_161 | ~v_693 | ~v_692 | ~v_3011 | ~v_3010 | ~v_3009 | ~v_3008 | ~v_691 | ~v_623 | ~v_2963 | ~v_2962 | ~v_690 | ~v_622 | ~v_2961 | ~v_2960 | ~v_3376 | ~v_3375 | ~v_3288 | ~v_3374 | ~v_3373 | ~v_3285 | ~v_3328 | ~v_3327 | ~v_3326 | ~v_3325 | ~v_4514 | ~v_4513 | v_4569;
assign x_32 = v_4568 | ~v_4565;
assign x_33 = v_4568 | ~v_4566;
assign x_34 = v_4568 | ~v_4567;
assign x_35 = v_103 | v_101 | v_100 | v_95 | v_92 | v_102 | v_171 | v_170 | v_169 | v_150 | v_149 | v_148 | ~v_3322 | ~v_3321 | ~v_2955 | ~v_2952 | ~v_435 | ~v_2951 | ~v_2950 | ~v_434 | ~v_2949 | ~v_2948 | ~v_653 | ~v_2973 | ~v_2972 | ~v_652 | ~v_2971 | ~v_2970 | ~v_687 | ~v_686 | ~v_685 | ~v_684 | ~v_3318 | ~v_3315 | ~v_3314 | ~v_3313 | ~v_3338 | ~v_3337 | ~v_3336 | ~v_3335 | ~v_4526 | ~v_4525 | ~v_4524 | ~v_4523 | v_4567;
assign x_36 = v_53 | v_61 | v_50 | v_60 | v_59 | v_58 | v_144 | v_145 | v_143 | v_167 | v_166 | v_165 | ~v_3307 | ~v_3306 | ~v_2940 | ~v_2937 | ~v_420 | ~v_2936 | ~v_2935 | ~v_419 | ~v_2934 | ~v_2933 | ~v_638 | ~v_2968 | ~v_2967 | ~v_637 | ~v_2966 | ~v_2965 | ~v_682 | ~v_681 | ~v_680 | ~v_679 | ~v_3303 | ~v_3300 | ~v_3299 | ~v_3298 | ~v_3333 | ~v_3332 | ~v_3331 | ~v_3330 | ~v_4521 | ~v_4520 | ~v_4519 | ~v_4518 | v_4566;
assign x_37 = v_7 | v_18 | v_17 | v_16 | v_15 | v_10 | ~v_4516 | ~v_2927 | ~v_4515 | ~v_2926 | v_136 | v_135 | v_137 | v_163 | v_162 | v_161 | ~v_3291 | ~v_3290 | ~v_405 | ~v_2921 | ~v_2920 | ~v_404 | ~v_2919 | ~v_2918 | ~v_623 | ~v_2963 | ~v_2962 | ~v_622 | ~v_2961 | ~v_2960 | ~v_677 | ~v_676 | ~v_675 | ~v_674 | ~v_3288 | ~v_3285 | ~v_3284 | ~v_3283 | ~v_3328 | ~v_3327 | ~v_3326 | ~v_3325 | ~v_4514 | ~v_4513 | v_4565;
assign x_38 = v_4564 | ~v_4561;
assign x_39 = v_4564 | ~v_4562;
assign x_40 = v_4564 | ~v_4563;
assign x_41 = v_98 | v_103 | v_101 | v_100 | v_94 | v_93 | v_92 | v_102 | v_150 | v_149 | v_148 | v_147 | ~v_609 | ~v_608 | ~v_3322 | ~v_3321 | ~v_299 | ~v_2957 | ~v_2956 | ~v_2955 | ~v_298 | ~v_2954 | ~v_2953 | ~v_2952 | ~v_435 | ~v_2951 | ~v_2950 | ~v_434 | ~v_2949 | ~v_2948 | ~v_607 | ~v_606 | ~v_3320 | ~v_3319 | ~v_3318 | ~v_3317 | ~v_3316 | ~v_3315 | ~v_3314 | ~v_3313 | ~v_4526 | ~v_4525 | ~v_4524 | ~v_4523 | v_4563;
assign x_42 = v_56 | v_61 | v_52 | v_50 | v_51 | v_60 | v_59 | v_58 | v_144 | v_145 | v_143 | v_142 | ~v_604 | ~v_603 | ~v_3307 | ~v_3306 | ~v_3305 | ~v_266 | ~v_2942 | ~v_2941 | ~v_2940 | ~v_265 | ~v_2939 | ~v_2938 | ~v_2937 | ~v_420 | ~v_2936 | ~v_2935 | ~v_419 | ~v_2934 | ~v_2933 | ~v_602 | ~v_601 | ~v_3304 | ~v_3303 | ~v_3302 | ~v_3301 | ~v_3300 | ~v_3299 | ~v_3298 | ~v_4521 | ~v_4520 | ~v_4519 | ~v_4518 | v_4562;
assign x_43 = v_13 | v_9 | v_7 | v_18 | v_17 | v_16 | v_8 | v_15 | ~v_4516 | ~v_2927 | ~v_4515 | ~v_2926 | v_136 | v_135 | v_134 | ~v_3292 | v_137 | ~v_599 | ~v_598 | ~v_3291 | ~v_3290 | ~v_233 | ~v_2925 | ~v_2924 | ~v_232 | ~v_2923 | ~v_2922 | ~v_405 | ~v_2921 | ~v_2920 | ~v_404 | ~v_2919 | ~v_2918 | ~v_597 | ~v_596 | ~v_3289 | ~v_3288 | ~v_3287 | ~v_3286 | ~v_3285 | ~v_3284 | ~v_3283 | ~v_4514 | ~v_4513 | v_4561;
assign x_44 = v_4560 | ~v_4557;
assign x_45 = v_4560 | ~v_4558;
assign x_46 = v_4560 | ~v_4559;
assign x_47 = v_103 | v_101 | v_97 | v_96 | v_99 | v_92 | v_102 | v_171 | v_170 | v_169 | v_147 | v_181 | ~v_483 | ~v_3021 | ~v_3020 | ~v_2955 | ~v_482 | ~v_3019 | ~v_3018 | ~v_2952 | ~v_481 | ~v_480 | ~v_345 | ~v_3073 | ~v_3072 | ~v_479 | ~v_478 | ~v_344 | ~v_3071 | ~v_3070 | ~v_3386 | ~v_3385 | ~v_3318 | ~v_3384 | ~v_3383 | ~v_3315 | ~v_3438 | ~v_3437 | ~v_3436 | ~v_3435 | ~v_4526 | ~v_4525 | ~v_4524 | ~v_4523 | v_4559;
assign x_48 = v_54 | v_55 | v_61 | v_50 | v_60 | v_59 | v_57 | ~v_3016 | v_180 | v_142 | v_167 | v_166 | v_165 | ~v_3381 | ~v_3015 | ~v_3380 | ~v_468 | ~v_2940 | ~v_467 | ~v_3014 | ~v_3013 | ~v_2937 | ~v_466 | ~v_465 | ~v_330 | ~v_3068 | ~v_3067 | ~v_464 | ~v_463 | ~v_329 | ~v_3066 | ~v_3065 | ~v_3303 | ~v_3379 | ~v_3378 | ~v_3300 | ~v_3433 | ~v_3432 | ~v_3431 | ~v_3430 | ~v_4521 | ~v_4520 | ~v_4519 | ~v_4518 | v_4558;
assign x_49 = v_7 | v_18 | v_17 | v_16 | v_14 | v_12 | v_11 | ~v_453 | ~v_4516 | ~v_2927 | ~v_452 | ~v_4515 | ~v_2926 | v_134 | v_179 | v_163 | v_162 | v_161 | ~v_3011 | ~v_3010 | ~v_3009 | ~v_3008 | ~v_451 | ~v_450 | ~v_315 | ~v_3063 | ~v_3062 | ~v_449 | ~v_448 | ~v_314 | ~v_3061 | ~v_3060 | ~v_3376 | ~v_3375 | ~v_3288 | ~v_3374 | ~v_3373 | ~v_3285 | ~v_3428 | ~v_3427 | ~v_3426 | ~v_3425 | ~v_4514 | ~v_4513 | v_4557;
assign x_50 = v_4556 | ~v_4553;
assign x_51 = v_4556 | ~v_4554;
assign x_52 = v_4556 | ~v_4555;
assign x_53 = v_103 | v_95 | v_92 | v_102 | v_171 | v_170 | v_169 | v_160 | v_150 | v_149 | v_148 | v_181 | ~v_2955 | ~v_2952 | ~v_297 | ~v_3005 | ~v_3004 | ~v_296 | ~v_3003 | ~v_3002 | ~v_345 | ~v_3073 | ~v_3072 | ~v_344 | ~v_3071 | ~v_3070 | ~v_343 | ~v_342 | ~v_341 | ~v_340 | ~v_3318 | ~v_3315 | ~v_3370 | ~v_3369 | ~v_3368 | ~v_3367 | ~v_3438 | ~v_3437 | ~v_3436 | ~v_3435 | ~v_4526 | ~v_4525 | ~v_4524 | ~v_4523 | v_4555;
assign x_54 = v_53 | v_61 | v_50 | v_60 | v_144 | v_180 | v_159 | v_145 | v_143 | v_167 | v_166 | v_165 | ~v_2940 | ~v_2937 | ~v_264 | ~v_3000 | ~v_2999 | ~v_263 | ~v_2998 | ~v_2997 | ~v_330 | ~v_3068 | ~v_3067 | ~v_329 | ~v_3066 | ~v_3065 | ~v_328 | ~v_327 | ~v_326 | ~v_325 | ~v_3303 | ~v_3300 | ~v_3365 | ~v_3364 | ~v_3363 | ~v_3362 | ~v_3433 | ~v_3432 | ~v_3431 | ~v_3430 | ~v_4521 | ~v_4520 | ~v_4519 | ~v_4518 | v_4554;
assign x_55 = v_7 | v_18 | v_17 | v_10 | ~v_4516 | ~v_2927 | ~v_4515 | ~v_2926 | v_136 | v_135 | v_137 | v_179 | v_163 | v_162 | v_161 | v_155 | ~v_231 | ~v_2995 | ~v_2994 | ~v_230 | ~v_2993 | ~v_2992 | ~v_315 | ~v_3063 | ~v_3062 | ~v_314 | ~v_3061 | ~v_3060 | ~v_313 | ~v_312 | ~v_311 | ~v_310 | ~v_3288 | ~v_3285 | ~v_3360 | ~v_3359 | ~v_3358 | ~v_3357 | ~v_3428 | ~v_3427 | ~v_3426 | ~v_3425 | ~v_4514 | ~v_4513 | v_4553;
assign x_56 = v_4552 | ~v_4549;
assign x_57 = v_4552 | ~v_4550;
assign x_58 = v_4552 | ~v_4551;
assign x_59 = v_98 | v_103 | v_100 | v_94 | v_93 | v_92 | v_102 | v_160 | v_150 | v_149 | v_148 | v_147 | ~v_299 | ~v_2957 | ~v_2956 | ~v_2955 | ~v_298 | ~v_2954 | ~v_2953 | ~v_2952 | ~v_297 | ~v_3005 | ~v_3004 | ~v_296 | ~v_3003 | ~v_3002 | ~v_295 | ~v_294 | ~v_293 | ~v_292 | ~v_3320 | ~v_3319 | ~v_3318 | ~v_3317 | ~v_3316 | ~v_3315 | ~v_3370 | ~v_3369 | ~v_3368 | ~v_3367 | ~v_4526 | ~v_4525 | ~v_4524 | ~v_4523 | v_4551;
assign x_60 = v_56 | v_61 | v_52 | v_50 | v_51 | v_60 | v_58 | v_144 | v_159 | v_145 | v_143 | v_142 | ~v_3305 | ~v_266 | ~v_2942 | ~v_2941 | ~v_2940 | ~v_265 | ~v_2939 | ~v_2938 | ~v_2937 | ~v_264 | ~v_3000 | ~v_2999 | ~v_263 | ~v_2998 | ~v_2997 | ~v_262 | ~v_261 | ~v_260 | ~v_259 | ~v_3304 | ~v_3303 | ~v_3302 | ~v_3301 | ~v_3300 | ~v_3365 | ~v_3364 | ~v_3363 | ~v_3362 | ~v_4521 | ~v_4520 | ~v_4519 | ~v_4518 | v_4550;
assign x_61 = v_13 | v_9 | v_7 | v_18 | v_17 | v_8 | v_15 | ~v_4516 | ~v_2927 | ~v_4515 | ~v_2926 | v_136 | v_135 | v_134 | ~v_3292 | v_137 | v_155 | ~v_233 | ~v_2925 | ~v_2924 | ~v_232 | ~v_2923 | ~v_2922 | ~v_231 | ~v_2995 | ~v_2994 | ~v_230 | ~v_2993 | ~v_2992 | ~v_229 | ~v_228 | ~v_227 | ~v_226 | ~v_3289 | ~v_3288 | ~v_3287 | ~v_3286 | ~v_3285 | ~v_3360 | ~v_3359 | ~v_3358 | ~v_3357 | ~v_4514 | ~v_4513 | v_4549;
assign x_62 = v_4548 | ~v_4545;
assign x_63 = v_4548 | ~v_4546;
assign x_64 = v_4548 | ~v_4547;
assign x_65 = v_103 | v_101 | v_100 | v_92 | v_151 | v_171 | v_170 | v_169 | v_150 | v_149 | v_148 | v_147 | ~v_3322 | ~v_3321 | ~v_577 | ~v_576 | ~v_2955 | ~v_2952 | ~v_545 | ~v_3041 | ~v_3040 | ~v_544 | ~v_3039 | ~v_3038 | ~v_575 | ~v_574 | ~v_435 | ~v_2951 | ~v_2950 | ~v_434 | ~v_2949 | ~v_2948 | ~v_3318 | ~v_3315 | ~v_3406 | ~v_3405 | ~v_3404 | ~v_3403 | ~v_3314 | ~v_3313 | ~v_4526 | ~v_4525 | ~v_4524 | ~v_4523 | v_4547;
assign x_66 = v_61 | v_50 | v_59 | v_58 | v_144 | v_145 | v_143 | v_142 | v_167 | v_166 | v_165 | v_146 | ~v_3307 | ~v_3306 | ~v_572 | ~v_571 | ~v_2940 | ~v_2937 | ~v_530 | ~v_3036 | ~v_3035 | ~v_529 | ~v_3034 | ~v_3033 | ~v_570 | ~v_569 | ~v_420 | ~v_2936 | ~v_2935 | ~v_419 | ~v_2934 | ~v_2933 | ~v_3303 | ~v_3300 | ~v_3401 | ~v_3400 | ~v_3399 | ~v_3398 | ~v_3299 | ~v_3298 | ~v_4521 | ~v_4520 | ~v_4519 | ~v_4518 | v_4546;
assign x_67 = v_7 | v_18 | v_16 | v_15 | ~v_4516 | ~v_2927 | ~v_4515 | ~v_2926 | v_136 | v_135 | v_134 | v_137 | v_138 | v_163 | v_162 | v_161 | ~v_3291 | ~v_3290 | ~v_567 | ~v_566 | ~v_515 | ~v_3031 | ~v_3030 | ~v_514 | ~v_3029 | ~v_3028 | ~v_565 | ~v_564 | ~v_405 | ~v_2921 | ~v_2920 | ~v_404 | ~v_2919 | ~v_2918 | ~v_3288 | ~v_3285 | ~v_3396 | ~v_3395 | ~v_3394 | ~v_3393 | ~v_3284 | ~v_3283 | ~v_4514 | ~v_4513 | v_4545;
assign x_68 = v_4544 | ~v_4541;
assign x_69 = v_4544 | ~v_4542;
assign x_70 = v_4544 | ~v_4543;
assign x_71 = v_101 | v_100 | v_92 | v_102 | v_172 | v_171 | v_170 | v_169 | v_150 | v_149 | v_148 | v_147 | ~v_671 | ~v_670 | ~v_2955 | ~v_2952 | ~v_387 | ~v_2989 | ~v_2988 | ~v_386 | ~v_2987 | ~v_2986 | ~v_653 | ~v_2973 | ~v_2972 | ~v_652 | ~v_2971 | ~v_2970 | ~v_669 | ~v_668 | ~v_3318 | ~v_3315 | ~v_3354 | ~v_3353 | ~v_3352 | ~v_3351 | ~v_3338 | ~v_3337 | ~v_3336 | ~v_3335 | ~v_4526 | ~v_4525 | ~v_4524 | ~v_4523 | v_4543;
assign x_72 = v_50 | v_60 | v_59 | v_58 | v_144 | v_145 | v_143 | v_142 | v_168 | v_167 | v_166 | v_165 | ~v_666 | ~v_665 | ~v_2940 | ~v_2937 | ~v_372 | ~v_2984 | ~v_2983 | ~v_371 | ~v_2982 | ~v_2981 | ~v_638 | ~v_2968 | ~v_2967 | ~v_637 | ~v_2966 | ~v_2965 | ~v_664 | ~v_663 | ~v_3303 | ~v_3300 | ~v_3349 | ~v_3348 | ~v_3347 | ~v_3346 | ~v_3333 | ~v_3332 | ~v_3331 | ~v_3330 | ~v_4521 | ~v_4520 | ~v_4519 | ~v_4518 | v_4542;
assign x_73 = v_7 | v_17 | v_16 | v_15 | ~v_4516 | ~v_2927 | ~v_4515 | ~v_2926 | v_136 | v_135 | v_134 | v_137 | v_164 | v_163 | v_162 | v_161 | ~v_661 | ~v_660 | ~v_357 | ~v_2979 | ~v_2978 | ~v_356 | ~v_2977 | ~v_2976 | ~v_623 | ~v_2963 | ~v_2962 | ~v_622 | ~v_2961 | ~v_2960 | ~v_659 | ~v_658 | ~v_3288 | ~v_3285 | ~v_3344 | ~v_3343 | ~v_3342 | ~v_3341 | ~v_3328 | ~v_3327 | ~v_3326 | ~v_3325 | ~v_4514 | ~v_4513 | v_4541;
assign x_74 = v_4540 | ~v_4537;
assign x_75 = v_4540 | ~v_4538;
assign x_76 = v_4540 | ~v_4539;
assign x_77 = v_103 | v_101 | v_92 | v_102 | v_171 | v_170 | v_169 | v_150 | v_149 | v_148 | v_147 | v_181 | ~v_391 | ~v_390 | ~v_2955 | ~v_2952 | ~v_387 | ~v_2989 | ~v_2988 | ~v_386 | ~v_2987 | ~v_2986 | ~v_345 | ~v_3073 | ~v_3072 | ~v_344 | ~v_3071 | ~v_3070 | ~v_385 | ~v_384 | ~v_3318 | ~v_3315 | ~v_3354 | ~v_3353 | ~v_3352 | ~v_3351 | ~v_3438 | ~v_3437 | ~v_3436 | ~v_3435 | ~v_4526 | ~v_4525 | ~v_4524 | ~v_4523 | v_4539;
assign x_78 = v_61 | v_50 | v_60 | v_59 | v_144 | v_180 | v_145 | v_143 | v_142 | v_167 | v_166 | v_165 | ~v_376 | ~v_375 | ~v_2940 | ~v_2937 | ~v_372 | ~v_2984 | ~v_2983 | ~v_371 | ~v_2982 | ~v_2981 | ~v_330 | ~v_3068 | ~v_3067 | ~v_329 | ~v_3066 | ~v_3065 | ~v_370 | ~v_369 | ~v_3303 | ~v_3300 | ~v_3349 | ~v_3348 | ~v_3347 | ~v_3346 | ~v_3433 | ~v_3432 | ~v_3431 | ~v_3430 | ~v_4521 | ~v_4520 | ~v_4519 | ~v_4518 | v_4538;
assign x_79 = v_7 | v_18 | v_17 | v_16 | ~v_4516 | ~v_2927 | ~v_4515 | ~v_2926 | v_136 | v_135 | v_134 | v_137 | v_179 | v_163 | v_162 | v_161 | ~v_361 | ~v_360 | ~v_357 | ~v_2979 | ~v_2978 | ~v_356 | ~v_2977 | ~v_2976 | ~v_315 | ~v_3063 | ~v_3062 | ~v_314 | ~v_3061 | ~v_3060 | ~v_355 | ~v_354 | ~v_3288 | ~v_3285 | ~v_3344 | ~v_3343 | ~v_3342 | ~v_3341 | ~v_3428 | ~v_3427 | ~v_3426 | ~v_3425 | ~v_4514 | ~v_4513 | v_4537;
assign x_80 = v_4536 | ~v_4533;
assign x_81 = v_4536 | ~v_4534;
assign x_82 = v_4536 | ~v_4535;
assign x_83 = v_103 | v_100 | v_92 | v_102 | v_171 | v_170 | v_169 | v_160 | v_150 | v_149 | v_148 | v_147 | ~v_2955 | ~v_2952 | ~v_545 | ~v_3041 | ~v_3040 | ~v_544 | ~v_3039 | ~v_3038 | ~v_543 | ~v_542 | ~v_541 | ~v_540 | ~v_297 | ~v_3005 | ~v_3004 | ~v_296 | ~v_3003 | ~v_3002 | ~v_3318 | ~v_3315 | ~v_3406 | ~v_3405 | ~v_3404 | ~v_3403 | ~v_3370 | ~v_3369 | ~v_3368 | ~v_3367 | ~v_4526 | ~v_4525 | ~v_4524 | ~v_4523 | v_4535;
assign x_84 = v_61 | v_50 | v_60 | v_58 | v_144 | v_159 | v_145 | v_143 | v_142 | v_167 | v_166 | v_165 | ~v_2940 | ~v_2937 | ~v_530 | ~v_3036 | ~v_3035 | ~v_529 | ~v_3034 | ~v_3033 | ~v_528 | ~v_527 | ~v_526 | ~v_525 | ~v_264 | ~v_3000 | ~v_2999 | ~v_263 | ~v_2998 | ~v_2997 | ~v_3303 | ~v_3300 | ~v_3401 | ~v_3400 | ~v_3399 | ~v_3398 | ~v_3365 | ~v_3364 | ~v_3363 | ~v_3362 | ~v_4521 | ~v_4520 | ~v_4519 | ~v_4518 | v_4534;
assign x_85 = v_7 | v_18 | v_17 | v_15 | ~v_4516 | ~v_2927 | ~v_4515 | ~v_2926 | v_136 | v_135 | v_134 | v_137 | v_163 | v_162 | v_161 | v_155 | ~v_515 | ~v_3031 | ~v_3030 | ~v_514 | ~v_3029 | ~v_3028 | ~v_513 | ~v_512 | ~v_511 | ~v_510 | ~v_231 | ~v_2995 | ~v_2994 | ~v_230 | ~v_2993 | ~v_2992 | ~v_3288 | ~v_3285 | ~v_3396 | ~v_3395 | ~v_3394 | ~v_3393 | ~v_3360 | ~v_3359 | ~v_3358 | ~v_3357 | ~v_4514 | ~v_4513 | v_4533;
assign x_86 = v_4532 | ~v_4529;
assign x_87 = v_4532 | ~v_4530;
assign x_88 = v_4532 | ~v_4531;
assign x_89 = v_103 | v_100 | v_92 | v_151 | v_171 | v_170 | v_169 | v_160 | v_150 | v_149 | v_148 | v_147 | ~v_655 | ~v_654 | ~v_2955 | ~v_2952 | ~v_297 | ~v_3005 | ~v_3004 | ~v_296 | ~v_3003 | ~v_3002 | ~v_653 | ~v_2973 | ~v_2972 | ~v_652 | ~v_2971 | ~v_2970 | ~v_651 | ~v_650 | ~v_3318 | ~v_3315 | ~v_3370 | ~v_3369 | ~v_3368 | ~v_3367 | ~v_3338 | ~v_3337 | ~v_3336 | ~v_3335 | ~v_4526 | ~v_4525 | ~v_4524 | ~v_4523 | v_4531;
assign x_90 = v_61 | v_50 | v_58 | v_144 | v_159 | v_145 | v_143 | v_142 | v_167 | v_166 | v_165 | v_146 | ~v_640 | ~v_639 | ~v_2940 | ~v_2937 | ~v_264 | ~v_3000 | ~v_2999 | ~v_263 | ~v_2998 | ~v_2997 | ~v_638 | ~v_2968 | ~v_2967 | ~v_637 | ~v_2966 | ~v_2965 | ~v_636 | ~v_635 | ~v_3303 | ~v_3300 | ~v_3365 | ~v_3364 | ~v_3363 | ~v_3362 | ~v_3333 | ~v_3332 | ~v_3331 | ~v_3330 | ~v_4521 | ~v_4520 | ~v_4519 | ~v_4518 | v_4530;
assign x_91 = v_7 | v_18 | v_15 | ~v_4516 | ~v_2927 | ~v_4515 | ~v_2926 | v_136 | v_135 | v_134 | v_137 | v_138 | v_163 | v_162 | v_161 | v_155 | ~v_625 | ~v_624 | ~v_231 | ~v_2995 | ~v_2994 | ~v_230 | ~v_2993 | ~v_2992 | ~v_623 | ~v_2963 | ~v_2962 | ~v_622 | ~v_2961 | ~v_2960 | ~v_621 | ~v_620 | ~v_3288 | ~v_3285 | ~v_3360 | ~v_3359 | ~v_3358 | ~v_3357 | ~v_3328 | ~v_3327 | ~v_3326 | ~v_3325 | ~v_4514 | ~v_4513 | v_4529;
assign x_92 = v_4528 | ~v_4517;
assign x_93 = v_4528 | ~v_4522;
assign x_94 = v_4528 | ~v_4527;
assign x_95 = v_101 | v_92 | v_102 | v_172 | v_171 | v_170 | v_169 | v_150 | v_149 | v_148 | v_147 | v_181 | ~v_3322 | ~v_3321 | ~v_437 | ~v_436 | ~v_2955 | ~v_2952 | ~v_435 | ~v_2951 | ~v_2950 | ~v_434 | ~v_2949 | ~v_2948 | ~v_345 | ~v_3073 | ~v_3072 | ~v_344 | ~v_3071 | ~v_3070 | ~v_433 | ~v_432 | ~v_3318 | ~v_3315 | ~v_3314 | ~v_3313 | ~v_3438 | ~v_3437 | ~v_3436 | ~v_3435 | ~v_4526 | ~v_4525 | ~v_4524 | ~v_4523 | v_4527;
assign x_96 = v_4526 | v_123;
assign x_97 = v_4526 | v_19;
assign x_98 = v_4525 | v_120;
assign x_99 = v_4525 | v_19;
assign x_100 = v_4524 | v_108;
assign x_101 = v_4524 | ~v_19;
assign x_102 = v_4523 | v_105;
assign x_103 = v_4523 | ~v_19;
assign x_104 = v_50 | v_60 | v_59 | v_144 | v_180 | v_145 | v_143 | v_142 | v_168 | v_167 | v_166 | v_165 | ~v_3307 | ~v_3306 | ~v_422 | ~v_421 | ~v_2940 | ~v_2937 | ~v_420 | ~v_2936 | ~v_2935 | ~v_419 | ~v_2934 | ~v_2933 | ~v_330 | ~v_3068 | ~v_3067 | ~v_329 | ~v_3066 | ~v_3065 | ~v_418 | ~v_417 | ~v_3303 | ~v_3300 | ~v_3299 | ~v_3298 | ~v_3433 | ~v_3432 | ~v_3431 | ~v_3430 | ~v_4521 | ~v_4520 | ~v_4519 | ~v_4518 | v_4522;
assign x_105 = v_4521 | v_81;
assign x_106 = v_4521 | v_19;
assign x_107 = v_4520 | v_78;
assign x_108 = v_4520 | v_19;
assign x_109 = v_4519 | v_66;
assign x_110 = v_4519 | ~v_19;
assign x_111 = v_4518 | v_63;
assign x_112 = v_4518 | ~v_19;
assign x_113 = v_7 | v_17 | v_16 | ~v_4516 | ~v_2927 | ~v_4515 | ~v_2926 | v_136 | v_135 | v_134 | v_137 | v_179 | v_164 | v_163 | v_162 | v_161 | ~v_3291 | ~v_3290 | ~v_407 | ~v_406 | ~v_405 | ~v_2921 | ~v_2920 | ~v_404 | ~v_2919 | ~v_2918 | ~v_315 | ~v_3063 | ~v_3062 | ~v_314 | ~v_3061 | ~v_3060 | ~v_403 | ~v_402 | ~v_3288 | ~v_3285 | ~v_3284 | ~v_3283 | ~v_3428 | ~v_3427 | ~v_3426 | ~v_3425 | ~v_4514 | ~v_4513 | v_4517;
assign x_114 = v_4516 | v_36;
assign x_115 = v_4516 | v_19;
assign x_116 = v_4515 | v_21;
assign x_117 = v_4515 | ~v_19;
assign x_118 = v_4514 | v_39;
assign x_119 = v_4514 | v_19;
assign x_120 = v_4513 | v_24;
assign x_121 = v_4513 | ~v_19;
assign x_122 = v_4512 | ~v_4509;
assign x_123 = v_4512 | ~v_4510;
assign x_124 = v_4512 | ~v_4511;
assign x_125 = v_98 | v_103 | v_101 | v_100 | v_95 | v_99 | v_92 | v_102 | ~v_719 | ~v_718 | v_170 | v_169 | v_149 | v_148 | ~v_2331 | ~v_2267 | ~v_2330 | ~v_2266 | ~v_2265 | ~v_2329 | ~v_2264 | ~v_2328 | ~v_2263 | ~v_2262 | ~v_483 | ~v_717 | ~v_299 | ~v_482 | ~v_716 | ~v_298 | ~v_1962 | ~v_1898 | ~v_1961 | ~v_1897 | ~v_1896 | ~v_1960 | ~v_1895 | ~v_1959 | ~v_1894 | ~v_1893 | ~v_4450 | ~v_4449 | ~v_4448 | ~v_4447 | v_4511;
assign x_126 = v_53 | v_56 | v_61 | v_50 | v_60 | v_59 | v_58 | v_57 | ~v_714 | ~v_713 | v_144 | v_143 | v_166 | v_165 | ~v_266 | ~v_2326 | ~v_2252 | ~v_2325 | ~v_2251 | ~v_2250 | ~v_2324 | ~v_2249 | ~v_2323 | ~v_2248 | ~v_2247 | ~v_468 | ~v_712 | ~v_467 | ~v_711 | ~v_265 | ~v_1957 | ~v_1883 | ~v_1956 | ~v_1882 | ~v_1881 | ~v_1955 | ~v_1880 | ~v_1954 | ~v_1879 | ~v_1878 | ~v_4445 | ~v_4444 | ~v_4443 | ~v_4442 | v_4510;
assign x_127 = v_13 | v_7 | v_18 | v_17 | v_16 | v_15 | v_14 | v_10 | ~v_453 | ~v_709 | ~v_452 | ~v_708 | v_136 | v_135 | ~v_707 | ~v_706 | v_162 | v_161 | ~v_2321 | ~v_2237 | ~v_2320 | ~v_2236 | ~v_2235 | ~v_2319 | ~v_2234 | ~v_2318 | ~v_2233 | ~v_2232 | ~v_233 | ~v_232 | ~v_1952 | ~v_1868 | ~v_1951 | ~v_1867 | ~v_1866 | ~v_1950 | ~v_1865 | ~v_1949 | ~v_1864 | ~v_1863 | ~v_4440 | ~v_4439 | ~v_4438 | ~v_4437 | v_4509;
assign x_128 = v_4508 | ~v_4505;
assign x_129 = v_4508 | ~v_4506;
assign x_130 = v_4508 | ~v_4507;
assign x_131 = v_101 | v_100 | v_94 | v_99 | v_93 | v_92 | v_102 | v_172 | v_171 | v_149 | v_148 | v_147 | ~v_2331 | ~v_2330 | ~v_2265 | ~v_2329 | ~v_2328 | ~v_2262 | ~v_483 | ~v_482 | ~v_2351 | ~v_2350 | ~v_2349 | ~v_2348 | ~v_593 | ~v_592 | ~v_545 | ~v_591 | ~v_590 | ~v_544 | ~v_1962 | ~v_1961 | ~v_1896 | ~v_1960 | ~v_1959 | ~v_1893 | ~v_2014 | ~v_2013 | ~v_2012 | ~v_2011 | ~v_4450 | ~v_4449 | ~v_4448 | ~v_4447 | v_4507;
assign x_132 = v_52 | v_50 | v_51 | v_60 | v_59 | v_58 | v_57 | v_144 | v_143 | v_142 | v_168 | v_167 | ~v_2326 | ~v_2325 | ~v_2250 | ~v_2324 | ~v_2323 | ~v_2247 | ~v_468 | ~v_467 | ~v_2346 | ~v_2345 | ~v_2344 | ~v_2343 | ~v_588 | ~v_587 | ~v_530 | ~v_586 | ~v_585 | ~v_529 | ~v_1957 | ~v_1956 | ~v_1881 | ~v_1955 | ~v_1954 | ~v_1878 | ~v_2009 | ~v_2008 | ~v_2007 | ~v_2006 | ~v_4445 | ~v_4444 | ~v_4443 | ~v_4442 | v_4506;
assign x_133 = v_9 | v_7 | v_17 | v_16 | v_8 | v_15 | v_14 | ~v_453 | ~v_452 | v_136 | v_135 | v_134 | v_164 | v_163 | ~v_2321 | ~v_2320 | ~v_2235 | ~v_2319 | ~v_2318 | ~v_2232 | ~v_2341 | ~v_2340 | ~v_2339 | ~v_2338 | ~v_583 | ~v_582 | ~v_515 | ~v_581 | ~v_580 | ~v_514 | ~v_1952 | ~v_1951 | ~v_1866 | ~v_1950 | ~v_1949 | ~v_1863 | ~v_2004 | ~v_2003 | ~v_2002 | ~v_2001 | ~v_4440 | ~v_4439 | ~v_4438 | ~v_4437 | v_4505;
assign x_134 = v_4504 | ~v_4501;
assign x_135 = v_4504 | ~v_4502;
assign x_136 = v_4504 | ~v_4503;
assign x_137 = v_103 | v_101 | v_97 | v_96 | v_100 | v_95 | v_94 | v_93 | v_92 | v_102 | v_171 | v_150 | ~v_2265 | ~v_2262 | ~v_2351 | ~v_2350 | ~v_2349 | ~v_2348 | ~v_545 | ~v_544 | ~v_2299 | ~v_2298 | ~v_2297 | ~v_2296 | ~v_561 | ~v_560 | ~v_559 | ~v_558 | ~v_387 | ~v_386 | ~v_1896 | ~v_1893 | ~v_2014 | ~v_2013 | ~v_2012 | ~v_2011 | ~v_1946 | ~v_1945 | ~v_1944 | ~v_1943 | ~v_4450 | ~v_4449 | ~v_4448 | ~v_4447 | v_4503;
assign x_138 = v_54 | v_53 | v_55 | v_61 | v_52 | v_50 | v_51 | v_60 | v_59 | v_58 | v_145 | v_167 | ~v_2250 | ~v_2247 | ~v_2346 | ~v_2345 | ~v_2344 | ~v_2343 | ~v_530 | ~v_529 | ~v_2294 | ~v_2293 | ~v_2292 | ~v_2291 | ~v_556 | ~v_555 | ~v_554 | ~v_553 | ~v_372 | ~v_371 | ~v_1881 | ~v_1878 | ~v_2009 | ~v_2008 | ~v_2007 | ~v_2006 | ~v_1941 | ~v_1940 | ~v_1939 | ~v_1938 | ~v_4445 | ~v_4444 | ~v_4443 | ~v_4442 | v_4502;
assign x_139 = v_9 | v_7 | v_18 | v_17 | v_16 | v_8 | v_15 | v_12 | v_11 | v_10 | v_137 | v_163 | ~v_2235 | ~v_2232 | ~v_2341 | ~v_2340 | ~v_2339 | ~v_2338 | ~v_515 | ~v_514 | ~v_2289 | ~v_2288 | ~v_2287 | ~v_2286 | ~v_551 | ~v_550 | ~v_549 | ~v_548 | ~v_357 | ~v_356 | ~v_1866 | ~v_1863 | ~v_2004 | ~v_2003 | ~v_2002 | ~v_2001 | ~v_1936 | ~v_1935 | ~v_1934 | ~v_1933 | ~v_4440 | ~v_4439 | ~v_4438 | ~v_4437 | v_4501;
assign x_140 = v_4500 | ~v_4497;
assign x_141 = v_4500 | ~v_4498;
assign x_142 = v_4500 | ~v_4499;
assign x_143 = v_103 | v_101 | v_100 | v_94 | v_93 | v_92 | v_151 | v_171 | v_150 | v_149 | v_148 | v_147 | ~v_577 | ~v_576 | ~v_2265 | ~v_2262 | ~v_2351 | ~v_2350 | ~v_2349 | ~v_2348 | ~v_545 | ~v_544 | ~v_2261 | ~v_2260 | ~v_2259 | ~v_2258 | ~v_575 | ~v_574 | ~v_435 | ~v_434 | ~v_1896 | ~v_1893 | ~v_2014 | ~v_2013 | ~v_2012 | ~v_2011 | ~v_1930 | ~v_1929 | ~v_1928 | ~v_1927 | ~v_4450 | ~v_4449 | ~v_4448 | ~v_4447 | v_4499;
assign x_144 = v_61 | v_52 | v_50 | v_51 | v_59 | v_58 | v_144 | v_145 | v_143 | v_142 | v_167 | v_146 | ~v_572 | ~v_571 | ~v_2250 | ~v_2247 | ~v_2346 | ~v_2345 | ~v_2344 | ~v_2343 | ~v_530 | ~v_529 | ~v_2246 | ~v_2245 | ~v_2244 | ~v_2243 | ~v_570 | ~v_569 | ~v_420 | ~v_419 | ~v_1881 | ~v_1878 | ~v_2009 | ~v_2008 | ~v_2007 | ~v_2006 | ~v_1925 | ~v_1924 | ~v_1923 | ~v_1922 | ~v_4445 | ~v_4444 | ~v_4443 | ~v_4442 | v_4498;
assign x_145 = v_9 | v_7 | v_18 | v_16 | v_8 | v_15 | v_136 | v_135 | v_134 | v_137 | v_138 | v_163 | ~v_567 | ~v_566 | ~v_2235 | ~v_2232 | ~v_2341 | ~v_2340 | ~v_2339 | ~v_2338 | ~v_515 | ~v_514 | ~v_2231 | ~v_2230 | ~v_2229 | ~v_2228 | ~v_565 | ~v_564 | ~v_405 | ~v_404 | ~v_1866 | ~v_1863 | ~v_2004 | ~v_2003 | ~v_2002 | ~v_2001 | ~v_1920 | ~v_1919 | ~v_1918 | ~v_1917 | ~v_4440 | ~v_4439 | ~v_4438 | ~v_4437 | v_4497;
assign x_146 = v_4496 | ~v_4493;
assign x_147 = v_4496 | ~v_4494;
assign x_148 = v_4496 | ~v_4495;
assign x_149 = v_103 | v_100 | v_94 | v_93 | v_92 | v_102 | v_171 | v_160 | v_150 | v_149 | v_148 | v_147 | ~v_2265 | ~v_2262 | ~v_2351 | ~v_2350 | ~v_2349 | ~v_2348 | ~v_545 | ~v_544 | ~v_2315 | ~v_2314 | ~v_2313 | ~v_2312 | ~v_543 | ~v_542 | ~v_541 | ~v_540 | ~v_297 | ~v_296 | ~v_1896 | ~v_1893 | ~v_2014 | ~v_2013 | ~v_2012 | ~v_2011 | ~v_1892 | ~v_1891 | ~v_1890 | ~v_1889 | ~v_4450 | ~v_4449 | ~v_4448 | ~v_4447 | v_4495;
assign x_150 = v_61 | v_52 | v_50 | v_51 | v_60 | v_58 | v_144 | v_159 | v_145 | v_143 | v_142 | v_167 | ~v_2250 | ~v_2247 | ~v_2346 | ~v_2345 | ~v_2344 | ~v_2343 | ~v_530 | ~v_529 | ~v_2310 | ~v_2309 | ~v_2308 | ~v_2307 | ~v_528 | ~v_527 | ~v_526 | ~v_525 | ~v_264 | ~v_263 | ~v_1881 | ~v_1878 | ~v_2009 | ~v_2008 | ~v_2007 | ~v_2006 | ~v_1877 | ~v_1876 | ~v_1875 | ~v_1874 | ~v_4445 | ~v_4444 | ~v_4443 | ~v_4442 | v_4494;
assign x_151 = v_9 | v_7 | v_18 | v_17 | v_8 | v_15 | v_136 | v_135 | v_134 | v_137 | v_163 | v_155 | ~v_2235 | ~v_2232 | ~v_2341 | ~v_2340 | ~v_2339 | ~v_2338 | ~v_515 | ~v_514 | ~v_2305 | ~v_2304 | ~v_2303 | ~v_2302 | ~v_513 | ~v_512 | ~v_511 | ~v_510 | ~v_231 | ~v_230 | ~v_1866 | ~v_1863 | ~v_2004 | ~v_2003 | ~v_2002 | ~v_2001 | ~v_1862 | ~v_1861 | ~v_1860 | ~v_1859 | ~v_4440 | ~v_4439 | ~v_4438 | ~v_4437 | v_4493;
assign x_152 = v_4492 | ~v_4489;
assign x_153 = v_4492 | ~v_4490;
assign x_154 = v_4492 | ~v_4491;
assign x_155 = v_98 | v_103 | v_101 | v_97 | v_96 | v_100 | v_92 | v_151 | v_170 | v_169 | v_150 | v_147 | ~v_2267 | ~v_2266 | ~v_2265 | ~v_2264 | ~v_2263 | ~v_2262 | ~v_299 | ~v_298 | ~v_2299 | ~v_2298 | ~v_2297 | ~v_2296 | ~v_387 | ~v_386 | ~v_499 | ~v_498 | ~v_497 | ~v_496 | ~v_1898 | ~v_1897 | ~v_1896 | ~v_1895 | ~v_1894 | ~v_1893 | ~v_1946 | ~v_1945 | ~v_1944 | ~v_1943 | ~v_4450 | ~v_4449 | ~v_4448 | ~v_4447 | v_4491;
assign x_156 = v_54 | v_56 | v_55 | v_61 | v_50 | v_59 | v_58 | v_145 | v_142 | v_166 | v_165 | v_146 | ~v_266 | ~v_2252 | ~v_2251 | ~v_2250 | ~v_2249 | ~v_2248 | ~v_2247 | ~v_265 | ~v_2294 | ~v_2293 | ~v_2292 | ~v_2291 | ~v_372 | ~v_371 | ~v_494 | ~v_493 | ~v_492 | ~v_491 | ~v_1883 | ~v_1882 | ~v_1881 | ~v_1880 | ~v_1879 | ~v_1878 | ~v_1941 | ~v_1940 | ~v_1939 | ~v_1938 | ~v_4445 | ~v_4444 | ~v_4443 | ~v_4442 | v_4490;
assign x_157 = v_13 | v_7 | v_18 | v_16 | v_15 | v_12 | v_11 | v_134 | v_137 | v_138 | v_162 | v_161 | ~v_2237 | ~v_2236 | ~v_2235 | ~v_2234 | ~v_2233 | ~v_2232 | ~v_233 | ~v_232 | ~v_2289 | ~v_2288 | ~v_2287 | ~v_2286 | ~v_357 | ~v_356 | ~v_489 | ~v_488 | ~v_487 | ~v_486 | ~v_1868 | ~v_1867 | ~v_1866 | ~v_1865 | ~v_1864 | ~v_1863 | ~v_1936 | ~v_1935 | ~v_1934 | ~v_1933 | ~v_4440 | ~v_4439 | ~v_4438 | ~v_4437 | v_4489;
assign x_158 = v_4488 | ~v_4485;
assign x_159 = v_4488 | ~v_4486;
assign x_160 = v_4488 | ~v_4487;
assign x_161 = v_103 | v_101 | v_100 | v_99 | v_92 | v_102 | v_171 | v_170 | v_169 | v_149 | v_148 | v_147 | ~v_703 | ~v_702 | ~v_2331 | ~v_2330 | ~v_2265 | ~v_2329 | ~v_2328 | ~v_2262 | ~v_483 | ~v_482 | ~v_2283 | ~v_2282 | ~v_2281 | ~v_2280 | ~v_701 | ~v_653 | ~v_700 | ~v_652 | ~v_1962 | ~v_1961 | ~v_1896 | ~v_1960 | ~v_1959 | ~v_1893 | ~v_1982 | ~v_1981 | ~v_1980 | ~v_1979 | ~v_4450 | ~v_4449 | ~v_4448 | ~v_4447 | v_4487;
assign x_162 = v_61 | v_50 | v_60 | v_59 | v_58 | v_57 | v_144 | v_143 | v_142 | v_167 | v_166 | v_165 | ~v_698 | ~v_697 | ~v_2326 | ~v_2325 | ~v_2250 | ~v_2324 | ~v_2323 | ~v_2247 | ~v_468 | ~v_467 | ~v_2278 | ~v_2277 | ~v_2276 | ~v_2275 | ~v_696 | ~v_638 | ~v_695 | ~v_637 | ~v_1957 | ~v_1956 | ~v_1881 | ~v_1955 | ~v_1954 | ~v_1878 | ~v_1977 | ~v_1976 | ~v_1975 | ~v_1974 | ~v_4445 | ~v_4444 | ~v_4443 | ~v_4442 | v_4486;
assign x_163 = v_7 | v_18 | v_17 | v_16 | v_15 | v_14 | ~v_453 | ~v_452 | v_136 | v_135 | v_134 | v_163 | v_162 | v_161 | ~v_693 | ~v_692 | ~v_2321 | ~v_2320 | ~v_2235 | ~v_2319 | ~v_2318 | ~v_2232 | ~v_2273 | ~v_2272 | ~v_2271 | ~v_2270 | ~v_691 | ~v_623 | ~v_690 | ~v_622 | ~v_1952 | ~v_1951 | ~v_1866 | ~v_1950 | ~v_1949 | ~v_1863 | ~v_1972 | ~v_1971 | ~v_1970 | ~v_1969 | ~v_4440 | ~v_4439 | ~v_4438 | ~v_4437 | v_4485;
assign x_164 = v_4484 | ~v_4481;
assign x_165 = v_4484 | ~v_4482;
assign x_166 = v_4484 | ~v_4483;
assign x_167 = v_101 | v_97 | v_96 | v_100 | v_92 | v_102 | v_172 | v_171 | v_170 | v_169 | v_150 | v_147 | ~v_671 | ~v_670 | ~v_2265 | ~v_2262 | ~v_2299 | ~v_2298 | ~v_2297 | ~v_2296 | ~v_387 | ~v_386 | ~v_2283 | ~v_2282 | ~v_2281 | ~v_2280 | ~v_653 | ~v_652 | ~v_669 | ~v_668 | ~v_1896 | ~v_1893 | ~v_1946 | ~v_1945 | ~v_1944 | ~v_1943 | ~v_1982 | ~v_1981 | ~v_1980 | ~v_1979 | ~v_4450 | ~v_4449 | ~v_4448 | ~v_4447 | v_4483;
assign x_168 = v_54 | v_55 | v_50 | v_60 | v_59 | v_58 | v_145 | v_142 | v_168 | v_167 | v_166 | v_165 | ~v_666 | ~v_665 | ~v_2250 | ~v_2247 | ~v_2294 | ~v_2293 | ~v_2292 | ~v_2291 | ~v_372 | ~v_371 | ~v_2278 | ~v_2277 | ~v_2276 | ~v_2275 | ~v_638 | ~v_637 | ~v_664 | ~v_663 | ~v_1881 | ~v_1878 | ~v_1941 | ~v_1940 | ~v_1939 | ~v_1938 | ~v_1977 | ~v_1976 | ~v_1975 | ~v_1974 | ~v_4445 | ~v_4444 | ~v_4443 | ~v_4442 | v_4482;
assign x_169 = v_7 | v_17 | v_16 | v_15 | v_12 | v_11 | v_134 | v_137 | v_164 | v_163 | v_162 | v_161 | ~v_661 | ~v_660 | ~v_2235 | ~v_2232 | ~v_2289 | ~v_2288 | ~v_2287 | ~v_2286 | ~v_357 | ~v_356 | ~v_2273 | ~v_2272 | ~v_2271 | ~v_2270 | ~v_623 | ~v_622 | ~v_659 | ~v_658 | ~v_1866 | ~v_1863 | ~v_1936 | ~v_1935 | ~v_1934 | ~v_1933 | ~v_1972 | ~v_1971 | ~v_1970 | ~v_1969 | ~v_4440 | ~v_4439 | ~v_4438 | ~v_4437 | v_4481;
assign x_170 = v_4480 | ~v_4477;
assign x_171 = v_4480 | ~v_4478;
assign x_172 = v_4480 | ~v_4479;
assign x_173 = v_103 | v_101 | v_100 | v_95 | v_92 | v_102 | v_171 | v_170 | v_169 | v_150 | v_149 | v_148 | ~v_2265 | ~v_2262 | ~v_2261 | ~v_2260 | ~v_2259 | ~v_2258 | ~v_435 | ~v_434 | ~v_2283 | ~v_2282 | ~v_2281 | ~v_2280 | ~v_653 | ~v_652 | ~v_687 | ~v_686 | ~v_685 | ~v_684 | ~v_1896 | ~v_1893 | ~v_1930 | ~v_1929 | ~v_1928 | ~v_1927 | ~v_1982 | ~v_1981 | ~v_1980 | ~v_1979 | ~v_4450 | ~v_4449 | ~v_4448 | ~v_4447 | v_4479;
assign x_174 = v_53 | v_61 | v_50 | v_60 | v_59 | v_58 | v_144 | v_145 | v_143 | v_167 | v_166 | v_165 | ~v_2250 | ~v_2247 | ~v_2246 | ~v_2245 | ~v_2244 | ~v_2243 | ~v_420 | ~v_419 | ~v_2278 | ~v_2277 | ~v_2276 | ~v_2275 | ~v_638 | ~v_637 | ~v_682 | ~v_681 | ~v_680 | ~v_679 | ~v_1881 | ~v_1878 | ~v_1925 | ~v_1924 | ~v_1923 | ~v_1922 | ~v_1977 | ~v_1976 | ~v_1975 | ~v_1974 | ~v_4445 | ~v_4444 | ~v_4443 | ~v_4442 | v_4478;
assign x_175 = v_7 | v_18 | v_17 | v_16 | v_15 | v_10 | v_136 | v_135 | v_137 | v_163 | v_162 | v_161 | ~v_2235 | ~v_2232 | ~v_2231 | ~v_2230 | ~v_2229 | ~v_2228 | ~v_405 | ~v_404 | ~v_2273 | ~v_2272 | ~v_2271 | ~v_2270 | ~v_623 | ~v_622 | ~v_677 | ~v_676 | ~v_675 | ~v_674 | ~v_1866 | ~v_1863 | ~v_1920 | ~v_1919 | ~v_1918 | ~v_1917 | ~v_1972 | ~v_1971 | ~v_1970 | ~v_1969 | ~v_4440 | ~v_4439 | ~v_4438 | ~v_4437 | v_4477;
assign x_176 = v_4476 | ~v_4473;
assign x_177 = v_4476 | ~v_4474;
assign x_178 = v_4476 | ~v_4475;
assign x_179 = v_103 | v_100 | v_92 | v_151 | v_171 | v_170 | v_169 | v_160 | v_150 | v_149 | v_148 | v_147 | ~v_655 | ~v_654 | ~v_2265 | ~v_2262 | ~v_2315 | ~v_2314 | ~v_2313 | ~v_2312 | ~v_297 | ~v_296 | ~v_2283 | ~v_2282 | ~v_2281 | ~v_2280 | ~v_653 | ~v_652 | ~v_651 | ~v_650 | ~v_1896 | ~v_1893 | ~v_1892 | ~v_1891 | ~v_1890 | ~v_1889 | ~v_1982 | ~v_1981 | ~v_1980 | ~v_1979 | ~v_4450 | ~v_4449 | ~v_4448 | ~v_4447 | v_4475;
assign x_180 = v_61 | v_50 | v_58 | v_144 | v_159 | v_145 | v_143 | v_142 | v_167 | v_166 | v_165 | v_146 | ~v_640 | ~v_639 | ~v_2250 | ~v_2247 | ~v_2310 | ~v_2309 | ~v_2308 | ~v_2307 | ~v_264 | ~v_263 | ~v_2278 | ~v_2277 | ~v_2276 | ~v_2275 | ~v_638 | ~v_637 | ~v_636 | ~v_635 | ~v_1881 | ~v_1878 | ~v_1877 | ~v_1876 | ~v_1875 | ~v_1874 | ~v_1977 | ~v_1976 | ~v_1975 | ~v_1974 | ~v_4445 | ~v_4444 | ~v_4443 | ~v_4442 | v_4474;
assign x_181 = v_7 | v_18 | v_15 | v_136 | v_135 | v_134 | v_137 | v_138 | v_163 | v_162 | v_161 | v_155 | ~v_625 | ~v_624 | ~v_2235 | ~v_2232 | ~v_2305 | ~v_2304 | ~v_2303 | ~v_2302 | ~v_231 | ~v_230 | ~v_2273 | ~v_2272 | ~v_2271 | ~v_2270 | ~v_623 | ~v_622 | ~v_621 | ~v_620 | ~v_1866 | ~v_1863 | ~v_1862 | ~v_1861 | ~v_1860 | ~v_1859 | ~v_1972 | ~v_1971 | ~v_1970 | ~v_1969 | ~v_4440 | ~v_4439 | ~v_4438 | ~v_4437 | v_4473;
assign x_182 = v_4472 | ~v_4469;
assign x_183 = v_4472 | ~v_4470;
assign x_184 = v_4472 | ~v_4471;
assign x_185 = v_98 | v_103 | v_101 | v_100 | v_92 | v_102 | v_170 | v_169 | v_150 | v_149 | v_148 | v_147 | ~v_609 | ~v_608 | ~v_2267 | ~v_2266 | ~v_2265 | ~v_2264 | ~v_2263 | ~v_2262 | ~v_299 | ~v_298 | ~v_2261 | ~v_2260 | ~v_2259 | ~v_2258 | ~v_435 | ~v_434 | ~v_607 | ~v_606 | ~v_1898 | ~v_1897 | ~v_1896 | ~v_1895 | ~v_1894 | ~v_1893 | ~v_1930 | ~v_1929 | ~v_1928 | ~v_1927 | ~v_4450 | ~v_4449 | ~v_4448 | ~v_4447 | v_4471;
assign x_186 = v_56 | v_61 | v_50 | v_60 | v_59 | v_58 | v_144 | v_145 | v_143 | v_142 | v_166 | v_165 | ~v_604 | ~v_603 | ~v_266 | ~v_2252 | ~v_2251 | ~v_2250 | ~v_2249 | ~v_2248 | ~v_2247 | ~v_265 | ~v_2246 | ~v_2245 | ~v_2244 | ~v_2243 | ~v_420 | ~v_419 | ~v_602 | ~v_601 | ~v_1883 | ~v_1882 | ~v_1881 | ~v_1880 | ~v_1879 | ~v_1878 | ~v_1925 | ~v_1924 | ~v_1923 | ~v_1922 | ~v_4445 | ~v_4444 | ~v_4443 | ~v_4442 | v_4470;
assign x_187 = v_13 | v_7 | v_18 | v_17 | v_16 | v_15 | v_136 | v_135 | v_134 | v_137 | v_162 | v_161 | ~v_599 | ~v_598 | ~v_2237 | ~v_2236 | ~v_2235 | ~v_2234 | ~v_2233 | ~v_2232 | ~v_233 | ~v_232 | ~v_2231 | ~v_2230 | ~v_2229 | ~v_2228 | ~v_405 | ~v_404 | ~v_597 | ~v_596 | ~v_1868 | ~v_1867 | ~v_1866 | ~v_1865 | ~v_1864 | ~v_1863 | ~v_1920 | ~v_1919 | ~v_1918 | ~v_1917 | ~v_4440 | ~v_4439 | ~v_4438 | ~v_4437 | v_4469;
assign x_188 = v_4468 | ~v_4465;
assign x_189 = v_4468 | ~v_4466;
assign x_190 = v_4468 | ~v_4467;
assign x_191 = v_103 | v_101 | v_99 | v_92 | v_102 | v_171 | v_170 | v_169 | v_149 | v_148 | v_147 | v_181 | ~v_2331 | ~v_2330 | ~v_2265 | ~v_2329 | ~v_2328 | ~v_2262 | ~v_483 | ~v_482 | ~v_2383 | ~v_2382 | ~v_2381 | ~v_2380 | ~v_481 | ~v_480 | ~v_345 | ~v_479 | ~v_478 | ~v_344 | ~v_1962 | ~v_1961 | ~v_1896 | ~v_1960 | ~v_1959 | ~v_1893 | ~v_1914 | ~v_1913 | ~v_1912 | ~v_1911 | ~v_4450 | ~v_4449 | ~v_4448 | ~v_4447 | v_4467;
assign x_192 = v_61 | v_50 | v_60 | v_59 | v_57 | v_144 | v_180 | v_143 | v_142 | v_167 | v_166 | v_165 | ~v_2326 | ~v_2325 | ~v_2250 | ~v_2324 | ~v_2323 | ~v_2247 | ~v_468 | ~v_467 | ~v_2378 | ~v_2377 | ~v_2376 | ~v_2375 | ~v_466 | ~v_465 | ~v_330 | ~v_464 | ~v_463 | ~v_329 | ~v_1957 | ~v_1956 | ~v_1881 | ~v_1955 | ~v_1954 | ~v_1878 | ~v_1909 | ~v_1908 | ~v_1907 | ~v_1906 | ~v_4445 | ~v_4444 | ~v_4443 | ~v_4442 | v_4466;
assign x_193 = v_7 | v_18 | v_17 | v_16 | v_14 | ~v_453 | ~v_452 | v_136 | v_135 | v_134 | v_179 | v_163 | v_162 | v_161 | ~v_2321 | ~v_2320 | ~v_2235 | ~v_2319 | ~v_2318 | ~v_2232 | ~v_2373 | ~v_2372 | ~v_2371 | ~v_2370 | ~v_451 | ~v_450 | ~v_315 | ~v_449 | ~v_448 | ~v_314 | ~v_1952 | ~v_1951 | ~v_1866 | ~v_1950 | ~v_1949 | ~v_1863 | ~v_1904 | ~v_1903 | ~v_1902 | ~v_1901 | ~v_4440 | ~v_4439 | ~v_4438 | ~v_4437 | v_4465;
assign x_194 = v_4464 | ~v_4461;
assign x_195 = v_4464 | ~v_4462;
assign x_196 = v_4464 | ~v_4463;
assign x_197 = v_103 | v_101 | v_97 | v_96 | v_92 | v_102 | v_171 | v_170 | v_169 | v_150 | v_147 | v_181 | ~v_391 | ~v_390 | ~v_2265 | ~v_2262 | ~v_2299 | ~v_2298 | ~v_2297 | ~v_2296 | ~v_387 | ~v_386 | ~v_2383 | ~v_2382 | ~v_2381 | ~v_2380 | ~v_345 | ~v_344 | ~v_385 | ~v_384 | ~v_1896 | ~v_1893 | ~v_1946 | ~v_1945 | ~v_1944 | ~v_1943 | ~v_1914 | ~v_1913 | ~v_1912 | ~v_1911 | ~v_4450 | ~v_4449 | ~v_4448 | ~v_4447 | v_4463;
assign x_198 = v_54 | v_55 | v_61 | v_50 | v_60 | v_59 | v_180 | v_145 | v_142 | v_167 | v_166 | v_165 | ~v_376 | ~v_375 | ~v_2250 | ~v_2247 | ~v_2294 | ~v_2293 | ~v_2292 | ~v_2291 | ~v_372 | ~v_371 | ~v_2378 | ~v_2377 | ~v_2376 | ~v_2375 | ~v_330 | ~v_329 | ~v_370 | ~v_369 | ~v_1881 | ~v_1878 | ~v_1941 | ~v_1940 | ~v_1939 | ~v_1938 | ~v_1909 | ~v_1908 | ~v_1907 | ~v_1906 | ~v_4445 | ~v_4444 | ~v_4443 | ~v_4442 | v_4462;
assign x_199 = v_7 | v_18 | v_17 | v_16 | v_12 | v_11 | v_134 | v_137 | v_179 | v_163 | v_162 | v_161 | ~v_361 | ~v_360 | ~v_2235 | ~v_2232 | ~v_2289 | ~v_2288 | ~v_2287 | ~v_2286 | ~v_357 | ~v_356 | ~v_2373 | ~v_2372 | ~v_2371 | ~v_2370 | ~v_315 | ~v_314 | ~v_355 | ~v_354 | ~v_1866 | ~v_1863 | ~v_1936 | ~v_1935 | ~v_1934 | ~v_1933 | ~v_1904 | ~v_1903 | ~v_1902 | ~v_1901 | ~v_4440 | ~v_4439 | ~v_4438 | ~v_4437 | v_4461;
assign x_200 = v_4460 | ~v_4457;
assign x_201 = v_4460 | ~v_4458;
assign x_202 = v_4460 | ~v_4459;
assign x_203 = v_101 | v_92 | v_102 | v_172 | v_171 | v_170 | v_169 | v_150 | v_149 | v_148 | v_147 | v_181 | ~v_437 | ~v_436 | ~v_2265 | ~v_2262 | ~v_2261 | ~v_2260 | ~v_2259 | ~v_2258 | ~v_435 | ~v_434 | ~v_2383 | ~v_2382 | ~v_2381 | ~v_2380 | ~v_345 | ~v_344 | ~v_433 | ~v_432 | ~v_1896 | ~v_1893 | ~v_1930 | ~v_1929 | ~v_1928 | ~v_1927 | ~v_1914 | ~v_1913 | ~v_1912 | ~v_1911 | ~v_4450 | ~v_4449 | ~v_4448 | ~v_4447 | v_4459;
assign x_204 = v_50 | v_60 | v_59 | v_144 | v_180 | v_145 | v_143 | v_142 | v_168 | v_167 | v_166 | v_165 | ~v_422 | ~v_421 | ~v_2250 | ~v_2247 | ~v_2246 | ~v_2245 | ~v_2244 | ~v_2243 | ~v_420 | ~v_419 | ~v_2378 | ~v_2377 | ~v_2376 | ~v_2375 | ~v_330 | ~v_329 | ~v_418 | ~v_417 | ~v_1881 | ~v_1878 | ~v_1925 | ~v_1924 | ~v_1923 | ~v_1922 | ~v_1909 | ~v_1908 | ~v_1907 | ~v_1906 | ~v_4445 | ~v_4444 | ~v_4443 | ~v_4442 | v_4458;
assign x_205 = v_7 | v_17 | v_16 | v_136 | v_135 | v_134 | v_137 | v_179 | v_164 | v_163 | v_162 | v_161 | ~v_407 | ~v_406 | ~v_2235 | ~v_2232 | ~v_2231 | ~v_2230 | ~v_2229 | ~v_2228 | ~v_405 | ~v_404 | ~v_2373 | ~v_2372 | ~v_2371 | ~v_2370 | ~v_315 | ~v_314 | ~v_403 | ~v_402 | ~v_1866 | ~v_1863 | ~v_1920 | ~v_1919 | ~v_1918 | ~v_1917 | ~v_1904 | ~v_1903 | ~v_1902 | ~v_1901 | ~v_4440 | ~v_4439 | ~v_4438 | ~v_4437 | v_4457;
assign x_206 = v_4456 | ~v_4453;
assign x_207 = v_4456 | ~v_4454;
assign x_208 = v_4456 | ~v_4455;
assign x_209 = v_103 | v_95 | v_92 | v_102 | v_171 | v_170 | v_169 | v_160 | v_150 | v_149 | v_148 | v_181 | ~v_2265 | ~v_2262 | ~v_2315 | ~v_2314 | ~v_2313 | ~v_2312 | ~v_297 | ~v_296 | ~v_2383 | ~v_2382 | ~v_2381 | ~v_2380 | ~v_345 | ~v_344 | ~v_343 | ~v_342 | ~v_341 | ~v_340 | ~v_1896 | ~v_1893 | ~v_1892 | ~v_1891 | ~v_1890 | ~v_1889 | ~v_1914 | ~v_1913 | ~v_1912 | ~v_1911 | ~v_4450 | ~v_4449 | ~v_4448 | ~v_4447 | v_4455;
assign x_210 = v_53 | v_61 | v_50 | v_60 | v_144 | v_180 | v_159 | v_145 | v_143 | v_167 | v_166 | v_165 | ~v_2250 | ~v_2247 | ~v_2310 | ~v_2309 | ~v_2308 | ~v_2307 | ~v_264 | ~v_263 | ~v_2378 | ~v_2377 | ~v_2376 | ~v_2375 | ~v_330 | ~v_329 | ~v_328 | ~v_327 | ~v_326 | ~v_325 | ~v_1881 | ~v_1878 | ~v_1877 | ~v_1876 | ~v_1875 | ~v_1874 | ~v_1909 | ~v_1908 | ~v_1907 | ~v_1906 | ~v_4445 | ~v_4444 | ~v_4443 | ~v_4442 | v_4454;
assign x_211 = v_7 | v_18 | v_17 | v_10 | v_136 | v_135 | v_137 | v_179 | v_163 | v_162 | v_161 | v_155 | ~v_2235 | ~v_2232 | ~v_2305 | ~v_2304 | ~v_2303 | ~v_2302 | ~v_231 | ~v_230 | ~v_2373 | ~v_2372 | ~v_2371 | ~v_2370 | ~v_315 | ~v_314 | ~v_313 | ~v_312 | ~v_311 | ~v_310 | ~v_1866 | ~v_1863 | ~v_1862 | ~v_1861 | ~v_1860 | ~v_1859 | ~v_1904 | ~v_1903 | ~v_1902 | ~v_1901 | ~v_4440 | ~v_4439 | ~v_4438 | ~v_4437 | v_4453;
assign x_212 = v_4452 | ~v_4441;
assign x_213 = v_4452 | ~v_4446;
assign x_214 = v_4452 | ~v_4451;
assign x_215 = v_98 | v_103 | v_100 | v_92 | v_102 | v_170 | v_169 | v_160 | v_150 | v_149 | v_148 | v_147 | ~v_2267 | ~v_2266 | ~v_2265 | ~v_2264 | ~v_2263 | ~v_2262 | ~v_299 | ~v_298 | ~v_2315 | ~v_2314 | ~v_2313 | ~v_2312 | ~v_297 | ~v_296 | ~v_295 | ~v_294 | ~v_293 | ~v_292 | ~v_1898 | ~v_1897 | ~v_1896 | ~v_1895 | ~v_1894 | ~v_1893 | ~v_1892 | ~v_1891 | ~v_1890 | ~v_1889 | ~v_4450 | ~v_4449 | ~v_4448 | ~v_4447 | v_4451;
assign x_216 = v_4450 | v_141;
assign x_217 = v_4450 | v_123;
assign x_218 = v_4449 | v_141;
assign x_219 = v_4449 | v_120;
assign x_220 = v_4448 | ~v_141;
assign x_221 = v_4448 | v_108;
assign x_222 = v_4447 | ~v_141;
assign x_223 = v_4447 | v_105;
assign x_224 = v_56 | v_61 | v_50 | v_60 | v_58 | v_144 | v_159 | v_145 | v_143 | v_142 | v_166 | v_165 | ~v_266 | ~v_2252 | ~v_2251 | ~v_2250 | ~v_2249 | ~v_2248 | ~v_2247 | ~v_265 | ~v_2310 | ~v_2309 | ~v_2308 | ~v_2307 | ~v_264 | ~v_263 | ~v_262 | ~v_261 | ~v_260 | ~v_259 | ~v_1883 | ~v_1882 | ~v_1881 | ~v_1880 | ~v_1879 | ~v_1878 | ~v_1877 | ~v_1876 | ~v_1875 | ~v_1874 | ~v_4445 | ~v_4444 | ~v_4443 | ~v_4442 | v_4446;
assign x_225 = v_4445 | v_141;
assign x_226 = v_4445 | v_81;
assign x_227 = v_4444 | v_141;
assign x_228 = v_4444 | v_78;
assign x_229 = v_4443 | ~v_141;
assign x_230 = v_4443 | v_66;
assign x_231 = v_4442 | ~v_141;
assign x_232 = v_4442 | v_63;
assign x_233 = v_13 | v_7 | v_18 | v_17 | v_15 | v_136 | v_135 | v_134 | v_137 | v_162 | v_161 | v_155 | ~v_2237 | ~v_2236 | ~v_2235 | ~v_2234 | ~v_2233 | ~v_2232 | ~v_233 | ~v_232 | ~v_2305 | ~v_2304 | ~v_2303 | ~v_2302 | ~v_231 | ~v_230 | ~v_229 | ~v_228 | ~v_227 | ~v_226 | ~v_1868 | ~v_1867 | ~v_1866 | ~v_1865 | ~v_1864 | ~v_1863 | ~v_1862 | ~v_1861 | ~v_1860 | ~v_1859 | ~v_4440 | ~v_4439 | ~v_4438 | ~v_4437 | v_4441;
assign x_234 = v_4440 | v_141;
assign x_235 = v_4440 | v_39;
assign x_236 = v_4439 | v_141;
assign x_237 = v_4439 | v_36;
assign x_238 = v_4438 | ~v_141;
assign x_239 = v_4438 | v_24;
assign x_240 = v_4437 | ~v_141;
assign x_241 = v_4437 | v_21;
assign x_242 = v_4436 | ~v_4433;
assign x_243 = v_4436 | ~v_4434;
assign x_244 = v_4436 | ~v_4435;
assign x_245 = v_98 | v_103 | v_101 | v_100 | v_95 | v_99 | v_92 | v_102 | ~v_719 | ~v_718 | v_170 | v_169 | v_149 | v_148 | ~v_483 | ~v_717 | ~v_299 | ~v_482 | ~v_716 | ~v_298 | ~v_1464 | ~v_1352 | ~v_1463 | ~v_1351 | ~v_1350 | ~v_1462 | ~v_1349 | ~v_1461 | ~v_1348 | ~v_1347 | ~v_477 | ~v_291 | ~v_476 | ~v_290 | ~v_289 | ~v_475 | ~v_288 | ~v_474 | ~v_287 | ~v_286 | ~v_4374 | ~v_4373 | ~v_4372 | ~v_4371 | v_4435;
assign x_246 = v_53 | v_56 | v_61 | v_50 | v_60 | v_59 | v_58 | v_57 | ~v_714 | ~v_713 | v_144 | v_143 | v_166 | v_165 | ~v_266 | ~v_468 | ~v_712 | ~v_467 | ~v_711 | ~v_265 | ~v_1455 | ~v_1327 | ~v_1454 | ~v_1326 | ~v_1325 | ~v_1453 | ~v_1324 | ~v_1452 | ~v_1323 | ~v_1322 | ~v_462 | ~v_258 | ~v_461 | ~v_257 | ~v_256 | ~v_460 | ~v_255 | ~v_459 | ~v_254 | ~v_253 | ~v_4369 | ~v_4368 | ~v_4367 | ~v_4366 | v_4434;
assign x_247 = v_13 | v_7 | v_18 | v_17 | v_16 | v_15 | v_14 | v_10 | ~v_453 | ~v_709 | ~v_452 | ~v_708 | v_136 | v_135 | ~v_707 | ~v_706 | v_162 | v_161 | ~v_233 | ~v_232 | ~v_1446 | ~v_1302 | ~v_1445 | ~v_1301 | ~v_1300 | ~v_1444 | ~v_1299 | ~v_1443 | ~v_1298 | ~v_1297 | ~v_447 | ~v_225 | ~v_446 | ~v_224 | ~v_223 | ~v_445 | ~v_222 | ~v_444 | ~v_221 | ~v_220 | ~v_4364 | ~v_4363 | ~v_4362 | ~v_4361 | v_4433;
assign x_248 = v_4432 | ~v_4429;
assign x_249 = v_4432 | ~v_4430;
assign x_250 = v_4432 | ~v_4431;
assign x_251 = v_103 | v_101 | v_100 | v_94 | v_99 | v_93 | v_92 | v_102 | v_171 | v_149 | v_148 | v_147 | ~v_703 | ~v_702 | ~v_483 | ~v_482 | ~v_701 | ~v_653 | ~v_700 | ~v_652 | ~v_1464 | ~v_1463 | ~v_1350 | ~v_1462 | ~v_1461 | ~v_1347 | ~v_1380 | ~v_1379 | ~v_1378 | ~v_1377 | ~v_477 | ~v_476 | ~v_289 | ~v_475 | ~v_474 | ~v_286 | ~v_649 | ~v_648 | ~v_647 | ~v_646 | ~v_4374 | ~v_4373 | ~v_4372 | ~v_4371 | v_4431;
assign x_252 = v_61 | v_52 | v_50 | v_51 | v_60 | v_59 | v_58 | v_57 | v_144 | v_143 | v_142 | v_167 | ~v_698 | ~v_697 | ~v_468 | ~v_467 | ~v_696 | ~v_638 | ~v_695 | ~v_637 | ~v_1455 | ~v_1454 | ~v_1325 | ~v_1453 | ~v_1452 | ~v_1322 | ~v_1371 | ~v_1370 | ~v_1369 | ~v_1368 | ~v_462 | ~v_461 | ~v_256 | ~v_460 | ~v_459 | ~v_253 | ~v_634 | ~v_633 | ~v_632 | ~v_631 | ~v_4369 | ~v_4368 | ~v_4367 | ~v_4366 | v_4430;
assign x_253 = v_9 | v_7 | v_18 | v_17 | v_16 | v_8 | v_15 | v_14 | ~v_453 | ~v_452 | v_136 | v_135 | v_134 | v_163 | ~v_693 | ~v_692 | ~v_691 | ~v_623 | ~v_690 | ~v_622 | ~v_1446 | ~v_1445 | ~v_1300 | ~v_1444 | ~v_1443 | ~v_1297 | ~v_1362 | ~v_1361 | ~v_1360 | ~v_1359 | ~v_447 | ~v_446 | ~v_223 | ~v_445 | ~v_444 | ~v_220 | ~v_619 | ~v_618 | ~v_617 | ~v_616 | ~v_4364 | ~v_4363 | ~v_4362 | ~v_4361 | v_4429;
assign x_254 = v_4428 | ~v_4425;
assign x_255 = v_4428 | ~v_4426;
assign x_256 = v_4428 | ~v_4427;
assign x_257 = v_103 | v_101 | v_97 | v_96 | v_100 | v_95 | v_94 | v_93 | v_92 | v_102 | v_171 | v_150 | ~v_435 | ~v_434 | ~v_653 | ~v_652 | ~v_687 | ~v_686 | ~v_685 | ~v_684 | ~v_1350 | ~v_1347 | ~v_1380 | ~v_1379 | ~v_1378 | ~v_1377 | ~v_1346 | ~v_1345 | ~v_1344 | ~v_1343 | ~v_289 | ~v_286 | ~v_649 | ~v_648 | ~v_647 | ~v_646 | ~v_431 | ~v_430 | ~v_429 | ~v_428 | ~v_4374 | ~v_4373 | ~v_4372 | ~v_4371 | v_4427;
assign x_258 = v_54 | v_53 | v_55 | v_61 | v_52 | v_50 | v_51 | v_60 | v_59 | v_58 | v_145 | v_167 | ~v_420 | ~v_419 | ~v_638 | ~v_637 | ~v_682 | ~v_681 | ~v_680 | ~v_679 | ~v_1325 | ~v_1322 | ~v_1371 | ~v_1370 | ~v_1369 | ~v_1368 | ~v_1321 | ~v_1320 | ~v_1319 | ~v_1318 | ~v_256 | ~v_253 | ~v_634 | ~v_633 | ~v_632 | ~v_631 | ~v_416 | ~v_415 | ~v_414 | ~v_413 | ~v_4369 | ~v_4368 | ~v_4367 | ~v_4366 | v_4426;
assign x_259 = v_9 | v_7 | v_18 | v_17 | v_16 | v_8 | v_15 | v_12 | v_11 | v_10 | v_137 | v_163 | ~v_405 | ~v_404 | ~v_623 | ~v_622 | ~v_677 | ~v_676 | ~v_675 | ~v_674 | ~v_1300 | ~v_1297 | ~v_1362 | ~v_1361 | ~v_1360 | ~v_1359 | ~v_1296 | ~v_1295 | ~v_1294 | ~v_1293 | ~v_223 | ~v_220 | ~v_619 | ~v_618 | ~v_617 | ~v_616 | ~v_401 | ~v_400 | ~v_399 | ~v_398 | ~v_4364 | ~v_4363 | ~v_4362 | ~v_4361 | v_4425;
assign x_260 = v_4424 | ~v_4421;
assign x_261 = v_4424 | ~v_4422;
assign x_262 = v_4424 | ~v_4423;
assign x_263 = v_101 | v_100 | v_94 | v_93 | v_92 | v_102 | v_172 | v_171 | v_150 | v_149 | v_148 | v_147 | ~v_671 | ~v_670 | ~v_387 | ~v_386 | ~v_653 | ~v_652 | ~v_669 | ~v_668 | ~v_1350 | ~v_1347 | ~v_1380 | ~v_1379 | ~v_1378 | ~v_1377 | ~v_1408 | ~v_1407 | ~v_1406 | ~v_1405 | ~v_289 | ~v_286 | ~v_649 | ~v_648 | ~v_647 | ~v_646 | ~v_383 | ~v_382 | ~v_381 | ~v_380 | ~v_4374 | ~v_4373 | ~v_4372 | ~v_4371 | v_4423;
assign x_264 = v_52 | v_50 | v_51 | v_60 | v_59 | v_58 | v_144 | v_145 | v_143 | v_142 | v_168 | v_167 | ~v_666 | ~v_665 | ~v_372 | ~v_371 | ~v_638 | ~v_637 | ~v_664 | ~v_663 | ~v_1325 | ~v_1322 | ~v_1371 | ~v_1370 | ~v_1369 | ~v_1368 | ~v_1399 | ~v_1398 | ~v_1397 | ~v_1396 | ~v_256 | ~v_253 | ~v_634 | ~v_633 | ~v_632 | ~v_631 | ~v_368 | ~v_367 | ~v_366 | ~v_365 | ~v_4369 | ~v_4368 | ~v_4367 | ~v_4366 | v_4422;
assign x_265 = v_9 | v_7 | v_17 | v_16 | v_8 | v_15 | v_136 | v_135 | v_134 | v_137 | v_164 | v_163 | ~v_661 | ~v_660 | ~v_357 | ~v_356 | ~v_623 | ~v_622 | ~v_659 | ~v_658 | ~v_1300 | ~v_1297 | ~v_1362 | ~v_1361 | ~v_1360 | ~v_1359 | ~v_1390 | ~v_1389 | ~v_1388 | ~v_1387 | ~v_223 | ~v_220 | ~v_619 | ~v_618 | ~v_617 | ~v_616 | ~v_353 | ~v_352 | ~v_351 | ~v_350 | ~v_4364 | ~v_4363 | ~v_4362 | ~v_4361 | v_4421;
assign x_266 = v_4420 | ~v_4417;
assign x_267 = v_4420 | ~v_4418;
assign x_268 = v_4420 | ~v_4419;
assign x_269 = v_103 | v_100 | v_94 | v_93 | v_92 | v_151 | v_171 | v_160 | v_150 | v_149 | v_148 | v_147 | ~v_655 | ~v_654 | ~v_297 | ~v_296 | ~v_653 | ~v_652 | ~v_651 | ~v_650 | ~v_1350 | ~v_1347 | ~v_1380 | ~v_1379 | ~v_1378 | ~v_1377 | ~v_1436 | ~v_1435 | ~v_1434 | ~v_1433 | ~v_289 | ~v_286 | ~v_649 | ~v_648 | ~v_647 | ~v_646 | ~v_285 | ~v_284 | ~v_283 | ~v_282 | ~v_4374 | ~v_4373 | ~v_4372 | ~v_4371 | v_4419;
assign x_270 = v_61 | v_52 | v_50 | v_51 | v_58 | v_144 | v_159 | v_145 | v_143 | v_142 | v_167 | v_146 | ~v_640 | ~v_639 | ~v_264 | ~v_263 | ~v_638 | ~v_637 | ~v_636 | ~v_635 | ~v_1325 | ~v_1322 | ~v_1371 | ~v_1370 | ~v_1369 | ~v_1368 | ~v_1427 | ~v_1426 | ~v_1425 | ~v_1424 | ~v_256 | ~v_253 | ~v_634 | ~v_633 | ~v_632 | ~v_631 | ~v_252 | ~v_251 | ~v_250 | ~v_249 | ~v_4369 | ~v_4368 | ~v_4367 | ~v_4366 | v_4418;
assign x_271 = v_9 | v_7 | v_18 | v_8 | v_15 | v_136 | v_135 | v_134 | v_137 | v_138 | v_163 | v_155 | ~v_625 | ~v_624 | ~v_231 | ~v_230 | ~v_623 | ~v_622 | ~v_621 | ~v_620 | ~v_1300 | ~v_1297 | ~v_1362 | ~v_1361 | ~v_1360 | ~v_1359 | ~v_1418 | ~v_1417 | ~v_1416 | ~v_1415 | ~v_223 | ~v_220 | ~v_619 | ~v_618 | ~v_617 | ~v_616 | ~v_219 | ~v_218 | ~v_217 | ~v_216 | ~v_4364 | ~v_4363 | ~v_4362 | ~v_4361 | v_4417;
assign x_272 = v_4416 | ~v_4413;
assign x_273 = v_4416 | ~v_4414;
assign x_274 = v_4416 | ~v_4415;
assign x_275 = v_98 | v_103 | v_101 | v_97 | v_96 | v_100 | v_92 | v_102 | v_170 | v_169 | v_150 | v_147 | ~v_609 | ~v_608 | ~v_299 | ~v_298 | ~v_435 | ~v_434 | ~v_607 | ~v_606 | ~v_1352 | ~v_1351 | ~v_1350 | ~v_1349 | ~v_1348 | ~v_1347 | ~v_1346 | ~v_1345 | ~v_1344 | ~v_1343 | ~v_291 | ~v_290 | ~v_289 | ~v_288 | ~v_287 | ~v_286 | ~v_431 | ~v_430 | ~v_429 | ~v_428 | ~v_4374 | ~v_4373 | ~v_4372 | ~v_4371 | v_4415;
assign x_276 = v_54 | v_56 | v_55 | v_61 | v_50 | v_60 | v_59 | v_58 | v_145 | v_142 | v_166 | v_165 | ~v_604 | ~v_603 | ~v_266 | ~v_265 | ~v_420 | ~v_419 | ~v_602 | ~v_601 | ~v_1327 | ~v_1326 | ~v_1325 | ~v_1324 | ~v_1323 | ~v_1322 | ~v_1321 | ~v_1320 | ~v_1319 | ~v_1318 | ~v_258 | ~v_257 | ~v_256 | ~v_255 | ~v_254 | ~v_253 | ~v_416 | ~v_415 | ~v_414 | ~v_413 | ~v_4369 | ~v_4368 | ~v_4367 | ~v_4366 | v_4414;
assign x_277 = v_13 | v_7 | v_18 | v_17 | v_16 | v_15 | v_12 | v_11 | v_134 | v_137 | v_162 | v_161 | ~v_599 | ~v_598 | ~v_233 | ~v_232 | ~v_405 | ~v_404 | ~v_597 | ~v_596 | ~v_1302 | ~v_1301 | ~v_1300 | ~v_1299 | ~v_1298 | ~v_1297 | ~v_1296 | ~v_1295 | ~v_1294 | ~v_1293 | ~v_225 | ~v_224 | ~v_223 | ~v_222 | ~v_221 | ~v_220 | ~v_401 | ~v_400 | ~v_399 | ~v_398 | ~v_4364 | ~v_4363 | ~v_4362 | ~v_4361 | v_4413;
assign x_278 = v_4412 | ~v_4409;
assign x_279 = v_4412 | ~v_4410;
assign x_280 = v_4412 | ~v_4411;
assign x_281 = v_101 | v_100 | v_99 | v_92 | v_102 | v_172 | v_171 | v_170 | v_169 | v_149 | v_148 | v_147 | ~v_483 | ~v_482 | ~v_593 | ~v_592 | ~v_545 | ~v_591 | ~v_590 | ~v_544 | ~v_1464 | ~v_1463 | ~v_1350 | ~v_1462 | ~v_1461 | ~v_1347 | ~v_1496 | ~v_1495 | ~v_1494 | ~v_1493 | ~v_477 | ~v_476 | ~v_289 | ~v_475 | ~v_474 | ~v_286 | ~v_539 | ~v_538 | ~v_537 | ~v_536 | ~v_4374 | ~v_4373 | ~v_4372 | ~v_4371 | v_4411;
assign x_282 = v_50 | v_60 | v_59 | v_58 | v_57 | v_144 | v_143 | v_142 | v_168 | v_167 | v_166 | v_165 | ~v_468 | ~v_467 | ~v_588 | ~v_587 | ~v_530 | ~v_586 | ~v_585 | ~v_529 | ~v_1455 | ~v_1454 | ~v_1325 | ~v_1453 | ~v_1452 | ~v_1322 | ~v_1487 | ~v_1486 | ~v_1485 | ~v_1484 | ~v_462 | ~v_461 | ~v_256 | ~v_460 | ~v_459 | ~v_253 | ~v_524 | ~v_523 | ~v_522 | ~v_521 | ~v_4369 | ~v_4368 | ~v_4367 | ~v_4366 | v_4410;
assign x_283 = v_7 | v_17 | v_16 | v_15 | v_14 | ~v_453 | ~v_452 | v_136 | v_135 | v_134 | v_164 | v_163 | v_162 | v_161 | ~v_583 | ~v_582 | ~v_515 | ~v_581 | ~v_580 | ~v_514 | ~v_1446 | ~v_1445 | ~v_1300 | ~v_1444 | ~v_1443 | ~v_1297 | ~v_1478 | ~v_1477 | ~v_1476 | ~v_1475 | ~v_447 | ~v_446 | ~v_223 | ~v_445 | ~v_444 | ~v_220 | ~v_509 | ~v_508 | ~v_507 | ~v_506 | ~v_4364 | ~v_4363 | ~v_4362 | ~v_4361 | v_4409;
assign x_284 = v_4408 | ~v_4405;
assign x_285 = v_4408 | ~v_4406;
assign x_286 = v_4408 | ~v_4407;
assign x_287 = v_103 | v_101 | v_97 | v_96 | v_100 | v_92 | v_151 | v_171 | v_170 | v_169 | v_150 | v_147 | ~v_577 | ~v_576 | ~v_545 | ~v_544 | ~v_575 | ~v_574 | ~v_435 | ~v_434 | ~v_1350 | ~v_1347 | ~v_1346 | ~v_1345 | ~v_1344 | ~v_1343 | ~v_1496 | ~v_1495 | ~v_1494 | ~v_1493 | ~v_289 | ~v_286 | ~v_431 | ~v_430 | ~v_429 | ~v_428 | ~v_539 | ~v_538 | ~v_537 | ~v_536 | ~v_4374 | ~v_4373 | ~v_4372 | ~v_4371 | v_4407;
assign x_288 = v_54 | v_55 | v_61 | v_50 | v_59 | v_58 | v_145 | v_142 | v_167 | v_166 | v_165 | v_146 | ~v_572 | ~v_571 | ~v_530 | ~v_529 | ~v_570 | ~v_569 | ~v_420 | ~v_419 | ~v_1325 | ~v_1322 | ~v_1321 | ~v_1320 | ~v_1319 | ~v_1318 | ~v_1487 | ~v_1486 | ~v_1485 | ~v_1484 | ~v_256 | ~v_253 | ~v_416 | ~v_415 | ~v_414 | ~v_413 | ~v_524 | ~v_523 | ~v_522 | ~v_521 | ~v_4369 | ~v_4368 | ~v_4367 | ~v_4366 | v_4406;
assign x_289 = v_7 | v_18 | v_16 | v_15 | v_12 | v_11 | v_134 | v_137 | v_138 | v_163 | v_162 | v_161 | ~v_567 | ~v_566 | ~v_515 | ~v_514 | ~v_565 | ~v_564 | ~v_405 | ~v_404 | ~v_1300 | ~v_1297 | ~v_1296 | ~v_1295 | ~v_1294 | ~v_1293 | ~v_1478 | ~v_1477 | ~v_1476 | ~v_1475 | ~v_223 | ~v_220 | ~v_401 | ~v_400 | ~v_399 | ~v_398 | ~v_509 | ~v_508 | ~v_507 | ~v_506 | ~v_4364 | ~v_4363 | ~v_4362 | ~v_4361 | v_4405;
assign x_290 = v_4404 | ~v_4401;
assign x_291 = v_4404 | ~v_4402;
assign x_292 = v_4404 | ~v_4403;
assign x_293 = v_103 | v_101 | v_100 | v_95 | v_92 | v_102 | v_171 | v_170 | v_169 | v_150 | v_149 | v_148 | ~v_545 | ~v_544 | ~v_561 | ~v_560 | ~v_559 | ~v_558 | ~v_387 | ~v_386 | ~v_1350 | ~v_1347 | ~v_1408 | ~v_1407 | ~v_1406 | ~v_1405 | ~v_1496 | ~v_1495 | ~v_1494 | ~v_1493 | ~v_289 | ~v_286 | ~v_383 | ~v_382 | ~v_381 | ~v_380 | ~v_539 | ~v_538 | ~v_537 | ~v_536 | ~v_4374 | ~v_4373 | ~v_4372 | ~v_4371 | v_4403;
assign x_294 = v_53 | v_61 | v_50 | v_60 | v_59 | v_58 | v_144 | v_145 | v_143 | v_167 | v_166 | v_165 | ~v_530 | ~v_529 | ~v_556 | ~v_555 | ~v_554 | ~v_553 | ~v_372 | ~v_371 | ~v_1325 | ~v_1322 | ~v_1399 | ~v_1398 | ~v_1397 | ~v_1396 | ~v_1487 | ~v_1486 | ~v_1485 | ~v_1484 | ~v_256 | ~v_253 | ~v_368 | ~v_367 | ~v_366 | ~v_365 | ~v_524 | ~v_523 | ~v_522 | ~v_521 | ~v_4369 | ~v_4368 | ~v_4367 | ~v_4366 | v_4402;
assign x_295 = v_7 | v_18 | v_17 | v_16 | v_15 | v_10 | v_136 | v_135 | v_137 | v_163 | v_162 | v_161 | ~v_515 | ~v_514 | ~v_551 | ~v_550 | ~v_549 | ~v_548 | ~v_357 | ~v_356 | ~v_1300 | ~v_1297 | ~v_1390 | ~v_1389 | ~v_1388 | ~v_1387 | ~v_1478 | ~v_1477 | ~v_1476 | ~v_1475 | ~v_223 | ~v_220 | ~v_353 | ~v_352 | ~v_351 | ~v_350 | ~v_509 | ~v_508 | ~v_507 | ~v_506 | ~v_4364 | ~v_4363 | ~v_4362 | ~v_4361 | v_4401;
assign x_296 = v_4400 | ~v_4397;
assign x_297 = v_4400 | ~v_4398;
assign x_298 = v_4400 | ~v_4399;
assign x_299 = v_103 | v_100 | v_92 | v_102 | v_171 | v_170 | v_169 | v_160 | v_150 | v_149 | v_148 | v_147 | ~v_545 | ~v_544 | ~v_543 | ~v_542 | ~v_541 | ~v_540 | ~v_297 | ~v_296 | ~v_1350 | ~v_1347 | ~v_1436 | ~v_1435 | ~v_1434 | ~v_1433 | ~v_1496 | ~v_1495 | ~v_1494 | ~v_1493 | ~v_289 | ~v_286 | ~v_285 | ~v_284 | ~v_283 | ~v_282 | ~v_539 | ~v_538 | ~v_537 | ~v_536 | ~v_4374 | ~v_4373 | ~v_4372 | ~v_4371 | v_4399;
assign x_300 = v_61 | v_50 | v_60 | v_58 | v_144 | v_159 | v_145 | v_143 | v_142 | v_167 | v_166 | v_165 | ~v_530 | ~v_529 | ~v_528 | ~v_527 | ~v_526 | ~v_525 | ~v_264 | ~v_263 | ~v_1325 | ~v_1322 | ~v_1427 | ~v_1426 | ~v_1425 | ~v_1424 | ~v_1487 | ~v_1486 | ~v_1485 | ~v_1484 | ~v_256 | ~v_253 | ~v_252 | ~v_251 | ~v_250 | ~v_249 | ~v_524 | ~v_523 | ~v_522 | ~v_521 | ~v_4369 | ~v_4368 | ~v_4367 | ~v_4366 | v_4398;
assign x_301 = v_7 | v_18 | v_17 | v_15 | v_136 | v_135 | v_134 | v_137 | v_163 | v_162 | v_161 | v_155 | ~v_515 | ~v_514 | ~v_513 | ~v_512 | ~v_511 | ~v_510 | ~v_231 | ~v_230 | ~v_1300 | ~v_1297 | ~v_1418 | ~v_1417 | ~v_1416 | ~v_1415 | ~v_1478 | ~v_1477 | ~v_1476 | ~v_1475 | ~v_223 | ~v_220 | ~v_219 | ~v_218 | ~v_217 | ~v_216 | ~v_509 | ~v_508 | ~v_507 | ~v_506 | ~v_4364 | ~v_4363 | ~v_4362 | ~v_4361 | v_4397;
assign x_302 = v_4396 | ~v_4393;
assign x_303 = v_4396 | ~v_4394;
assign x_304 = v_4396 | ~v_4395;
assign x_305 = v_98 | v_103 | v_101 | v_100 | v_92 | v_151 | v_170 | v_169 | v_150 | v_149 | v_148 | v_147 | ~v_299 | ~v_298 | ~v_387 | ~v_386 | ~v_499 | ~v_498 | ~v_497 | ~v_496 | ~v_1352 | ~v_1351 | ~v_1350 | ~v_1349 | ~v_1348 | ~v_1347 | ~v_1408 | ~v_1407 | ~v_1406 | ~v_1405 | ~v_291 | ~v_290 | ~v_289 | ~v_288 | ~v_287 | ~v_286 | ~v_383 | ~v_382 | ~v_381 | ~v_380 | ~v_4374 | ~v_4373 | ~v_4372 | ~v_4371 | v_4395;
assign x_306 = v_56 | v_61 | v_50 | v_59 | v_58 | v_144 | v_145 | v_143 | v_142 | v_166 | v_165 | v_146 | ~v_266 | ~v_265 | ~v_372 | ~v_371 | ~v_494 | ~v_493 | ~v_492 | ~v_491 | ~v_1327 | ~v_1326 | ~v_1325 | ~v_1324 | ~v_1323 | ~v_1322 | ~v_1399 | ~v_1398 | ~v_1397 | ~v_1396 | ~v_258 | ~v_257 | ~v_256 | ~v_255 | ~v_254 | ~v_253 | ~v_368 | ~v_367 | ~v_366 | ~v_365 | ~v_4369 | ~v_4368 | ~v_4367 | ~v_4366 | v_4394;
assign x_307 = v_13 | v_7 | v_18 | v_16 | v_15 | v_136 | v_135 | v_134 | v_137 | v_138 | v_162 | v_161 | ~v_233 | ~v_232 | ~v_357 | ~v_356 | ~v_489 | ~v_488 | ~v_487 | ~v_486 | ~v_1302 | ~v_1301 | ~v_1300 | ~v_1299 | ~v_1298 | ~v_1297 | ~v_1390 | ~v_1389 | ~v_1388 | ~v_1387 | ~v_225 | ~v_224 | ~v_223 | ~v_222 | ~v_221 | ~v_220 | ~v_353 | ~v_352 | ~v_351 | ~v_350 | ~v_4364 | ~v_4363 | ~v_4362 | ~v_4361 | v_4393;
assign x_308 = v_4392 | ~v_4389;
assign x_309 = v_4392 | ~v_4390;
assign x_310 = v_4392 | ~v_4391;
assign x_311 = v_103 | v_101 | v_99 | v_92 | v_102 | v_171 | v_170 | v_169 | v_149 | v_148 | v_147 | v_181 | ~v_483 | ~v_482 | ~v_481 | ~v_480 | ~v_345 | ~v_479 | ~v_478 | ~v_344 | ~v_1464 | ~v_1463 | ~v_1350 | ~v_1462 | ~v_1461 | ~v_1347 | ~v_1540 | ~v_1539 | ~v_1538 | ~v_1537 | ~v_477 | ~v_476 | ~v_289 | ~v_475 | ~v_474 | ~v_286 | ~v_339 | ~v_338 | ~v_337 | ~v_336 | ~v_4374 | ~v_4373 | ~v_4372 | ~v_4371 | v_4391;
assign x_312 = v_61 | v_50 | v_60 | v_59 | v_57 | v_144 | v_180 | v_143 | v_142 | v_167 | v_166 | v_165 | ~v_468 | ~v_467 | ~v_466 | ~v_465 | ~v_330 | ~v_464 | ~v_463 | ~v_329 | ~v_1455 | ~v_1454 | ~v_1325 | ~v_1453 | ~v_1452 | ~v_1322 | ~v_1531 | ~v_1530 | ~v_1529 | ~v_1528 | ~v_462 | ~v_461 | ~v_256 | ~v_460 | ~v_459 | ~v_253 | ~v_324 | ~v_323 | ~v_322 | ~v_321 | ~v_4369 | ~v_4368 | ~v_4367 | ~v_4366 | v_4390;
assign x_313 = v_7 | v_18 | v_17 | v_16 | v_14 | ~v_453 | ~v_452 | v_136 | v_135 | v_134 | v_179 | v_163 | v_162 | v_161 | ~v_451 | ~v_450 | ~v_315 | ~v_449 | ~v_448 | ~v_314 | ~v_1446 | ~v_1445 | ~v_1300 | ~v_1444 | ~v_1443 | ~v_1297 | ~v_1522 | ~v_1521 | ~v_1520 | ~v_1519 | ~v_447 | ~v_446 | ~v_223 | ~v_445 | ~v_444 | ~v_220 | ~v_309 | ~v_308 | ~v_307 | ~v_306 | ~v_4364 | ~v_4363 | ~v_4362 | ~v_4361 | v_4389;
assign x_314 = v_4388 | ~v_4385;
assign x_315 = v_4388 | ~v_4386;
assign x_316 = v_4388 | ~v_4387;
assign x_317 = v_101 | v_97 | v_96 | v_92 | v_102 | v_172 | v_171 | v_170 | v_169 | v_150 | v_147 | v_181 | ~v_437 | ~v_436 | ~v_435 | ~v_434 | ~v_345 | ~v_344 | ~v_433 | ~v_432 | ~v_1350 | ~v_1347 | ~v_1346 | ~v_1345 | ~v_1344 | ~v_1343 | ~v_1540 | ~v_1539 | ~v_1538 | ~v_1537 | ~v_289 | ~v_286 | ~v_431 | ~v_430 | ~v_429 | ~v_428 | ~v_339 | ~v_338 | ~v_337 | ~v_336 | ~v_4374 | ~v_4373 | ~v_4372 | ~v_4371 | v_4387;
assign x_318 = v_54 | v_55 | v_50 | v_60 | v_59 | v_180 | v_145 | v_142 | v_168 | v_167 | v_166 | v_165 | ~v_422 | ~v_421 | ~v_420 | ~v_419 | ~v_330 | ~v_329 | ~v_418 | ~v_417 | ~v_1325 | ~v_1322 | ~v_1321 | ~v_1320 | ~v_1319 | ~v_1318 | ~v_1531 | ~v_1530 | ~v_1529 | ~v_1528 | ~v_256 | ~v_253 | ~v_416 | ~v_415 | ~v_414 | ~v_413 | ~v_324 | ~v_323 | ~v_322 | ~v_321 | ~v_4369 | ~v_4368 | ~v_4367 | ~v_4366 | v_4386;
assign x_319 = v_7 | v_17 | v_16 | v_12 | v_11 | v_134 | v_137 | v_179 | v_164 | v_163 | v_162 | v_161 | ~v_407 | ~v_406 | ~v_405 | ~v_404 | ~v_315 | ~v_314 | ~v_403 | ~v_402 | ~v_1300 | ~v_1297 | ~v_1296 | ~v_1295 | ~v_1294 | ~v_1293 | ~v_1522 | ~v_1521 | ~v_1520 | ~v_1519 | ~v_223 | ~v_220 | ~v_401 | ~v_400 | ~v_399 | ~v_398 | ~v_309 | ~v_308 | ~v_307 | ~v_306 | ~v_4364 | ~v_4363 | ~v_4362 | ~v_4361 | v_4385;
assign x_320 = v_4384 | ~v_4381;
assign x_321 = v_4384 | ~v_4382;
assign x_322 = v_4384 | ~v_4383;
assign x_323 = v_103 | v_101 | v_92 | v_102 | v_171 | v_170 | v_169 | v_150 | v_149 | v_148 | v_147 | v_181 | ~v_391 | ~v_390 | ~v_387 | ~v_386 | ~v_345 | ~v_344 | ~v_385 | ~v_384 | ~v_1350 | ~v_1347 | ~v_1408 | ~v_1407 | ~v_1406 | ~v_1405 | ~v_1540 | ~v_1539 | ~v_1538 | ~v_1537 | ~v_289 | ~v_286 | ~v_383 | ~v_382 | ~v_381 | ~v_380 | ~v_339 | ~v_338 | ~v_337 | ~v_336 | ~v_4374 | ~v_4373 | ~v_4372 | ~v_4371 | v_4383;
assign x_324 = v_61 | v_50 | v_60 | v_59 | v_144 | v_180 | v_145 | v_143 | v_142 | v_167 | v_166 | v_165 | ~v_376 | ~v_375 | ~v_372 | ~v_371 | ~v_330 | ~v_329 | ~v_370 | ~v_369 | ~v_1325 | ~v_1322 | ~v_1399 | ~v_1398 | ~v_1397 | ~v_1396 | ~v_1531 | ~v_1530 | ~v_1529 | ~v_1528 | ~v_256 | ~v_253 | ~v_368 | ~v_367 | ~v_366 | ~v_365 | ~v_324 | ~v_323 | ~v_322 | ~v_321 | ~v_4369 | ~v_4368 | ~v_4367 | ~v_4366 | v_4382;
assign x_325 = v_7 | v_18 | v_17 | v_16 | v_136 | v_135 | v_134 | v_137 | v_179 | v_163 | v_162 | v_161 | ~v_361 | ~v_360 | ~v_357 | ~v_356 | ~v_315 | ~v_314 | ~v_355 | ~v_354 | ~v_1300 | ~v_1297 | ~v_1390 | ~v_1389 | ~v_1388 | ~v_1387 | ~v_1522 | ~v_1521 | ~v_1520 | ~v_1519 | ~v_223 | ~v_220 | ~v_353 | ~v_352 | ~v_351 | ~v_350 | ~v_309 | ~v_308 | ~v_307 | ~v_306 | ~v_4364 | ~v_4363 | ~v_4362 | ~v_4361 | v_4381;
assign x_326 = v_4380 | ~v_4377;
assign x_327 = v_4380 | ~v_4378;
assign x_328 = v_4380 | ~v_4379;
assign x_329 = v_103 | v_95 | v_92 | v_102 | v_171 | v_170 | v_169 | v_160 | v_150 | v_149 | v_148 | v_181 | ~v_297 | ~v_296 | ~v_345 | ~v_344 | ~v_343 | ~v_342 | ~v_341 | ~v_340 | ~v_1350 | ~v_1347 | ~v_1436 | ~v_1435 | ~v_1434 | ~v_1433 | ~v_1540 | ~v_1539 | ~v_1538 | ~v_1537 | ~v_289 | ~v_286 | ~v_285 | ~v_284 | ~v_283 | ~v_282 | ~v_339 | ~v_338 | ~v_337 | ~v_336 | ~v_4374 | ~v_4373 | ~v_4372 | ~v_4371 | v_4379;
assign x_330 = v_53 | v_61 | v_50 | v_60 | v_144 | v_180 | v_159 | v_145 | v_143 | v_167 | v_166 | v_165 | ~v_264 | ~v_263 | ~v_330 | ~v_329 | ~v_328 | ~v_327 | ~v_326 | ~v_325 | ~v_1325 | ~v_1322 | ~v_1427 | ~v_1426 | ~v_1425 | ~v_1424 | ~v_1531 | ~v_1530 | ~v_1529 | ~v_1528 | ~v_256 | ~v_253 | ~v_252 | ~v_251 | ~v_250 | ~v_249 | ~v_324 | ~v_323 | ~v_322 | ~v_321 | ~v_4369 | ~v_4368 | ~v_4367 | ~v_4366 | v_4378;
assign x_331 = v_7 | v_18 | v_17 | v_10 | v_136 | v_135 | v_137 | v_179 | v_163 | v_162 | v_161 | v_155 | ~v_231 | ~v_230 | ~v_315 | ~v_314 | ~v_313 | ~v_312 | ~v_311 | ~v_310 | ~v_1300 | ~v_1297 | ~v_1418 | ~v_1417 | ~v_1416 | ~v_1415 | ~v_1522 | ~v_1521 | ~v_1520 | ~v_1519 | ~v_223 | ~v_220 | ~v_219 | ~v_218 | ~v_217 | ~v_216 | ~v_309 | ~v_308 | ~v_307 | ~v_306 | ~v_4364 | ~v_4363 | ~v_4362 | ~v_4361 | v_4377;
assign x_332 = v_4376 | ~v_4365;
assign x_333 = v_4376 | ~v_4370;
assign x_334 = v_4376 | ~v_4375;
assign x_335 = v_98 | v_103 | v_100 | v_92 | v_102 | v_170 | v_169 | v_160 | v_150 | v_149 | v_148 | v_147 | ~v_299 | ~v_298 | ~v_297 | ~v_296 | ~v_295 | ~v_294 | ~v_293 | ~v_292 | ~v_1352 | ~v_1351 | ~v_1350 | ~v_1349 | ~v_1348 | ~v_1347 | ~v_1436 | ~v_1435 | ~v_1434 | ~v_1433 | ~v_291 | ~v_290 | ~v_289 | ~v_288 | ~v_287 | ~v_286 | ~v_285 | ~v_284 | ~v_283 | ~v_282 | ~v_4374 | ~v_4373 | ~v_4372 | ~v_4371 | v_4375;
assign x_336 = v_4374 | v_154;
assign x_337 = v_4374 | v_123;
assign x_338 = v_4373 | v_154;
assign x_339 = v_4373 | v_120;
assign x_340 = v_4372 | ~v_154;
assign x_341 = v_4372 | v_108;
assign x_342 = v_4371 | ~v_154;
assign x_343 = v_4371 | v_105;
assign x_344 = v_56 | v_61 | v_50 | v_60 | v_58 | v_144 | v_159 | v_145 | v_143 | v_142 | v_166 | v_165 | ~v_266 | ~v_265 | ~v_264 | ~v_263 | ~v_262 | ~v_261 | ~v_260 | ~v_259 | ~v_1327 | ~v_1326 | ~v_1325 | ~v_1324 | ~v_1323 | ~v_1322 | ~v_1427 | ~v_1426 | ~v_1425 | ~v_1424 | ~v_258 | ~v_257 | ~v_256 | ~v_255 | ~v_254 | ~v_253 | ~v_252 | ~v_251 | ~v_250 | ~v_249 | ~v_4369 | ~v_4368 | ~v_4367 | ~v_4366 | v_4370;
assign x_345 = v_4369 | v_154;
assign x_346 = v_4369 | v_81;
assign x_347 = v_4368 | v_154;
assign x_348 = v_4368 | v_78;
assign x_349 = v_4367 | ~v_154;
assign x_350 = v_4367 | v_66;
assign x_351 = v_4366 | ~v_154;
assign x_352 = v_4366 | v_63;
assign x_353 = v_13 | v_7 | v_18 | v_17 | v_15 | v_136 | v_135 | v_134 | v_137 | v_162 | v_161 | v_155 | ~v_233 | ~v_232 | ~v_231 | ~v_230 | ~v_229 | ~v_228 | ~v_227 | ~v_226 | ~v_1302 | ~v_1301 | ~v_1300 | ~v_1299 | ~v_1298 | ~v_1297 | ~v_1418 | ~v_1417 | ~v_1416 | ~v_1415 | ~v_225 | ~v_224 | ~v_223 | ~v_222 | ~v_221 | ~v_220 | ~v_219 | ~v_218 | ~v_217 | ~v_216 | ~v_4364 | ~v_4363 | ~v_4362 | ~v_4361 | v_4365;
assign x_354 = v_4364 | v_154;
assign x_355 = v_4364 | v_39;
assign x_356 = v_4363 | v_154;
assign x_357 = v_4363 | v_36;
assign x_358 = v_4362 | ~v_154;
assign x_359 = v_4362 | v_24;
assign x_360 = v_4361 | ~v_154;
assign x_361 = v_4361 | v_21;
assign x_362 = v_4360 | ~v_4357;
assign x_363 = v_4360 | ~v_4358;
assign x_364 = v_4360 | ~v_4359;
assign x_365 = v_98 | v_103 | v_101 | v_100 | v_95 | v_99 | v_92 | v_102 | ~v_719 | ~v_718 | v_170 | v_169 | v_149 | v_148 | ~v_483 | ~v_717 | ~v_299 | ~v_482 | ~v_716 | ~v_298 | ~v_473 | ~v_281 | ~v_472 | ~v_280 | ~v_279 | ~v_471 | ~v_278 | ~v_470 | ~v_277 | ~v_276 | ~v_1460 | ~v_1342 | ~v_1459 | ~v_1341 | ~v_1340 | ~v_1458 | ~v_1339 | ~v_1457 | ~v_1338 | ~v_1337 | ~v_4298 | ~v_4297 | ~v_4296 | ~v_4295 | v_4359;
assign x_366 = v_53 | v_56 | v_61 | v_50 | v_60 | v_59 | v_58 | v_57 | ~v_714 | ~v_713 | v_144 | v_143 | v_166 | v_165 | ~v_266 | ~v_468 | ~v_712 | ~v_467 | ~v_711 | ~v_265 | ~v_458 | ~v_248 | ~v_457 | ~v_247 | ~v_246 | ~v_456 | ~v_245 | ~v_455 | ~v_244 | ~v_243 | ~v_1451 | ~v_1317 | ~v_1450 | ~v_1316 | ~v_1315 | ~v_1449 | ~v_1314 | ~v_1448 | ~v_1313 | ~v_1312 | ~v_4293 | ~v_4292 | ~v_4291 | ~v_4290 | v_4358;
assign x_367 = v_13 | v_7 | v_18 | v_17 | v_16 | v_15 | v_14 | v_10 | ~v_453 | ~v_709 | ~v_452 | ~v_708 | v_136 | v_135 | ~v_707 | ~v_706 | v_162 | v_161 | ~v_233 | ~v_232 | ~v_443 | ~v_215 | ~v_442 | ~v_214 | ~v_213 | ~v_441 | ~v_212 | ~v_440 | ~v_211 | ~v_210 | ~v_1442 | ~v_1292 | ~v_1441 | ~v_1291 | ~v_1290 | ~v_1440 | ~v_1289 | ~v_1439 | ~v_1288 | ~v_1287 | ~v_4288 | ~v_4287 | ~v_4286 | ~v_4285 | v_4357;
assign x_368 = v_4356 | ~v_4353;
assign x_369 = v_4356 | ~v_4354;
assign x_370 = v_4356 | ~v_4355;
assign x_371 = v_103 | v_101 | v_94 | v_99 | v_93 | v_92 | v_102 | v_171 | v_149 | v_148 | v_147 | v_181 | ~v_483 | ~v_482 | ~v_481 | ~v_480 | ~v_345 | ~v_479 | ~v_478 | ~v_344 | ~v_473 | ~v_472 | ~v_279 | ~v_471 | ~v_470 | ~v_276 | ~v_335 | ~v_334 | ~v_333 | ~v_332 | ~v_1460 | ~v_1459 | ~v_1340 | ~v_1458 | ~v_1457 | ~v_1337 | ~v_1536 | ~v_1535 | ~v_1534 | ~v_1533 | ~v_4298 | ~v_4297 | ~v_4296 | ~v_4295 | v_4355;
assign x_372 = v_61 | v_52 | v_50 | v_51 | v_60 | v_59 | v_57 | v_144 | v_180 | v_143 | v_142 | v_167 | ~v_468 | ~v_467 | ~v_466 | ~v_465 | ~v_330 | ~v_464 | ~v_463 | ~v_329 | ~v_458 | ~v_457 | ~v_246 | ~v_456 | ~v_455 | ~v_243 | ~v_320 | ~v_319 | ~v_318 | ~v_317 | ~v_1451 | ~v_1450 | ~v_1315 | ~v_1449 | ~v_1448 | ~v_1312 | ~v_1527 | ~v_1526 | ~v_1525 | ~v_1524 | ~v_4293 | ~v_4292 | ~v_4291 | ~v_4290 | v_4354;
assign x_373 = v_9 | v_7 | v_18 | v_17 | v_16 | v_8 | v_14 | ~v_453 | ~v_452 | v_136 | v_135 | v_134 | v_179 | v_163 | ~v_451 | ~v_450 | ~v_315 | ~v_449 | ~v_448 | ~v_314 | ~v_443 | ~v_442 | ~v_213 | ~v_441 | ~v_440 | ~v_210 | ~v_305 | ~v_304 | ~v_303 | ~v_302 | ~v_1442 | ~v_1441 | ~v_1290 | ~v_1440 | ~v_1439 | ~v_1287 | ~v_1518 | ~v_1517 | ~v_1516 | ~v_1515 | ~v_4288 | ~v_4287 | ~v_4286 | ~v_4285 | v_4353;
assign x_374 = v_4352 | ~v_4349;
assign x_375 = v_4352 | ~v_4350;
assign x_376 = v_4352 | ~v_4351;
assign x_377 = v_103 | v_97 | v_96 | v_95 | v_94 | v_93 | v_92 | v_102 | v_171 | v_160 | v_150 | v_181 | ~v_297 | ~v_296 | ~v_345 | ~v_344 | ~v_343 | ~v_342 | ~v_341 | ~v_340 | ~v_279 | ~v_276 | ~v_335 | ~v_334 | ~v_333 | ~v_332 | ~v_275 | ~v_274 | ~v_273 | ~v_272 | ~v_1340 | ~v_1337 | ~v_1536 | ~v_1535 | ~v_1534 | ~v_1533 | ~v_1432 | ~v_1431 | ~v_1430 | ~v_1429 | ~v_4298 | ~v_4297 | ~v_4296 | ~v_4295 | v_4351;
assign x_378 = v_54 | v_53 | v_55 | v_61 | v_52 | v_50 | v_51 | v_60 | v_180 | v_159 | v_145 | v_167 | ~v_264 | ~v_263 | ~v_330 | ~v_329 | ~v_328 | ~v_327 | ~v_326 | ~v_325 | ~v_246 | ~v_243 | ~v_320 | ~v_319 | ~v_318 | ~v_317 | ~v_242 | ~v_241 | ~v_240 | ~v_239 | ~v_1315 | ~v_1312 | ~v_1527 | ~v_1526 | ~v_1525 | ~v_1524 | ~v_1423 | ~v_1422 | ~v_1421 | ~v_1420 | ~v_4293 | ~v_4292 | ~v_4291 | ~v_4290 | v_4350;
assign x_379 = v_9 | v_7 | v_18 | v_17 | v_8 | v_12 | v_11 | v_10 | v_137 | v_179 | v_163 | v_155 | ~v_231 | ~v_230 | ~v_315 | ~v_314 | ~v_313 | ~v_312 | ~v_311 | ~v_310 | ~v_213 | ~v_210 | ~v_305 | ~v_304 | ~v_303 | ~v_302 | ~v_209 | ~v_208 | ~v_207 | ~v_206 | ~v_1290 | ~v_1287 | ~v_1518 | ~v_1517 | ~v_1516 | ~v_1515 | ~v_1414 | ~v_1413 | ~v_1412 | ~v_1411 | ~v_4288 | ~v_4287 | ~v_4286 | ~v_4285 | v_4349;
assign x_380 = v_4348 | ~v_4345;
assign x_381 = v_4348 | ~v_4346;
assign x_382 = v_4348 | ~v_4347;
assign x_383 = v_103 | v_101 | v_94 | v_93 | v_92 | v_102 | v_171 | v_150 | v_149 | v_148 | v_147 | v_181 | ~v_391 | ~v_390 | ~v_389 | ~v_388 | ~v_387 | ~v_386 | ~v_345 | ~v_344 | ~v_385 | ~v_384 | ~v_279 | ~v_276 | ~v_335 | ~v_334 | ~v_333 | ~v_332 | ~v_379 | ~v_378 | ~v_1340 | ~v_1337 | ~v_1536 | ~v_1535 | ~v_1534 | ~v_1533 | ~v_1404 | ~v_1403 | ~v_1402 | ~v_1401 | ~v_4298 | ~v_4297 | ~v_4296 | ~v_4295 | v_4347;
assign x_384 = v_61 | v_52 | v_50 | v_51 | v_60 | v_59 | v_144 | v_180 | v_145 | v_143 | v_142 | v_167 | ~v_376 | ~v_375 | ~v_374 | ~v_373 | ~v_372 | ~v_371 | ~v_330 | ~v_329 | ~v_370 | ~v_369 | ~v_246 | ~v_243 | ~v_320 | ~v_319 | ~v_318 | ~v_317 | ~v_364 | ~v_363 | ~v_1315 | ~v_1312 | ~v_1527 | ~v_1526 | ~v_1525 | ~v_1524 | ~v_1395 | ~v_1394 | ~v_1393 | ~v_1392 | ~v_4293 | ~v_4292 | ~v_4291 | ~v_4290 | v_4346;
assign x_385 = v_9 | v_7 | v_18 | v_17 | v_16 | v_8 | v_136 | v_135 | v_134 | v_137 | v_179 | v_163 | ~v_361 | ~v_360 | ~v_359 | ~v_358 | ~v_357 | ~v_356 | ~v_315 | ~v_314 | ~v_355 | ~v_354 | ~v_213 | ~v_210 | ~v_305 | ~v_304 | ~v_303 | ~v_302 | ~v_349 | ~v_348 | ~v_1290 | ~v_1287 | ~v_1518 | ~v_1517 | ~v_1516 | ~v_1515 | ~v_1386 | ~v_1385 | ~v_1384 | ~v_1383 | ~v_4288 | ~v_4287 | ~v_4286 | ~v_4285 | v_4345;
assign x_386 = v_4344 | ~v_4341;
assign x_387 = v_4344 | ~v_4342;
assign x_388 = v_4344 | ~v_4343;
assign x_389 = v_101 | v_94 | v_93 | v_92 | v_102 | v_172 | v_171 | v_150 | v_149 | v_148 | v_147 | v_181 | ~v_437 | ~v_436 | ~v_435 | ~v_434 | ~v_345 | ~v_344 | ~v_433 | ~v_432 | ~v_279 | ~v_276 | ~v_335 | ~v_334 | ~v_333 | ~v_332 | ~v_427 | ~v_426 | ~v_425 | ~v_424 | ~v_1340 | ~v_1337 | ~v_1536 | ~v_1535 | ~v_1534 | ~v_1533 | ~v_1336 | ~v_1335 | ~v_1334 | ~v_1333 | ~v_4298 | ~v_4297 | ~v_4296 | ~v_4295 | v_4343;
assign x_390 = v_52 | v_50 | v_51 | v_60 | v_59 | v_144 | v_180 | v_145 | v_143 | v_142 | v_168 | v_167 | ~v_422 | ~v_421 | ~v_420 | ~v_419 | ~v_330 | ~v_329 | ~v_418 | ~v_417 | ~v_246 | ~v_243 | ~v_320 | ~v_319 | ~v_318 | ~v_317 | ~v_412 | ~v_411 | ~v_410 | ~v_409 | ~v_1315 | ~v_1312 | ~v_1527 | ~v_1526 | ~v_1525 | ~v_1524 | ~v_1311 | ~v_1310 | ~v_1309 | ~v_1308 | ~v_4293 | ~v_4292 | ~v_4291 | ~v_4290 | v_4342;
assign x_391 = v_9 | v_7 | v_17 | v_16 | v_8 | v_136 | v_135 | v_134 | v_137 | v_179 | v_164 | v_163 | ~v_407 | ~v_406 | ~v_405 | ~v_404 | ~v_315 | ~v_314 | ~v_403 | ~v_402 | ~v_213 | ~v_210 | ~v_305 | ~v_304 | ~v_303 | ~v_302 | ~v_397 | ~v_396 | ~v_395 | ~v_394 | ~v_1290 | ~v_1287 | ~v_1518 | ~v_1517 | ~v_1516 | ~v_1515 | ~v_1286 | ~v_1285 | ~v_1284 | ~v_1283 | ~v_4288 | ~v_4287 | ~v_4286 | ~v_4285 | v_4341;
assign x_392 = v_4340 | ~v_4337;
assign x_393 = v_4340 | ~v_4338;
assign x_394 = v_4340 | ~v_4339;
assign x_395 = v_98 | v_103 | v_97 | v_96 | v_100 | v_92 | v_102 | v_170 | v_169 | v_160 | v_150 | v_147 | ~v_299 | ~v_298 | ~v_297 | ~v_296 | ~v_295 | ~v_294 | ~v_293 | ~v_292 | ~v_281 | ~v_280 | ~v_279 | ~v_278 | ~v_277 | ~v_276 | ~v_275 | ~v_274 | ~v_273 | ~v_272 | ~v_1342 | ~v_1341 | ~v_1340 | ~v_1339 | ~v_1338 | ~v_1337 | ~v_1432 | ~v_1431 | ~v_1430 | ~v_1429 | ~v_4298 | ~v_4297 | ~v_4296 | ~v_4295 | v_4339;
assign x_396 = v_54 | v_56 | v_55 | v_61 | v_50 | v_60 | v_58 | v_159 | v_145 | v_142 | v_166 | v_165 | ~v_266 | ~v_265 | ~v_264 | ~v_263 | ~v_262 | ~v_261 | ~v_260 | ~v_259 | ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_244 | ~v_243 | ~v_242 | ~v_241 | ~v_240 | ~v_239 | ~v_1317 | ~v_1316 | ~v_1315 | ~v_1314 | ~v_1313 | ~v_1312 | ~v_1423 | ~v_1422 | ~v_1421 | ~v_1420 | ~v_4293 | ~v_4292 | ~v_4291 | ~v_4290 | v_4338;
assign x_397 = v_13 | v_7 | v_18 | v_17 | v_15 | v_12 | v_11 | v_134 | v_137 | v_162 | v_161 | v_155 | ~v_233 | ~v_232 | ~v_231 | ~v_230 | ~v_229 | ~v_228 | ~v_227 | ~v_226 | ~v_215 | ~v_214 | ~v_213 | ~v_212 | ~v_211 | ~v_210 | ~v_209 | ~v_208 | ~v_207 | ~v_206 | ~v_1292 | ~v_1291 | ~v_1290 | ~v_1289 | ~v_1288 | ~v_1287 | ~v_1414 | ~v_1413 | ~v_1412 | ~v_1411 | ~v_4288 | ~v_4287 | ~v_4286 | ~v_4285 | v_4337;
assign x_398 = v_4336 | ~v_4333;
assign x_399 = v_4336 | ~v_4334;
assign x_400 = v_4336 | ~v_4335;
assign x_401 = v_101 | v_100 | v_99 | v_92 | v_102 | v_172 | v_171 | v_170 | v_169 | v_149 | v_148 | v_147 | ~v_483 | ~v_482 | ~v_593 | ~v_592 | ~v_545 | ~v_591 | ~v_590 | ~v_544 | ~v_473 | ~v_472 | ~v_279 | ~v_471 | ~v_470 | ~v_276 | ~v_535 | ~v_534 | ~v_533 | ~v_532 | ~v_1460 | ~v_1459 | ~v_1340 | ~v_1458 | ~v_1457 | ~v_1337 | ~v_1492 | ~v_1491 | ~v_1490 | ~v_1489 | ~v_4298 | ~v_4297 | ~v_4296 | ~v_4295 | v_4335;
assign x_402 = v_50 | v_60 | v_59 | v_58 | v_57 | v_144 | v_143 | v_142 | v_168 | v_167 | v_166 | v_165 | ~v_468 | ~v_467 | ~v_588 | ~v_587 | ~v_530 | ~v_586 | ~v_585 | ~v_529 | ~v_458 | ~v_457 | ~v_246 | ~v_456 | ~v_455 | ~v_243 | ~v_520 | ~v_519 | ~v_518 | ~v_517 | ~v_1451 | ~v_1450 | ~v_1315 | ~v_1449 | ~v_1448 | ~v_1312 | ~v_1483 | ~v_1482 | ~v_1481 | ~v_1480 | ~v_4293 | ~v_4292 | ~v_4291 | ~v_4290 | v_4334;
assign x_403 = v_7 | v_17 | v_16 | v_15 | v_14 | ~v_453 | ~v_452 | v_136 | v_135 | v_134 | v_164 | v_163 | v_162 | v_161 | ~v_583 | ~v_582 | ~v_515 | ~v_581 | ~v_580 | ~v_514 | ~v_443 | ~v_442 | ~v_213 | ~v_441 | ~v_440 | ~v_210 | ~v_505 | ~v_504 | ~v_503 | ~v_502 | ~v_1442 | ~v_1441 | ~v_1290 | ~v_1440 | ~v_1439 | ~v_1287 | ~v_1474 | ~v_1473 | ~v_1472 | ~v_1471 | ~v_4288 | ~v_4287 | ~v_4286 | ~v_4285 | v_4333;
assign x_404 = v_4332 | ~v_4329;
assign x_405 = v_4332 | ~v_4330;
assign x_406 = v_4332 | ~v_4331;
assign x_407 = v_103 | v_97 | v_96 | v_100 | v_92 | v_102 | v_171 | v_170 | v_169 | v_160 | v_150 | v_147 | ~v_545 | ~v_544 | ~v_543 | ~v_542 | ~v_541 | ~v_540 | ~v_297 | ~v_296 | ~v_279 | ~v_276 | ~v_275 | ~v_274 | ~v_273 | ~v_272 | ~v_535 | ~v_534 | ~v_533 | ~v_532 | ~v_1340 | ~v_1337 | ~v_1432 | ~v_1431 | ~v_1430 | ~v_1429 | ~v_1492 | ~v_1491 | ~v_1490 | ~v_1489 | ~v_4298 | ~v_4297 | ~v_4296 | ~v_4295 | v_4331;
assign x_408 = v_54 | v_55 | v_61 | v_50 | v_60 | v_58 | v_159 | v_145 | v_142 | v_167 | v_166 | v_165 | ~v_530 | ~v_529 | ~v_528 | ~v_527 | ~v_526 | ~v_525 | ~v_264 | ~v_263 | ~v_246 | ~v_243 | ~v_242 | ~v_241 | ~v_240 | ~v_239 | ~v_520 | ~v_519 | ~v_518 | ~v_517 | ~v_1315 | ~v_1312 | ~v_1423 | ~v_1422 | ~v_1421 | ~v_1420 | ~v_1483 | ~v_1482 | ~v_1481 | ~v_1480 | ~v_4293 | ~v_4292 | ~v_4291 | ~v_4290 | v_4330;
assign x_409 = v_7 | v_18 | v_17 | v_15 | v_12 | v_11 | v_134 | v_137 | v_163 | v_162 | v_161 | v_155 | ~v_515 | ~v_514 | ~v_513 | ~v_512 | ~v_511 | ~v_510 | ~v_231 | ~v_230 | ~v_213 | ~v_210 | ~v_209 | ~v_208 | ~v_207 | ~v_206 | ~v_505 | ~v_504 | ~v_503 | ~v_502 | ~v_1290 | ~v_1287 | ~v_1414 | ~v_1413 | ~v_1412 | ~v_1411 | ~v_1474 | ~v_1473 | ~v_1472 | ~v_1471 | ~v_4288 | ~v_4287 | ~v_4286 | ~v_4285 | v_4329;
assign x_410 = v_4328 | ~v_4325;
assign x_411 = v_4328 | ~v_4326;
assign x_412 = v_4328 | ~v_4327;
assign x_413 = v_103 | v_101 | v_100 | v_95 | v_92 | v_102 | v_171 | v_170 | v_169 | v_150 | v_149 | v_148 | ~v_389 | ~v_388 | ~v_545 | ~v_544 | ~v_561 | ~v_560 | ~v_559 | ~v_558 | ~v_387 | ~v_386 | ~v_279 | ~v_276 | ~v_379 | ~v_378 | ~v_535 | ~v_534 | ~v_533 | ~v_532 | ~v_1340 | ~v_1337 | ~v_1404 | ~v_1403 | ~v_1402 | ~v_1401 | ~v_1492 | ~v_1491 | ~v_1490 | ~v_1489 | ~v_4298 | ~v_4297 | ~v_4296 | ~v_4295 | v_4327;
assign x_414 = v_53 | v_61 | v_50 | v_60 | v_59 | v_58 | v_144 | v_145 | v_143 | v_167 | v_166 | v_165 | ~v_374 | ~v_373 | ~v_530 | ~v_529 | ~v_556 | ~v_555 | ~v_554 | ~v_553 | ~v_372 | ~v_371 | ~v_246 | ~v_243 | ~v_364 | ~v_363 | ~v_520 | ~v_519 | ~v_518 | ~v_517 | ~v_1315 | ~v_1312 | ~v_1395 | ~v_1394 | ~v_1393 | ~v_1392 | ~v_1483 | ~v_1482 | ~v_1481 | ~v_1480 | ~v_4293 | ~v_4292 | ~v_4291 | ~v_4290 | v_4326;
assign x_415 = v_7 | v_18 | v_17 | v_16 | v_15 | v_10 | v_136 | v_135 | v_137 | v_163 | v_162 | v_161 | ~v_359 | ~v_358 | ~v_515 | ~v_514 | ~v_551 | ~v_550 | ~v_549 | ~v_548 | ~v_357 | ~v_356 | ~v_213 | ~v_210 | ~v_349 | ~v_348 | ~v_505 | ~v_504 | ~v_503 | ~v_502 | ~v_1290 | ~v_1287 | ~v_1386 | ~v_1385 | ~v_1384 | ~v_1383 | ~v_1474 | ~v_1473 | ~v_1472 | ~v_1471 | ~v_4288 | ~v_4287 | ~v_4286 | ~v_4285 | v_4325;
assign x_416 = v_4324 | ~v_4321;
assign x_417 = v_4324 | ~v_4322;
assign x_418 = v_4324 | ~v_4323;
assign x_419 = v_103 | v_101 | v_100 | v_92 | v_151 | v_171 | v_170 | v_169 | v_150 | v_149 | v_148 | v_147 | ~v_577 | ~v_576 | ~v_545 | ~v_544 | ~v_575 | ~v_574 | ~v_435 | ~v_434 | ~v_279 | ~v_276 | ~v_427 | ~v_426 | ~v_425 | ~v_424 | ~v_535 | ~v_534 | ~v_533 | ~v_532 | ~v_1340 | ~v_1337 | ~v_1336 | ~v_1335 | ~v_1334 | ~v_1333 | ~v_1492 | ~v_1491 | ~v_1490 | ~v_1489 | ~v_4298 | ~v_4297 | ~v_4296 | ~v_4295 | v_4323;
assign x_420 = v_61 | v_50 | v_59 | v_58 | v_144 | v_145 | v_143 | v_142 | v_167 | v_166 | v_165 | v_146 | ~v_572 | ~v_571 | ~v_530 | ~v_529 | ~v_570 | ~v_569 | ~v_420 | ~v_419 | ~v_246 | ~v_243 | ~v_412 | ~v_411 | ~v_410 | ~v_409 | ~v_520 | ~v_519 | ~v_518 | ~v_517 | ~v_1315 | ~v_1312 | ~v_1311 | ~v_1310 | ~v_1309 | ~v_1308 | ~v_1483 | ~v_1482 | ~v_1481 | ~v_1480 | ~v_4293 | ~v_4292 | ~v_4291 | ~v_4290 | v_4322;
assign x_421 = v_7 | v_18 | v_16 | v_15 | v_136 | v_135 | v_134 | v_137 | v_138 | v_163 | v_162 | v_161 | ~v_567 | ~v_566 | ~v_515 | ~v_514 | ~v_565 | ~v_564 | ~v_405 | ~v_404 | ~v_213 | ~v_210 | ~v_397 | ~v_396 | ~v_395 | ~v_394 | ~v_505 | ~v_504 | ~v_503 | ~v_502 | ~v_1290 | ~v_1287 | ~v_1286 | ~v_1285 | ~v_1284 | ~v_1283 | ~v_1474 | ~v_1473 | ~v_1472 | ~v_1471 | ~v_4288 | ~v_4287 | ~v_4286 | ~v_4285 | v_4321;
assign x_422 = v_4320 | ~v_4317;
assign x_423 = v_4320 | ~v_4318;
assign x_424 = v_4320 | ~v_4319;
assign x_425 = v_98 | v_103 | v_101 | v_100 | v_92 | v_151 | v_170 | v_169 | v_150 | v_149 | v_148 | v_147 | ~v_389 | ~v_388 | ~v_299 | ~v_298 | ~v_387 | ~v_386 | ~v_499 | ~v_498 | ~v_497 | ~v_496 | ~v_281 | ~v_280 | ~v_279 | ~v_278 | ~v_277 | ~v_276 | ~v_379 | ~v_378 | ~v_1342 | ~v_1341 | ~v_1340 | ~v_1339 | ~v_1338 | ~v_1337 | ~v_1404 | ~v_1403 | ~v_1402 | ~v_1401 | ~v_4298 | ~v_4297 | ~v_4296 | ~v_4295 | v_4319;
assign x_426 = v_56 | v_61 | v_50 | v_59 | v_58 | v_144 | v_145 | v_143 | v_142 | v_166 | v_165 | v_146 | ~v_374 | ~v_373 | ~v_266 | ~v_265 | ~v_372 | ~v_371 | ~v_494 | ~v_493 | ~v_492 | ~v_491 | ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_244 | ~v_243 | ~v_364 | ~v_363 | ~v_1317 | ~v_1316 | ~v_1315 | ~v_1314 | ~v_1313 | ~v_1312 | ~v_1395 | ~v_1394 | ~v_1393 | ~v_1392 | ~v_4293 | ~v_4292 | ~v_4291 | ~v_4290 | v_4318;
assign x_427 = v_13 | v_7 | v_18 | v_16 | v_15 | v_136 | v_135 | v_134 | v_137 | v_138 | v_162 | v_161 | ~v_359 | ~v_358 | ~v_233 | ~v_232 | ~v_357 | ~v_356 | ~v_489 | ~v_488 | ~v_487 | ~v_486 | ~v_215 | ~v_214 | ~v_213 | ~v_212 | ~v_211 | ~v_210 | ~v_349 | ~v_348 | ~v_1292 | ~v_1291 | ~v_1290 | ~v_1289 | ~v_1288 | ~v_1287 | ~v_1386 | ~v_1385 | ~v_1384 | ~v_1383 | ~v_4288 | ~v_4287 | ~v_4286 | ~v_4285 | v_4317;
assign x_428 = v_4316 | ~v_4313;
assign x_429 = v_4316 | ~v_4314;
assign x_430 = v_4316 | ~v_4315;
assign x_431 = v_103 | v_101 | v_100 | v_99 | v_92 | v_102 | v_171 | v_170 | v_169 | v_149 | v_148 | v_147 | ~v_703 | ~v_702 | ~v_483 | ~v_482 | ~v_701 | ~v_653 | ~v_700 | ~v_652 | ~v_473 | ~v_472 | ~v_279 | ~v_471 | ~v_470 | ~v_276 | ~v_645 | ~v_644 | ~v_643 | ~v_642 | ~v_1460 | ~v_1459 | ~v_1340 | ~v_1458 | ~v_1457 | ~v_1337 | ~v_1376 | ~v_1375 | ~v_1374 | ~v_1373 | ~v_4298 | ~v_4297 | ~v_4296 | ~v_4295 | v_4315;
assign x_432 = v_61 | v_50 | v_60 | v_59 | v_58 | v_57 | v_144 | v_143 | v_142 | v_167 | v_166 | v_165 | ~v_698 | ~v_697 | ~v_468 | ~v_467 | ~v_696 | ~v_638 | ~v_695 | ~v_637 | ~v_458 | ~v_457 | ~v_246 | ~v_456 | ~v_455 | ~v_243 | ~v_630 | ~v_629 | ~v_628 | ~v_627 | ~v_1451 | ~v_1450 | ~v_1315 | ~v_1449 | ~v_1448 | ~v_1312 | ~v_1367 | ~v_1366 | ~v_1365 | ~v_1364 | ~v_4293 | ~v_4292 | ~v_4291 | ~v_4290 | v_4314;
assign x_433 = v_7 | v_18 | v_17 | v_16 | v_15 | v_14 | ~v_453 | ~v_452 | v_136 | v_135 | v_134 | v_163 | v_162 | v_161 | ~v_693 | ~v_692 | ~v_691 | ~v_623 | ~v_690 | ~v_622 | ~v_443 | ~v_442 | ~v_213 | ~v_441 | ~v_440 | ~v_210 | ~v_615 | ~v_614 | ~v_613 | ~v_612 | ~v_1442 | ~v_1441 | ~v_1290 | ~v_1440 | ~v_1439 | ~v_1287 | ~v_1358 | ~v_1357 | ~v_1356 | ~v_1355 | ~v_4288 | ~v_4287 | ~v_4286 | ~v_4285 | v_4313;
assign x_434 = v_4312 | ~v_4309;
assign x_435 = v_4312 | ~v_4310;
assign x_436 = v_4312 | ~v_4311;
assign x_437 = v_103 | v_97 | v_96 | v_100 | v_92 | v_151 | v_171 | v_170 | v_169 | v_160 | v_150 | v_147 | ~v_655 | ~v_654 | ~v_297 | ~v_296 | ~v_653 | ~v_652 | ~v_651 | ~v_650 | ~v_279 | ~v_276 | ~v_275 | ~v_274 | ~v_273 | ~v_272 | ~v_645 | ~v_644 | ~v_643 | ~v_642 | ~v_1340 | ~v_1337 | ~v_1432 | ~v_1431 | ~v_1430 | ~v_1429 | ~v_1376 | ~v_1375 | ~v_1374 | ~v_1373 | ~v_4298 | ~v_4297 | ~v_4296 | ~v_4295 | v_4311;
assign x_438 = v_54 | v_55 | v_61 | v_50 | v_58 | v_159 | v_145 | v_142 | v_167 | v_166 | v_165 | v_146 | ~v_640 | ~v_639 | ~v_264 | ~v_263 | ~v_638 | ~v_637 | ~v_636 | ~v_635 | ~v_246 | ~v_243 | ~v_242 | ~v_241 | ~v_240 | ~v_239 | ~v_630 | ~v_629 | ~v_628 | ~v_627 | ~v_1315 | ~v_1312 | ~v_1423 | ~v_1422 | ~v_1421 | ~v_1420 | ~v_1367 | ~v_1366 | ~v_1365 | ~v_1364 | ~v_4293 | ~v_4292 | ~v_4291 | ~v_4290 | v_4310;
assign x_439 = v_7 | v_18 | v_15 | v_12 | v_11 | v_134 | v_137 | v_138 | v_163 | v_162 | v_161 | v_155 | ~v_625 | ~v_624 | ~v_231 | ~v_230 | ~v_623 | ~v_622 | ~v_621 | ~v_620 | ~v_213 | ~v_210 | ~v_209 | ~v_208 | ~v_207 | ~v_206 | ~v_615 | ~v_614 | ~v_613 | ~v_612 | ~v_1290 | ~v_1287 | ~v_1414 | ~v_1413 | ~v_1412 | ~v_1411 | ~v_1358 | ~v_1357 | ~v_1356 | ~v_1355 | ~v_4288 | ~v_4287 | ~v_4286 | ~v_4285 | v_4309;
assign x_440 = v_4308 | ~v_4305;
assign x_441 = v_4308 | ~v_4306;
assign x_442 = v_4308 | ~v_4307;
assign x_443 = v_101 | v_100 | v_92 | v_102 | v_172 | v_171 | v_170 | v_169 | v_150 | v_149 | v_148 | v_147 | ~v_389 | ~v_388 | ~v_671 | ~v_670 | ~v_387 | ~v_386 | ~v_653 | ~v_652 | ~v_669 | ~v_668 | ~v_279 | ~v_276 | ~v_379 | ~v_378 | ~v_645 | ~v_644 | ~v_643 | ~v_642 | ~v_1340 | ~v_1337 | ~v_1404 | ~v_1403 | ~v_1402 | ~v_1401 | ~v_1376 | ~v_1375 | ~v_1374 | ~v_1373 | ~v_4298 | ~v_4297 | ~v_4296 | ~v_4295 | v_4307;
assign x_444 = v_50 | v_60 | v_59 | v_58 | v_144 | v_145 | v_143 | v_142 | v_168 | v_167 | v_166 | v_165 | ~v_374 | ~v_373 | ~v_666 | ~v_665 | ~v_372 | ~v_371 | ~v_638 | ~v_637 | ~v_664 | ~v_663 | ~v_246 | ~v_243 | ~v_364 | ~v_363 | ~v_630 | ~v_629 | ~v_628 | ~v_627 | ~v_1315 | ~v_1312 | ~v_1395 | ~v_1394 | ~v_1393 | ~v_1392 | ~v_1367 | ~v_1366 | ~v_1365 | ~v_1364 | ~v_4293 | ~v_4292 | ~v_4291 | ~v_4290 | v_4306;
assign x_445 = v_7 | v_17 | v_16 | v_15 | v_136 | v_135 | v_134 | v_137 | v_164 | v_163 | v_162 | v_161 | ~v_359 | ~v_358 | ~v_661 | ~v_660 | ~v_357 | ~v_356 | ~v_623 | ~v_622 | ~v_659 | ~v_658 | ~v_213 | ~v_210 | ~v_349 | ~v_348 | ~v_615 | ~v_614 | ~v_613 | ~v_612 | ~v_1290 | ~v_1287 | ~v_1386 | ~v_1385 | ~v_1384 | ~v_1383 | ~v_1358 | ~v_1357 | ~v_1356 | ~v_1355 | ~v_4288 | ~v_4287 | ~v_4286 | ~v_4285 | v_4305;
assign x_446 = v_4304 | ~v_4301;
assign x_447 = v_4304 | ~v_4302;
assign x_448 = v_4304 | ~v_4303;
assign x_449 = v_103 | v_101 | v_100 | v_95 | v_92 | v_102 | v_171 | v_170 | v_169 | v_150 | v_149 | v_148 | ~v_435 | ~v_434 | ~v_653 | ~v_652 | ~v_687 | ~v_686 | ~v_685 | ~v_684 | ~v_279 | ~v_276 | ~v_427 | ~v_426 | ~v_425 | ~v_424 | ~v_645 | ~v_644 | ~v_643 | ~v_642 | ~v_1340 | ~v_1337 | ~v_1336 | ~v_1335 | ~v_1334 | ~v_1333 | ~v_1376 | ~v_1375 | ~v_1374 | ~v_1373 | ~v_4298 | ~v_4297 | ~v_4296 | ~v_4295 | v_4303;
assign x_450 = v_53 | v_61 | v_50 | v_60 | v_59 | v_58 | v_144 | v_145 | v_143 | v_167 | v_166 | v_165 | ~v_420 | ~v_419 | ~v_638 | ~v_637 | ~v_682 | ~v_681 | ~v_680 | ~v_679 | ~v_246 | ~v_243 | ~v_412 | ~v_411 | ~v_410 | ~v_409 | ~v_630 | ~v_629 | ~v_628 | ~v_627 | ~v_1315 | ~v_1312 | ~v_1311 | ~v_1310 | ~v_1309 | ~v_1308 | ~v_1367 | ~v_1366 | ~v_1365 | ~v_1364 | ~v_4293 | ~v_4292 | ~v_4291 | ~v_4290 | v_4302;
assign x_451 = v_7 | v_18 | v_17 | v_16 | v_15 | v_10 | v_136 | v_135 | v_137 | v_163 | v_162 | v_161 | ~v_405 | ~v_404 | ~v_623 | ~v_622 | ~v_677 | ~v_676 | ~v_675 | ~v_674 | ~v_213 | ~v_210 | ~v_397 | ~v_396 | ~v_395 | ~v_394 | ~v_615 | ~v_614 | ~v_613 | ~v_612 | ~v_1290 | ~v_1287 | ~v_1286 | ~v_1285 | ~v_1284 | ~v_1283 | ~v_1358 | ~v_1357 | ~v_1356 | ~v_1355 | ~v_4288 | ~v_4287 | ~v_4286 | ~v_4285 | v_4301;
assign x_452 = v_4300 | ~v_4289;
assign x_453 = v_4300 | ~v_4294;
assign x_454 = v_4300 | ~v_4299;
assign x_455 = v_98 | v_103 | v_101 | v_100 | v_92 | v_102 | v_170 | v_169 | v_150 | v_149 | v_148 | v_147 | ~v_609 | ~v_608 | ~v_299 | ~v_298 | ~v_435 | ~v_434 | ~v_607 | ~v_606 | ~v_281 | ~v_280 | ~v_279 | ~v_278 | ~v_277 | ~v_276 | ~v_427 | ~v_426 | ~v_425 | ~v_424 | ~v_1342 | ~v_1341 | ~v_1340 | ~v_1339 | ~v_1338 | ~v_1337 | ~v_1336 | ~v_1335 | ~v_1334 | ~v_1333 | ~v_4298 | ~v_4297 | ~v_4296 | ~v_4295 | v_4299;
assign x_456 = v_4298 | v_158;
assign x_457 = v_4298 | v_123;
assign x_458 = v_4297 | v_158;
assign x_459 = v_4297 | v_120;
assign x_460 = v_4296 | ~v_158;
assign x_461 = v_4296 | v_108;
assign x_462 = v_4295 | ~v_158;
assign x_463 = v_4295 | v_105;
assign x_464 = v_56 | v_61 | v_50 | v_60 | v_59 | v_58 | v_144 | v_145 | v_143 | v_142 | v_166 | v_165 | ~v_604 | ~v_603 | ~v_266 | ~v_265 | ~v_420 | ~v_419 | ~v_602 | ~v_601 | ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_244 | ~v_243 | ~v_412 | ~v_411 | ~v_410 | ~v_409 | ~v_1317 | ~v_1316 | ~v_1315 | ~v_1314 | ~v_1313 | ~v_1312 | ~v_1311 | ~v_1310 | ~v_1309 | ~v_1308 | ~v_4293 | ~v_4292 | ~v_4291 | ~v_4290 | v_4294;
assign x_465 = v_4293 | v_158;
assign x_466 = v_4293 | v_81;
assign x_467 = v_4292 | v_158;
assign x_468 = v_4292 | v_78;
assign x_469 = v_4291 | ~v_158;
assign x_470 = v_4291 | v_66;
assign x_471 = v_4290 | ~v_158;
assign x_472 = v_4290 | v_63;
assign x_473 = v_13 | v_7 | v_18 | v_17 | v_16 | v_15 | v_136 | v_135 | v_134 | v_137 | v_162 | v_161 | ~v_599 | ~v_598 | ~v_233 | ~v_232 | ~v_405 | ~v_404 | ~v_597 | ~v_596 | ~v_215 | ~v_214 | ~v_213 | ~v_212 | ~v_211 | ~v_210 | ~v_397 | ~v_396 | ~v_395 | ~v_394 | ~v_1292 | ~v_1291 | ~v_1290 | ~v_1289 | ~v_1288 | ~v_1287 | ~v_1286 | ~v_1285 | ~v_1284 | ~v_1283 | ~v_4288 | ~v_4287 | ~v_4286 | ~v_4285 | v_4289;
assign x_474 = v_4288 | v_158;
assign x_475 = v_4288 | v_39;
assign x_476 = v_4287 | v_158;
assign x_477 = v_4287 | v_36;
assign x_478 = v_4286 | ~v_158;
assign x_479 = v_4286 | v_24;
assign x_480 = v_4285 | ~v_158;
assign x_481 = v_4285 | v_21;
assign x_482 = v_4284 | ~v_4203;
assign x_483 = v_4284 | ~v_4283;
assign x_484 = v_140 | v_139 | ~v_4282 | ~v_2405 | ~v_2404 | ~v_4205 | ~v_4204 | v_4283;
assign x_485 = v_4282 | ~v_4221;
assign x_486 = v_4282 | ~v_4225;
assign x_487 = v_4282 | ~v_4229;
assign x_488 = v_4282 | ~v_4233;
assign x_489 = v_4282 | ~v_4237;
assign x_490 = v_4282 | ~v_4241;
assign x_491 = v_4282 | ~v_4245;
assign x_492 = v_4282 | ~v_4249;
assign x_493 = v_4282 | ~v_4253;
assign x_494 = v_4282 | ~v_4257;
assign x_495 = v_4282 | ~v_4261;
assign x_496 = v_4282 | ~v_4265;
assign x_497 = v_4282 | ~v_4269;
assign x_498 = v_4282 | ~v_4273;
assign x_499 = v_4282 | ~v_4277;
assign x_500 = v_4282 | ~v_4281;
assign x_501 = v_4282 | ~v_1263;
assign x_502 = v_4282 | ~v_1264;
assign x_503 = v_4282 | ~v_1265;
assign x_504 = v_4282 | ~v_1266;
assign x_505 = ~v_4280 | ~v_4279 | ~v_4278 | v_4281;
assign x_506 = v_4280 | ~v_3496;
assign x_507 = v_4280 | ~v_3497;
assign x_508 = v_4280 | ~v_3564;
assign x_509 = v_4280 | ~v_3498;
assign x_510 = v_4280 | ~v_3565;
assign x_511 = v_4280 | ~v_3499;
assign x_512 = v_4280 | ~v_3500;
assign x_513 = v_4280 | ~v_3566;
assign x_514 = v_4280 | ~v_3501;
assign x_515 = v_4280 | ~v_3567;
assign x_516 = v_4280 | ~v_2075;
assign x_517 = v_4280 | ~v_4216;
assign x_518 = v_4280 | ~v_2076;
assign x_519 = v_4280 | ~v_2141;
assign x_520 = v_4280 | ~v_4217;
assign x_521 = v_4280 | ~v_2077;
assign x_522 = v_4280 | ~v_2142;
assign x_523 = v_4280 | ~v_2078;
assign x_524 = v_4280 | ~v_4218;
assign x_525 = v_4280 | ~v_2079;
assign x_526 = v_4280 | ~v_2143;
assign x_527 = v_4280 | ~v_4219;
assign x_528 = v_4280 | ~v_2080;
assign x_529 = v_4280 | ~v_2144;
assign x_530 = v_4280 | ~v_839;
assign x_531 = v_4280 | ~v_1257;
assign x_532 = v_4280 | ~v_1023;
assign x_533 = v_4280 | ~v_840;
assign x_534 = v_4280 | ~v_1258;
assign x_535 = v_4280 | ~v_1024;
assign x_536 = v_4280 | ~v_184;
assign x_537 = v_4280 | ~v_169;
assign x_538 = v_4280 | ~v_148;
assign x_539 = v_4280 | ~v_1259;
assign x_540 = v_4280 | ~v_1260;
assign x_541 = v_4280 | ~v_103;
assign x_542 = v_4280 | ~v_102;
assign x_543 = v_4280 | ~v_101;
assign x_544 = v_4280 | ~v_100;
assign x_545 = v_4280 | ~v_99;
assign x_546 = v_4280 | ~v_98;
assign x_547 = v_4280 | ~v_97;
assign x_548 = v_4280 | ~v_95;
assign x_549 = v_4280 | ~v_94;
assign x_550 = v_4279 | ~v_3481;
assign x_551 = v_4279 | ~v_3482;
assign x_552 = v_4279 | ~v_3559;
assign x_553 = v_4279 | ~v_3483;
assign x_554 = v_4279 | ~v_3560;
assign x_555 = v_4279 | ~v_3484;
assign x_556 = v_4279 | ~v_3485;
assign x_557 = v_4279 | ~v_2060;
assign x_558 = v_4279 | ~v_4211;
assign x_559 = v_4279 | ~v_2061;
assign x_560 = v_4279 | ~v_2136;
assign x_561 = v_4279 | ~v_4212;
assign x_562 = v_4279 | ~v_2062;
assign x_563 = v_4279 | ~v_2137;
assign x_564 = v_4279 | ~v_2063;
assign x_565 = v_4279 | ~v_4213;
assign x_566 = v_4279 | ~v_2064;
assign x_567 = v_4279 | ~v_2138;
assign x_568 = v_4279 | ~v_4214;
assign x_569 = v_4279 | ~v_2065;
assign x_570 = v_4279 | ~v_2139;
assign x_571 = v_4279 | ~v_806;
assign x_572 = v_4279 | ~v_1252;
assign x_573 = v_4279 | ~v_1008;
assign x_574 = v_4279 | ~v_1253;
assign x_575 = v_4279 | ~v_1009;
assign x_576 = v_4279 | ~v_3561;
assign x_577 = v_4279 | ~v_807;
assign x_578 = v_4279 | ~v_3486;
assign x_579 = v_4279 | ~v_3562;
assign x_580 = v_4279 | ~v_183;
assign x_581 = v_4279 | ~v_165;
assign x_582 = v_4279 | ~v_143;
assign x_583 = v_4279 | ~v_1254;
assign x_584 = v_4279 | ~v_1255;
assign x_585 = v_4279 | ~v_61;
assign x_586 = v_4279 | ~v_60;
assign x_587 = v_4279 | ~v_59;
assign x_588 = v_4279 | ~v_58;
assign x_589 = v_4279 | ~v_57;
assign x_590 = v_4279 | ~v_56;
assign x_591 = v_4279 | ~v_55;
assign x_592 = v_4279 | ~v_53;
assign x_593 = v_4279 | ~v_52;
assign x_594 = v_4278 | ~v_3466;
assign x_595 = v_4278 | ~v_3467;
assign x_596 = v_4278 | ~v_3554;
assign x_597 = v_4278 | ~v_3468;
assign x_598 = v_4278 | ~v_3555;
assign x_599 = v_4278 | ~v_3469;
assign x_600 = v_4278 | ~v_3556;
assign x_601 = v_4278 | ~v_3470;
assign x_602 = v_4278 | ~v_3557;
assign x_603 = v_4278 | ~v_2045;
assign x_604 = v_4278 | ~v_4206;
assign x_605 = v_4278 | ~v_2046;
assign x_606 = v_4278 | ~v_2131;
assign x_607 = v_4278 | ~v_4207;
assign x_608 = v_4278 | ~v_2047;
assign x_609 = v_4278 | ~v_2132;
assign x_610 = v_4278 | ~v_2048;
assign x_611 = v_4278 | ~v_4208;
assign x_612 = v_4278 | ~v_2049;
assign x_613 = v_4278 | ~v_2133;
assign x_614 = v_4278 | ~v_4209;
assign x_615 = v_4278 | ~v_2050;
assign x_616 = v_4278 | ~v_2134;
assign x_617 = v_4278 | ~v_773;
assign x_618 = v_4278 | ~v_774;
assign x_619 = v_4278 | ~v_182;
assign x_620 = v_4278 | ~v_161;
assign x_621 = v_4278 | ~v_3473;
assign x_622 = v_4278 | ~v_1247;
assign x_623 = v_4278 | ~v_1248;
assign x_624 = v_4278 | ~v_135;
assign x_625 = v_4278 | ~v_1249;
assign x_626 = v_4278 | ~v_993;
assign x_627 = v_4278 | ~v_1250;
assign x_628 = v_4278 | ~v_994;
assign x_629 = v_4278 | ~v_18;
assign x_630 = v_4278 | ~v_17;
assign x_631 = v_4278 | ~v_16;
assign x_632 = v_4278 | ~v_15;
assign x_633 = v_4278 | ~v_14;
assign x_634 = v_4278 | ~v_13;
assign x_635 = v_4278 | ~v_12;
assign x_636 = v_4278 | ~v_10;
assign x_637 = v_4278 | ~v_9;
assign x_638 = ~v_4276 | ~v_4275 | ~v_4274 | v_4277;
assign x_639 = v_4276 | ~v_3584;
assign x_640 = v_4276 | ~v_3585;
assign x_641 = v_4276 | ~v_3586;
assign x_642 = v_4276 | ~v_3587;
assign x_643 = v_4276 | ~v_2193;
assign x_644 = v_4276 | ~v_2194;
assign x_645 = v_4276 | ~v_2195;
assign x_646 = v_4276 | ~v_2196;
assign x_647 = v_4276 | ~v_3496;
assign x_648 = v_4276 | ~v_3564;
assign x_649 = v_4276 | ~v_3565;
assign x_650 = v_4276 | ~v_3499;
assign x_651 = v_4276 | ~v_3566;
assign x_652 = v_4276 | ~v_3567;
assign x_653 = v_4276 | ~v_2075;
assign x_654 = v_4276 | ~v_4216;
assign x_655 = v_4276 | ~v_2141;
assign x_656 = v_4276 | ~v_4217;
assign x_657 = v_4276 | ~v_2142;
assign x_658 = v_4276 | ~v_2078;
assign x_659 = v_4276 | ~v_4218;
assign x_660 = v_4276 | ~v_2143;
assign x_661 = v_4276 | ~v_4219;
assign x_662 = v_4276 | ~v_2144;
assign x_663 = v_4276 | ~v_1085;
assign x_664 = v_4276 | ~v_1131;
assign x_665 = v_4276 | ~v_1132;
assign x_666 = v_4276 | ~v_1086;
assign x_667 = v_4276 | ~v_1133;
assign x_668 = v_4276 | ~v_1134;
assign x_669 = v_4276 | ~v_1023;
assign x_670 = v_4276 | ~v_1024;
assign x_671 = v_4276 | ~v_184;
assign x_672 = v_4276 | ~v_172;
assign x_673 = v_4276 | ~v_171;
assign x_674 = v_4276 | ~v_170;
assign x_675 = v_4276 | ~v_148;
assign x_676 = v_4276 | ~v_147;
assign x_677 = v_4276 | ~v_102;
assign x_678 = v_4276 | ~v_101;
assign x_679 = v_4276 | ~v_100;
assign x_680 = v_4276 | ~v_99;
assign x_681 = v_4276 | ~v_97;
assign x_682 = v_4276 | ~v_93;
assign x_683 = v_4275 | ~v_3579;
assign x_684 = v_4275 | ~v_3580;
assign x_685 = v_4275 | ~v_3581;
assign x_686 = v_4275 | ~v_3582;
assign x_687 = v_4275 | ~v_2188;
assign x_688 = v_4275 | ~v_2189;
assign x_689 = v_4275 | ~v_2190;
assign x_690 = v_4275 | ~v_2191;
assign x_691 = v_4275 | ~v_3481;
assign x_692 = v_4275 | ~v_3559;
assign x_693 = v_4275 | ~v_3560;
assign x_694 = v_4275 | ~v_3484;
assign x_695 = v_4275 | ~v_2060;
assign x_696 = v_4275 | ~v_4211;
assign x_697 = v_4275 | ~v_2136;
assign x_698 = v_4275 | ~v_4212;
assign x_699 = v_4275 | ~v_2137;
assign x_700 = v_4275 | ~v_2063;
assign x_701 = v_4275 | ~v_4213;
assign x_702 = v_4275 | ~v_2138;
assign x_703 = v_4275 | ~v_4214;
assign x_704 = v_4275 | ~v_2139;
assign x_705 = v_4275 | ~v_1070;
assign x_706 = v_4275 | ~v_1126;
assign x_707 = v_4275 | ~v_1127;
assign x_708 = v_4275 | ~v_1071;
assign x_709 = v_4275 | ~v_1128;
assign x_710 = v_4275 | ~v_1129;
assign x_711 = v_4275 | ~v_1008;
assign x_712 = v_4275 | ~v_1009;
assign x_713 = v_4275 | ~v_3561;
assign x_714 = v_4275 | ~v_3562;
assign x_715 = v_4275 | ~v_183;
assign x_716 = v_4275 | ~v_168;
assign x_717 = v_4275 | ~v_167;
assign x_718 = v_4275 | ~v_166;
assign x_719 = v_4275 | ~v_143;
assign x_720 = v_4275 | ~v_142;
assign x_721 = v_4275 | ~v_60;
assign x_722 = v_4275 | ~v_59;
assign x_723 = v_4275 | ~v_58;
assign x_724 = v_4275 | ~v_57;
assign x_725 = v_4275 | ~v_55;
assign x_726 = v_4275 | ~v_51;
assign x_727 = v_4274 | ~v_3574;
assign x_728 = v_4274 | ~v_3575;
assign x_729 = v_4274 | ~v_3576;
assign x_730 = v_4274 | ~v_3577;
assign x_731 = v_4274 | ~v_2183;
assign x_732 = v_4274 | ~v_2184;
assign x_733 = v_4274 | ~v_2185;
assign x_734 = v_4274 | ~v_2186;
assign x_735 = v_4274 | ~v_3466;
assign x_736 = v_4274 | ~v_3554;
assign x_737 = v_4274 | ~v_3555;
assign x_738 = v_4274 | ~v_3469;
assign x_739 = v_4274 | ~v_3556;
assign x_740 = v_4274 | ~v_3557;
assign x_741 = v_4274 | ~v_2045;
assign x_742 = v_4274 | ~v_4206;
assign x_743 = v_4274 | ~v_2131;
assign x_744 = v_4274 | ~v_4207;
assign x_745 = v_4274 | ~v_2132;
assign x_746 = v_4274 | ~v_2048;
assign x_747 = v_4274 | ~v_4208;
assign x_748 = v_4274 | ~v_2133;
assign x_749 = v_4274 | ~v_4209;
assign x_750 = v_4274 | ~v_2134;
assign x_751 = v_4274 | ~v_1055;
assign x_752 = v_4274 | ~v_1121;
assign x_753 = v_4274 | ~v_1122;
assign x_754 = v_4274 | ~v_1056;
assign x_755 = v_4274 | ~v_1123;
assign x_756 = v_4274 | ~v_1124;
assign x_757 = v_4274 | ~v_182;
assign x_758 = v_4274 | ~v_164;
assign x_759 = v_4274 | ~v_163;
assign x_760 = v_4274 | ~v_162;
assign x_761 = v_4274 | ~v_135;
assign x_762 = v_4274 | ~v_134;
assign x_763 = v_4274 | ~v_993;
assign x_764 = v_4274 | ~v_994;
assign x_765 = v_4274 | ~v_17;
assign x_766 = v_4274 | ~v_16;
assign x_767 = v_4274 | ~v_15;
assign x_768 = v_4274 | ~v_14;
assign x_769 = v_4274 | ~v_12;
assign x_770 = v_4274 | ~v_8;
assign x_771 = ~v_4272 | ~v_4271 | ~v_4270 | v_4273;
assign x_772 = v_4272 | ~v_3532;
assign x_773 = v_4272 | ~v_3533;
assign x_774 = v_4272 | ~v_3534;
assign x_775 = v_4272 | ~v_3535;
assign x_776 = v_4272 | ~v_2125;
assign x_777 = v_4272 | ~v_2126;
assign x_778 = v_4272 | ~v_2127;
assign x_779 = v_4272 | ~v_2128;
assign x_780 = v_4272 | ~v_3584;
assign x_781 = v_4272 | ~v_3585;
assign x_782 = v_4272 | ~v_3586;
assign x_783 = v_4272 | ~v_3587;
assign x_784 = v_4272 | ~v_2193;
assign x_785 = v_4272 | ~v_2194;
assign x_786 = v_4272 | ~v_2195;
assign x_787 = v_4272 | ~v_2196;
assign x_788 = v_4272 | ~v_3496;
assign x_789 = v_4272 | ~v_3499;
assign x_790 = v_4272 | ~v_2075;
assign x_791 = v_4272 | ~v_4216;
assign x_792 = v_4272 | ~v_4217;
assign x_793 = v_4272 | ~v_2078;
assign x_794 = v_4272 | ~v_4218;
assign x_795 = v_4272 | ~v_4219;
assign x_796 = v_4272 | ~v_927;
assign x_797 = v_4272 | ~v_928;
assign x_798 = v_4272 | ~v_1099;
assign x_799 = v_4272 | ~v_1100;
assign x_800 = v_4272 | ~v_1101;
assign x_801 = v_4272 | ~v_1102;
assign x_802 = v_4272 | ~v_1085;
assign x_803 = v_4272 | ~v_1086;
assign x_804 = v_4272 | ~v_184;
assign x_805 = v_4272 | ~v_171;
assign x_806 = v_4272 | ~v_170;
assign x_807 = v_4272 | ~v_150;
assign x_808 = v_4272 | ~v_149;
assign x_809 = v_4272 | ~v_103;
assign x_810 = v_4272 | ~v_102;
assign x_811 = v_4272 | ~v_101;
assign x_812 = v_4272 | ~v_100;
assign x_813 = v_4272 | ~v_96;
assign x_814 = v_4272 | ~v_95;
assign x_815 = v_4272 | ~v_93;
assign x_816 = v_4271 | ~v_3527;
assign x_817 = v_4271 | ~v_3528;
assign x_818 = v_4271 | ~v_3529;
assign x_819 = v_4271 | ~v_3530;
assign x_820 = v_4271 | ~v_2120;
assign x_821 = v_4271 | ~v_2121;
assign x_822 = v_4271 | ~v_2122;
assign x_823 = v_4271 | ~v_2123;
assign x_824 = v_4271 | ~v_3579;
assign x_825 = v_4271 | ~v_3580;
assign x_826 = v_4271 | ~v_3581;
assign x_827 = v_4271 | ~v_3582;
assign x_828 = v_4271 | ~v_2188;
assign x_829 = v_4271 | ~v_2189;
assign x_830 = v_4271 | ~v_2190;
assign x_831 = v_4271 | ~v_2191;
assign x_832 = v_4271 | ~v_3481;
assign x_833 = v_4271 | ~v_3484;
assign x_834 = v_4271 | ~v_2060;
assign x_835 = v_4271 | ~v_4211;
assign x_836 = v_4271 | ~v_4212;
assign x_837 = v_4271 | ~v_2063;
assign x_838 = v_4271 | ~v_4213;
assign x_839 = v_4271 | ~v_4214;
assign x_840 = v_4271 | ~v_912;
assign x_841 = v_4271 | ~v_913;
assign x_842 = v_4271 | ~v_1094;
assign x_843 = v_4271 | ~v_1095;
assign x_844 = v_4271 | ~v_1096;
assign x_845 = v_4271 | ~v_1097;
assign x_846 = v_4271 | ~v_1070;
assign x_847 = v_4271 | ~v_1071;
assign x_848 = v_4271 | ~v_183;
assign x_849 = v_4271 | ~v_167;
assign x_850 = v_4271 | ~v_166;
assign x_851 = v_4271 | ~v_145;
assign x_852 = v_4271 | ~v_144;
assign x_853 = v_4271 | ~v_61;
assign x_854 = v_4271 | ~v_60;
assign x_855 = v_4271 | ~v_59;
assign x_856 = v_4271 | ~v_58;
assign x_857 = v_4271 | ~v_54;
assign x_858 = v_4271 | ~v_53;
assign x_859 = v_4271 | ~v_51;
assign x_860 = v_4270 | ~v_3522;
assign x_861 = v_4270 | ~v_3523;
assign x_862 = v_4270 | ~v_3524;
assign x_863 = v_4270 | ~v_3525;
assign x_864 = v_4270 | ~v_2115;
assign x_865 = v_4270 | ~v_2116;
assign x_866 = v_4270 | ~v_2117;
assign x_867 = v_4270 | ~v_2118;
assign x_868 = v_4270 | ~v_3574;
assign x_869 = v_4270 | ~v_3575;
assign x_870 = v_4270 | ~v_3576;
assign x_871 = v_4270 | ~v_3577;
assign x_872 = v_4270 | ~v_2183;
assign x_873 = v_4270 | ~v_2184;
assign x_874 = v_4270 | ~v_2185;
assign x_875 = v_4270 | ~v_2186;
assign x_876 = v_4270 | ~v_3466;
assign x_877 = v_4270 | ~v_3469;
assign x_878 = v_4270 | ~v_2045;
assign x_879 = v_4270 | ~v_4206;
assign x_880 = v_4270 | ~v_4207;
assign x_881 = v_4270 | ~v_2048;
assign x_882 = v_4270 | ~v_4208;
assign x_883 = v_4270 | ~v_4209;
assign x_884 = v_4270 | ~v_897;
assign x_885 = v_4270 | ~v_898;
assign x_886 = v_4270 | ~v_1089;
assign x_887 = v_4270 | ~v_1090;
assign x_888 = v_4270 | ~v_1091;
assign x_889 = v_4270 | ~v_1092;
assign x_890 = v_4270 | ~v_1055;
assign x_891 = v_4270 | ~v_1056;
assign x_892 = v_4270 | ~v_182;
assign x_893 = v_4270 | ~v_163;
assign x_894 = v_4270 | ~v_162;
assign x_895 = v_4270 | ~v_137;
assign x_896 = v_4270 | ~v_136;
assign x_897 = v_4270 | ~v_18;
assign x_898 = v_4270 | ~v_17;
assign x_899 = v_4270 | ~v_16;
assign x_900 = v_4270 | ~v_15;
assign x_901 = v_4270 | ~v_11;
assign x_902 = v_4270 | ~v_10;
assign x_903 = v_4270 | ~v_8;
assign x_904 = ~v_4268 | ~v_4267 | ~v_4266 | v_4269;
assign x_905 = v_4268 | ~v_3494;
assign x_906 = v_4268 | ~v_3495;
assign x_907 = v_4268 | ~v_2109;
assign x_908 = v_4268 | ~v_2110;
assign x_909 = v_4268 | ~v_2111;
assign x_910 = v_4268 | ~v_2112;
assign x_911 = v_4268 | ~v_3584;
assign x_912 = v_4268 | ~v_3585;
assign x_913 = v_4268 | ~v_3586;
assign x_914 = v_4268 | ~v_3587;
assign x_915 = v_4268 | ~v_2193;
assign x_916 = v_4268 | ~v_2194;
assign x_917 = v_4268 | ~v_2195;
assign x_918 = v_4268 | ~v_2196;
assign x_919 = v_4268 | ~v_3496;
assign x_920 = v_4268 | ~v_3499;
assign x_921 = v_4268 | ~v_2075;
assign x_922 = v_4268 | ~v_4216;
assign x_923 = v_4268 | ~v_4217;
assign x_924 = v_4268 | ~v_2078;
assign x_925 = v_4268 | ~v_4218;
assign x_926 = v_4268 | ~v_4219;
assign x_927 = v_4268 | ~v_975;
assign x_928 = v_4268 | ~v_976;
assign x_929 = v_4268 | ~v_1115;
assign x_930 = v_4268 | ~v_1116;
assign x_931 = v_4268 | ~v_1085;
assign x_932 = v_4268 | ~v_1086;
assign x_933 = v_4268 | ~v_1117;
assign x_934 = v_4268 | ~v_1118;
assign x_935 = v_4268 | ~v_3502;
assign x_936 = v_4268 | ~v_3503;
assign x_937 = v_4268 | ~v_184;
assign x_938 = v_4268 | ~v_171;
assign x_939 = v_4268 | ~v_170;
assign x_940 = v_4268 | ~v_151;
assign x_941 = v_4268 | ~v_150;
assign x_942 = v_4268 | ~v_149;
assign x_943 = v_4268 | ~v_148;
assign x_944 = v_4268 | ~v_147;
assign x_945 = v_4268 | ~v_103;
assign x_946 = v_4268 | ~v_101;
assign x_947 = v_4268 | ~v_100;
assign x_948 = v_4268 | ~v_93;
assign x_949 = v_4267 | ~v_3479;
assign x_950 = v_4267 | ~v_3480;
assign x_951 = v_4267 | ~v_2104;
assign x_952 = v_4267 | ~v_2105;
assign x_953 = v_4267 | ~v_2106;
assign x_954 = v_4267 | ~v_2107;
assign x_955 = v_4267 | ~v_3579;
assign x_956 = v_4267 | ~v_3580;
assign x_957 = v_4267 | ~v_3581;
assign x_958 = v_4267 | ~v_3582;
assign x_959 = v_4267 | ~v_2188;
assign x_960 = v_4267 | ~v_2189;
assign x_961 = v_4267 | ~v_2190;
assign x_962 = v_4267 | ~v_2191;
assign x_963 = v_4267 | ~v_3481;
assign x_964 = v_4267 | ~v_3484;
assign x_965 = v_4267 | ~v_2060;
assign x_966 = v_4267 | ~v_4211;
assign x_967 = v_4267 | ~v_4212;
assign x_968 = v_4267 | ~v_2063;
assign x_969 = v_4267 | ~v_4213;
assign x_970 = v_4267 | ~v_4214;
assign x_971 = v_4267 | ~v_960;
assign x_972 = v_4267 | ~v_961;
assign x_973 = v_4267 | ~v_1110;
assign x_974 = v_4267 | ~v_1111;
assign x_975 = v_4267 | ~v_1070;
assign x_976 = v_4267 | ~v_1071;
assign x_977 = v_4267 | ~v_1112;
assign x_978 = v_4267 | ~v_1113;
assign x_979 = v_4267 | ~v_3487;
assign x_980 = v_4267 | ~v_3488;
assign x_981 = v_4267 | ~v_183;
assign x_982 = v_4267 | ~v_167;
assign x_983 = v_4267 | ~v_166;
assign x_984 = v_4267 | ~v_146;
assign x_985 = v_4267 | ~v_145;
assign x_986 = v_4267 | ~v_144;
assign x_987 = v_4267 | ~v_143;
assign x_988 = v_4267 | ~v_142;
assign x_989 = v_4267 | ~v_61;
assign x_990 = v_4267 | ~v_59;
assign x_991 = v_4267 | ~v_58;
assign x_992 = v_4267 | ~v_51;
assign x_993 = v_4266 | ~v_3464;
assign x_994 = v_4266 | ~v_3465;
assign x_995 = v_4266 | ~v_2099;
assign x_996 = v_4266 | ~v_2100;
assign x_997 = v_4266 | ~v_2101;
assign x_998 = v_4266 | ~v_2102;
assign x_999 = v_4266 | ~v_3574;
assign x_1000 = v_4266 | ~v_3575;
assign x_1001 = v_4266 | ~v_3576;
assign x_1002 = v_4266 | ~v_3577;
assign x_1003 = v_4266 | ~v_2183;
assign x_1004 = v_4266 | ~v_2184;
assign x_1005 = v_4266 | ~v_2185;
assign x_1006 = v_4266 | ~v_2186;
assign x_1007 = v_4266 | ~v_3466;
assign x_1008 = v_4266 | ~v_3469;
assign x_1009 = v_4266 | ~v_2045;
assign x_1010 = v_4266 | ~v_4206;
assign x_1011 = v_4266 | ~v_4207;
assign x_1012 = v_4266 | ~v_2048;
assign x_1013 = v_4266 | ~v_4208;
assign x_1014 = v_4266 | ~v_4209;
assign x_1015 = v_4266 | ~v_945;
assign x_1016 = v_4266 | ~v_946;
assign x_1017 = v_4266 | ~v_1105;
assign x_1018 = v_4266 | ~v_1106;
assign x_1019 = v_4266 | ~v_1055;
assign x_1020 = v_4266 | ~v_1056;
assign x_1021 = v_4266 | ~v_1107;
assign x_1022 = v_4266 | ~v_1108;
assign x_1023 = v_4266 | ~v_3471;
assign x_1024 = v_4266 | ~v_3472;
assign x_1025 = v_4266 | ~v_182;
assign x_1026 = v_4266 | ~v_163;
assign x_1027 = v_4266 | ~v_162;
assign x_1028 = v_4266 | ~v_138;
assign x_1029 = v_4266 | ~v_137;
assign x_1030 = v_4266 | ~v_136;
assign x_1031 = v_4266 | ~v_135;
assign x_1032 = v_4266 | ~v_134;
assign x_1033 = v_4266 | ~v_18;
assign x_1034 = v_4266 | ~v_16;
assign x_1035 = v_4266 | ~v_15;
assign x_1036 = v_4266 | ~v_8;
assign x_1037 = ~v_4264 | ~v_4263 | ~v_4262 | v_4265;
assign x_1038 = v_4264 | ~v_3548;
assign x_1039 = v_4264 | ~v_3549;
assign x_1040 = v_4264 | ~v_3550;
assign x_1041 = v_4264 | ~v_3551;
assign x_1042 = v_4264 | ~v_2071;
assign x_1043 = v_4264 | ~v_2072;
assign x_1044 = v_4264 | ~v_2073;
assign x_1045 = v_4264 | ~v_2074;
assign x_1046 = v_4264 | ~v_3584;
assign x_1047 = v_4264 | ~v_3585;
assign x_1048 = v_4264 | ~v_3586;
assign x_1049 = v_4264 | ~v_3587;
assign x_1050 = v_4264 | ~v_2193;
assign x_1051 = v_4264 | ~v_2194;
assign x_1052 = v_4264 | ~v_2195;
assign x_1053 = v_4264 | ~v_2196;
assign x_1054 = v_4264 | ~v_3496;
assign x_1055 = v_4264 | ~v_3499;
assign x_1056 = v_4264 | ~v_2075;
assign x_1057 = v_4264 | ~v_4216;
assign x_1058 = v_4264 | ~v_4217;
assign x_1059 = v_4264 | ~v_2078;
assign x_1060 = v_4264 | ~v_4218;
assign x_1061 = v_4264 | ~v_4219;
assign x_1062 = v_4264 | ~v_837;
assign x_1063 = v_4264 | ~v_838;
assign x_1064 = v_4264 | ~v_1081;
assign x_1065 = v_4264 | ~v_1082;
assign x_1066 = v_4264 | ~v_1083;
assign x_1067 = v_4264 | ~v_1084;
assign x_1068 = v_4264 | ~v_1085;
assign x_1069 = v_4264 | ~v_1086;
assign x_1070 = v_4264 | ~v_184;
assign x_1071 = v_4264 | ~v_171;
assign x_1072 = v_4264 | ~v_170;
assign x_1073 = v_4264 | ~v_160;
assign x_1074 = v_4264 | ~v_150;
assign x_1075 = v_4264 | ~v_149;
assign x_1076 = v_4264 | ~v_148;
assign x_1077 = v_4264 | ~v_147;
assign x_1078 = v_4264 | ~v_103;
assign x_1079 = v_4264 | ~v_102;
assign x_1080 = v_4264 | ~v_100;
assign x_1081 = v_4264 | ~v_93;
assign x_1082 = v_4263 | ~v_3543;
assign x_1083 = v_4263 | ~v_3544;
assign x_1084 = v_4263 | ~v_3545;
assign x_1085 = v_4263 | ~v_3546;
assign x_1086 = v_4263 | ~v_2056;
assign x_1087 = v_4263 | ~v_2057;
assign x_1088 = v_4263 | ~v_2058;
assign x_1089 = v_4263 | ~v_2059;
assign x_1090 = v_4263 | ~v_3579;
assign x_1091 = v_4263 | ~v_3580;
assign x_1092 = v_4263 | ~v_3581;
assign x_1093 = v_4263 | ~v_3582;
assign x_1094 = v_4263 | ~v_2188;
assign x_1095 = v_4263 | ~v_2189;
assign x_1096 = v_4263 | ~v_2190;
assign x_1097 = v_4263 | ~v_2191;
assign x_1098 = v_4263 | ~v_3481;
assign x_1099 = v_4263 | ~v_3484;
assign x_1100 = v_4263 | ~v_2060;
assign x_1101 = v_4263 | ~v_4211;
assign x_1102 = v_4263 | ~v_4212;
assign x_1103 = v_4263 | ~v_2063;
assign x_1104 = v_4263 | ~v_4213;
assign x_1105 = v_4263 | ~v_4214;
assign x_1106 = v_4263 | ~v_804;
assign x_1107 = v_4263 | ~v_805;
assign x_1108 = v_4263 | ~v_1066;
assign x_1109 = v_4263 | ~v_1067;
assign x_1110 = v_4263 | ~v_1068;
assign x_1111 = v_4263 | ~v_1069;
assign x_1112 = v_4263 | ~v_1070;
assign x_1113 = v_4263 | ~v_1071;
assign x_1114 = v_4263 | ~v_183;
assign x_1115 = v_4263 | ~v_167;
assign x_1116 = v_4263 | ~v_166;
assign x_1117 = v_4263 | ~v_159;
assign x_1118 = v_4263 | ~v_145;
assign x_1119 = v_4263 | ~v_144;
assign x_1120 = v_4263 | ~v_143;
assign x_1121 = v_4263 | ~v_142;
assign x_1122 = v_4263 | ~v_61;
assign x_1123 = v_4263 | ~v_60;
assign x_1124 = v_4263 | ~v_58;
assign x_1125 = v_4263 | ~v_51;
assign x_1126 = v_4262 | ~v_3538;
assign x_1127 = v_4262 | ~v_3539;
assign x_1128 = v_4262 | ~v_3540;
assign x_1129 = v_4262 | ~v_3541;
assign x_1130 = v_4262 | ~v_2041;
assign x_1131 = v_4262 | ~v_2042;
assign x_1132 = v_4262 | ~v_2043;
assign x_1133 = v_4262 | ~v_2044;
assign x_1134 = v_4262 | ~v_3574;
assign x_1135 = v_4262 | ~v_3575;
assign x_1136 = v_4262 | ~v_3576;
assign x_1137 = v_4262 | ~v_3577;
assign x_1138 = v_4262 | ~v_2183;
assign x_1139 = v_4262 | ~v_2184;
assign x_1140 = v_4262 | ~v_2185;
assign x_1141 = v_4262 | ~v_2186;
assign x_1142 = v_4262 | ~v_3466;
assign x_1143 = v_4262 | ~v_3469;
assign x_1144 = v_4262 | ~v_2045;
assign x_1145 = v_4262 | ~v_4206;
assign x_1146 = v_4262 | ~v_4207;
assign x_1147 = v_4262 | ~v_2048;
assign x_1148 = v_4262 | ~v_4208;
assign x_1149 = v_4262 | ~v_4209;
assign x_1150 = v_4262 | ~v_771;
assign x_1151 = v_4262 | ~v_772;
assign x_1152 = v_4262 | ~v_1051;
assign x_1153 = v_4262 | ~v_1052;
assign x_1154 = v_4262 | ~v_1053;
assign x_1155 = v_4262 | ~v_1054;
assign x_1156 = v_4262 | ~v_1055;
assign x_1157 = v_4262 | ~v_1056;
assign x_1158 = v_4262 | ~v_182;
assign x_1159 = v_4262 | ~v_163;
assign x_1160 = v_4262 | ~v_162;
assign x_1161 = v_4262 | ~v_155;
assign x_1162 = v_4262 | ~v_137;
assign x_1163 = v_4262 | ~v_136;
assign x_1164 = v_4262 | ~v_135;
assign x_1165 = v_4262 | ~v_134;
assign x_1166 = v_4262 | ~v_18;
assign x_1167 = v_4262 | ~v_17;
assign x_1168 = v_4262 | ~v_15;
assign x_1169 = v_4262 | ~v_8;
assign x_1170 = ~v_4260 | ~v_4259 | ~v_4258 | v_4261;
assign x_1171 = v_4260 | ~v_3532;
assign x_1172 = v_4260 | ~v_3533;
assign x_1173 = v_4260 | ~v_3534;
assign x_1174 = v_4260 | ~v_3535;
assign x_1175 = v_4260 | ~v_2125;
assign x_1176 = v_4260 | ~v_2126;
assign x_1177 = v_4260 | ~v_2127;
assign x_1178 = v_4260 | ~v_2128;
assign x_1179 = v_4260 | ~v_3496;
assign x_1180 = v_4260 | ~v_3497;
assign x_1181 = v_4260 | ~v_3498;
assign x_1182 = v_4260 | ~v_3499;
assign x_1183 = v_4260 | ~v_3500;
assign x_1184 = v_4260 | ~v_3501;
assign x_1185 = v_4260 | ~v_2075;
assign x_1186 = v_4260 | ~v_4216;
assign x_1187 = v_4260 | ~v_2076;
assign x_1188 = v_4260 | ~v_4217;
assign x_1189 = v_4260 | ~v_2077;
assign x_1190 = v_4260 | ~v_2078;
assign x_1191 = v_4260 | ~v_4218;
assign x_1192 = v_4260 | ~v_2079;
assign x_1193 = v_4260 | ~v_4219;
assign x_1194 = v_4260 | ~v_2080;
assign x_1195 = v_4260 | ~v_1037;
assign x_1196 = v_4260 | ~v_1038;
assign x_1197 = v_4260 | ~v_1039;
assign x_1198 = v_4260 | ~v_1040;
assign x_1199 = v_4260 | ~v_927;
assign x_1200 = v_4260 | ~v_928;
assign x_1201 = v_4260 | ~v_839;
assign x_1202 = v_4260 | ~v_840;
assign x_1203 = v_4260 | ~v_184;
assign x_1204 = v_4260 | ~v_169;
assign x_1205 = v_4260 | ~v_151;
assign x_1206 = v_4260 | ~v_150;
assign x_1207 = v_4260 | ~v_149;
assign x_1208 = v_4260 | ~v_147;
assign x_1209 = v_4260 | ~v_103;
assign x_1210 = v_4260 | ~v_101;
assign x_1211 = v_4260 | ~v_100;
assign x_1212 = v_4260 | ~v_98;
assign x_1213 = v_4260 | ~v_96;
assign x_1214 = v_4260 | ~v_94;
assign x_1215 = v_4259 | ~v_3527;
assign x_1216 = v_4259 | ~v_3528;
assign x_1217 = v_4259 | ~v_3529;
assign x_1218 = v_4259 | ~v_3530;
assign x_1219 = v_4259 | ~v_2120;
assign x_1220 = v_4259 | ~v_2121;
assign x_1221 = v_4259 | ~v_2122;
assign x_1222 = v_4259 | ~v_2123;
assign x_1223 = v_4259 | ~v_3481;
assign x_1224 = v_4259 | ~v_3482;
assign x_1225 = v_4259 | ~v_3483;
assign x_1226 = v_4259 | ~v_3484;
assign x_1227 = v_4259 | ~v_3485;
assign x_1228 = v_4259 | ~v_2060;
assign x_1229 = v_4259 | ~v_4211;
assign x_1230 = v_4259 | ~v_2061;
assign x_1231 = v_4259 | ~v_4212;
assign x_1232 = v_4259 | ~v_2062;
assign x_1233 = v_4259 | ~v_2063;
assign x_1234 = v_4259 | ~v_4213;
assign x_1235 = v_4259 | ~v_2064;
assign x_1236 = v_4259 | ~v_4214;
assign x_1237 = v_4259 | ~v_2065;
assign x_1238 = v_4259 | ~v_1032;
assign x_1239 = v_4259 | ~v_1033;
assign x_1240 = v_4259 | ~v_1034;
assign x_1241 = v_4259 | ~v_1035;
assign x_1242 = v_4259 | ~v_912;
assign x_1243 = v_4259 | ~v_913;
assign x_1244 = v_4259 | ~v_806;
assign x_1245 = v_4259 | ~v_807;
assign x_1246 = v_4259 | ~v_3486;
assign x_1247 = v_4259 | ~v_183;
assign x_1248 = v_4259 | ~v_165;
assign x_1249 = v_4259 | ~v_146;
assign x_1250 = v_4259 | ~v_145;
assign x_1251 = v_4259 | ~v_144;
assign x_1252 = v_4259 | ~v_142;
assign x_1253 = v_4259 | ~v_61;
assign x_1254 = v_4259 | ~v_59;
assign x_1255 = v_4259 | ~v_58;
assign x_1256 = v_4259 | ~v_56;
assign x_1257 = v_4259 | ~v_54;
assign x_1258 = v_4259 | ~v_52;
assign x_1259 = v_4258 | ~v_3522;
assign x_1260 = v_4258 | ~v_3523;
assign x_1261 = v_4258 | ~v_3524;
assign x_1262 = v_4258 | ~v_3525;
assign x_1263 = v_4258 | ~v_2115;
assign x_1264 = v_4258 | ~v_2116;
assign x_1265 = v_4258 | ~v_2117;
assign x_1266 = v_4258 | ~v_2118;
assign x_1267 = v_4258 | ~v_3466;
assign x_1268 = v_4258 | ~v_3467;
assign x_1269 = v_4258 | ~v_3468;
assign x_1270 = v_4258 | ~v_3469;
assign x_1271 = v_4258 | ~v_3470;
assign x_1272 = v_4258 | ~v_2045;
assign x_1273 = v_4258 | ~v_4206;
assign x_1274 = v_4258 | ~v_2046;
assign x_1275 = v_4258 | ~v_4207;
assign x_1276 = v_4258 | ~v_2047;
assign x_1277 = v_4258 | ~v_2048;
assign x_1278 = v_4258 | ~v_4208;
assign x_1279 = v_4258 | ~v_2049;
assign x_1280 = v_4258 | ~v_4209;
assign x_1281 = v_4258 | ~v_2050;
assign x_1282 = v_4258 | ~v_1027;
assign x_1283 = v_4258 | ~v_1028;
assign x_1284 = v_4258 | ~v_1029;
assign x_1285 = v_4258 | ~v_1030;
assign x_1286 = v_4258 | ~v_897;
assign x_1287 = v_4258 | ~v_898;
assign x_1288 = v_4258 | ~v_773;
assign x_1289 = v_4258 | ~v_774;
assign x_1290 = v_4258 | ~v_182;
assign x_1291 = v_4258 | ~v_161;
assign x_1292 = v_4258 | ~v_138;
assign x_1293 = v_4258 | ~v_137;
assign x_1294 = v_4258 | ~v_3473;
assign x_1295 = v_4258 | ~v_136;
assign x_1296 = v_4258 | ~v_134;
assign x_1297 = v_4258 | ~v_18;
assign x_1298 = v_4258 | ~v_16;
assign x_1299 = v_4258 | ~v_15;
assign x_1300 = v_4258 | ~v_13;
assign x_1301 = v_4258 | ~v_11;
assign x_1302 = v_4258 | ~v_9;
assign x_1303 = ~v_4256 | ~v_4255 | ~v_4254 | v_4257;
assign x_1304 = v_4256 | ~v_3516;
assign x_1305 = v_4256 | ~v_3517;
assign x_1306 = v_4256 | ~v_3518;
assign x_1307 = v_4256 | ~v_3519;
assign x_1308 = v_4256 | ~v_2161;
assign x_1309 = v_4256 | ~v_2162;
assign x_1310 = v_4256 | ~v_2163;
assign x_1311 = v_4256 | ~v_2164;
assign x_1312 = v_4256 | ~v_3496;
assign x_1313 = v_4256 | ~v_3564;
assign x_1314 = v_4256 | ~v_3565;
assign x_1315 = v_4256 | ~v_3499;
assign x_1316 = v_4256 | ~v_3566;
assign x_1317 = v_4256 | ~v_3567;
assign x_1318 = v_4256 | ~v_2075;
assign x_1319 = v_4256 | ~v_4216;
assign x_1320 = v_4256 | ~v_2141;
assign x_1321 = v_4256 | ~v_4217;
assign x_1322 = v_4256 | ~v_2142;
assign x_1323 = v_4256 | ~v_2078;
assign x_1324 = v_4256 | ~v_4218;
assign x_1325 = v_4256 | ~v_2143;
assign x_1326 = v_4256 | ~v_4219;
assign x_1327 = v_4256 | ~v_2144;
assign x_1328 = v_4256 | ~v_1193;
assign x_1329 = v_4256 | ~v_1241;
assign x_1330 = v_4256 | ~v_1194;
assign x_1331 = v_4256 | ~v_1242;
assign x_1332 = v_4256 | ~v_1023;
assign x_1333 = v_4256 | ~v_1024;
assign x_1334 = v_4256 | ~v_1243;
assign x_1335 = v_4256 | ~v_1244;
assign x_1336 = v_4256 | ~v_184;
assign x_1337 = v_4256 | ~v_171;
assign x_1338 = v_4256 | ~v_170;
assign x_1339 = v_4256 | ~v_169;
assign x_1340 = v_4256 | ~v_148;
assign x_1341 = v_4256 | ~v_147;
assign x_1342 = v_4256 | ~v_103;
assign x_1343 = v_4256 | ~v_102;
assign x_1344 = v_4256 | ~v_101;
assign x_1345 = v_4256 | ~v_100;
assign x_1346 = v_4256 | ~v_99;
assign x_1347 = v_4256 | ~v_97;
assign x_1348 = v_4255 | ~v_3511;
assign x_1349 = v_4255 | ~v_3512;
assign x_1350 = v_4255 | ~v_3513;
assign x_1351 = v_4255 | ~v_3514;
assign x_1352 = v_4255 | ~v_2156;
assign x_1353 = v_4255 | ~v_2157;
assign x_1354 = v_4255 | ~v_2158;
assign x_1355 = v_4255 | ~v_2159;
assign x_1356 = v_4255 | ~v_3481;
assign x_1357 = v_4255 | ~v_3559;
assign x_1358 = v_4255 | ~v_3560;
assign x_1359 = v_4255 | ~v_3484;
assign x_1360 = v_4255 | ~v_2060;
assign x_1361 = v_4255 | ~v_4211;
assign x_1362 = v_4255 | ~v_2136;
assign x_1363 = v_4255 | ~v_4212;
assign x_1364 = v_4255 | ~v_2137;
assign x_1365 = v_4255 | ~v_2063;
assign x_1366 = v_4255 | ~v_4213;
assign x_1367 = v_4255 | ~v_2138;
assign x_1368 = v_4255 | ~v_4214;
assign x_1369 = v_4255 | ~v_2139;
assign x_1370 = v_4255 | ~v_1178;
assign x_1371 = v_4255 | ~v_1236;
assign x_1372 = v_4255 | ~v_1179;
assign x_1373 = v_4255 | ~v_1237;
assign x_1374 = v_4255 | ~v_1008;
assign x_1375 = v_4255 | ~v_1009;
assign x_1376 = v_4255 | ~v_3561;
assign x_1377 = v_4255 | ~v_3562;
assign x_1378 = v_4255 | ~v_1238;
assign x_1379 = v_4255 | ~v_1239;
assign x_1380 = v_4255 | ~v_183;
assign x_1381 = v_4255 | ~v_167;
assign x_1382 = v_4255 | ~v_166;
assign x_1383 = v_4255 | ~v_165;
assign x_1384 = v_4255 | ~v_143;
assign x_1385 = v_4255 | ~v_142;
assign x_1386 = v_4255 | ~v_61;
assign x_1387 = v_4255 | ~v_60;
assign x_1388 = v_4255 | ~v_59;
assign x_1389 = v_4255 | ~v_58;
assign x_1390 = v_4255 | ~v_57;
assign x_1391 = v_4255 | ~v_55;
assign x_1392 = v_4254 | ~v_3506;
assign x_1393 = v_4254 | ~v_3507;
assign x_1394 = v_4254 | ~v_3508;
assign x_1395 = v_4254 | ~v_3509;
assign x_1396 = v_4254 | ~v_2151;
assign x_1397 = v_4254 | ~v_2152;
assign x_1398 = v_4254 | ~v_2153;
assign x_1399 = v_4254 | ~v_2154;
assign x_1400 = v_4254 | ~v_3466;
assign x_1401 = v_4254 | ~v_3554;
assign x_1402 = v_4254 | ~v_3555;
assign x_1403 = v_4254 | ~v_3469;
assign x_1404 = v_4254 | ~v_3556;
assign x_1405 = v_4254 | ~v_3557;
assign x_1406 = v_4254 | ~v_2045;
assign x_1407 = v_4254 | ~v_4206;
assign x_1408 = v_4254 | ~v_2131;
assign x_1409 = v_4254 | ~v_4207;
assign x_1410 = v_4254 | ~v_2132;
assign x_1411 = v_4254 | ~v_2048;
assign x_1412 = v_4254 | ~v_4208;
assign x_1413 = v_4254 | ~v_2133;
assign x_1414 = v_4254 | ~v_4209;
assign x_1415 = v_4254 | ~v_2134;
assign x_1416 = v_4254 | ~v_1163;
assign x_1417 = v_4254 | ~v_1231;
assign x_1418 = v_4254 | ~v_1164;
assign x_1419 = v_4254 | ~v_1232;
assign x_1420 = v_4254 | ~v_1233;
assign x_1421 = v_4254 | ~v_1234;
assign x_1422 = v_4254 | ~v_182;
assign x_1423 = v_4254 | ~v_163;
assign x_1424 = v_4254 | ~v_162;
assign x_1425 = v_4254 | ~v_161;
assign x_1426 = v_4254 | ~v_135;
assign x_1427 = v_4254 | ~v_134;
assign x_1428 = v_4254 | ~v_993;
assign x_1429 = v_4254 | ~v_994;
assign x_1430 = v_4254 | ~v_18;
assign x_1431 = v_4254 | ~v_17;
assign x_1432 = v_4254 | ~v_16;
assign x_1433 = v_4254 | ~v_15;
assign x_1434 = v_4254 | ~v_14;
assign x_1435 = v_4254 | ~v_12;
assign x_1436 = ~v_4252 | ~v_4251 | ~v_4250 | v_4253;
assign x_1437 = v_4252 | ~v_3516;
assign x_1438 = v_4252 | ~v_3517;
assign x_1439 = v_4252 | ~v_3518;
assign x_1440 = v_4252 | ~v_3519;
assign x_1441 = v_4252 | ~v_2161;
assign x_1442 = v_4252 | ~v_2162;
assign x_1443 = v_4252 | ~v_2163;
assign x_1444 = v_4252 | ~v_2164;
assign x_1445 = v_4252 | ~v_3532;
assign x_1446 = v_4252 | ~v_3533;
assign x_1447 = v_4252 | ~v_3534;
assign x_1448 = v_4252 | ~v_3535;
assign x_1449 = v_4252 | ~v_2125;
assign x_1450 = v_4252 | ~v_2126;
assign x_1451 = v_4252 | ~v_2127;
assign x_1452 = v_4252 | ~v_2128;
assign x_1453 = v_4252 | ~v_3496;
assign x_1454 = v_4252 | ~v_3499;
assign x_1455 = v_4252 | ~v_2075;
assign x_1456 = v_4252 | ~v_4216;
assign x_1457 = v_4252 | ~v_4217;
assign x_1458 = v_4252 | ~v_2078;
assign x_1459 = v_4252 | ~v_4218;
assign x_1460 = v_4252 | ~v_4219;
assign x_1461 = v_4252 | ~v_1209;
assign x_1462 = v_4252 | ~v_1210;
assign x_1463 = v_4252 | ~v_1193;
assign x_1464 = v_4252 | ~v_1194;
assign x_1465 = v_4252 | ~v_927;
assign x_1466 = v_4252 | ~v_928;
assign x_1467 = v_4252 | ~v_1211;
assign x_1468 = v_4252 | ~v_1212;
assign x_1469 = v_4252 | ~v_184;
assign x_1470 = v_4252 | ~v_172;
assign x_1471 = v_4252 | ~v_171;
assign x_1472 = v_4252 | ~v_170;
assign x_1473 = v_4252 | ~v_169;
assign x_1474 = v_4252 | ~v_150;
assign x_1475 = v_4252 | ~v_149;
assign x_1476 = v_4252 | ~v_147;
assign x_1477 = v_4252 | ~v_102;
assign x_1478 = v_4252 | ~v_101;
assign x_1479 = v_4252 | ~v_100;
assign x_1480 = v_4252 | ~v_96;
assign x_1481 = v_4251 | ~v_3511;
assign x_1482 = v_4251 | ~v_3512;
assign x_1483 = v_4251 | ~v_3513;
assign x_1484 = v_4251 | ~v_3514;
assign x_1485 = v_4251 | ~v_2156;
assign x_1486 = v_4251 | ~v_2157;
assign x_1487 = v_4251 | ~v_2158;
assign x_1488 = v_4251 | ~v_2159;
assign x_1489 = v_4251 | ~v_3527;
assign x_1490 = v_4251 | ~v_3528;
assign x_1491 = v_4251 | ~v_3529;
assign x_1492 = v_4251 | ~v_3530;
assign x_1493 = v_4251 | ~v_2120;
assign x_1494 = v_4251 | ~v_2121;
assign x_1495 = v_4251 | ~v_2122;
assign x_1496 = v_4251 | ~v_2123;
assign x_1497 = v_4251 | ~v_3481;
assign x_1498 = v_4251 | ~v_3484;
assign x_1499 = v_4251 | ~v_2060;
assign x_1500 = v_4251 | ~v_4211;
assign x_1501 = v_4251 | ~v_4212;
assign x_1502 = v_4251 | ~v_2063;
assign x_1503 = v_4251 | ~v_4213;
assign x_1504 = v_4251 | ~v_4214;
assign x_1505 = v_4251 | ~v_1204;
assign x_1506 = v_4251 | ~v_1205;
assign x_1507 = v_4251 | ~v_1178;
assign x_1508 = v_4251 | ~v_1179;
assign x_1509 = v_4251 | ~v_912;
assign x_1510 = v_4251 | ~v_913;
assign x_1511 = v_4251 | ~v_1206;
assign x_1512 = v_4251 | ~v_1207;
assign x_1513 = v_4251 | ~v_183;
assign x_1514 = v_4251 | ~v_168;
assign x_1515 = v_4251 | ~v_167;
assign x_1516 = v_4251 | ~v_166;
assign x_1517 = v_4251 | ~v_165;
assign x_1518 = v_4251 | ~v_145;
assign x_1519 = v_4251 | ~v_144;
assign x_1520 = v_4251 | ~v_142;
assign x_1521 = v_4251 | ~v_60;
assign x_1522 = v_4251 | ~v_59;
assign x_1523 = v_4251 | ~v_58;
assign x_1524 = v_4251 | ~v_54;
assign x_1525 = v_4250 | ~v_3506;
assign x_1526 = v_4250 | ~v_3507;
assign x_1527 = v_4250 | ~v_3508;
assign x_1528 = v_4250 | ~v_3509;
assign x_1529 = v_4250 | ~v_2151;
assign x_1530 = v_4250 | ~v_2152;
assign x_1531 = v_4250 | ~v_2153;
assign x_1532 = v_4250 | ~v_2154;
assign x_1533 = v_4250 | ~v_3522;
assign x_1534 = v_4250 | ~v_3523;
assign x_1535 = v_4250 | ~v_3524;
assign x_1536 = v_4250 | ~v_3525;
assign x_1537 = v_4250 | ~v_2115;
assign x_1538 = v_4250 | ~v_2116;
assign x_1539 = v_4250 | ~v_2117;
assign x_1540 = v_4250 | ~v_2118;
assign x_1541 = v_4250 | ~v_3466;
assign x_1542 = v_4250 | ~v_3469;
assign x_1543 = v_4250 | ~v_2045;
assign x_1544 = v_4250 | ~v_4206;
assign x_1545 = v_4250 | ~v_4207;
assign x_1546 = v_4250 | ~v_2048;
assign x_1547 = v_4250 | ~v_4208;
assign x_1548 = v_4250 | ~v_4209;
assign x_1549 = v_4250 | ~v_1199;
assign x_1550 = v_4250 | ~v_1200;
assign x_1551 = v_4250 | ~v_1163;
assign x_1552 = v_4250 | ~v_1164;
assign x_1553 = v_4250 | ~v_897;
assign x_1554 = v_4250 | ~v_898;
assign x_1555 = v_4250 | ~v_1201;
assign x_1556 = v_4250 | ~v_1202;
assign x_1557 = v_4250 | ~v_182;
assign x_1558 = v_4250 | ~v_164;
assign x_1559 = v_4250 | ~v_163;
assign x_1560 = v_4250 | ~v_162;
assign x_1561 = v_4250 | ~v_161;
assign x_1562 = v_4250 | ~v_137;
assign x_1563 = v_4250 | ~v_136;
assign x_1564 = v_4250 | ~v_134;
assign x_1565 = v_4250 | ~v_17;
assign x_1566 = v_4250 | ~v_16;
assign x_1567 = v_4250 | ~v_15;
assign x_1568 = v_4250 | ~v_11;
assign x_1569 = ~v_4248 | ~v_4247 | ~v_4246 | v_4249;
assign x_1570 = v_4248 | ~v_3516;
assign x_1571 = v_4248 | ~v_3517;
assign x_1572 = v_4248 | ~v_3518;
assign x_1573 = v_4248 | ~v_3519;
assign x_1574 = v_4248 | ~v_2161;
assign x_1575 = v_4248 | ~v_2162;
assign x_1576 = v_4248 | ~v_2163;
assign x_1577 = v_4248 | ~v_2164;
assign x_1578 = v_4248 | ~v_3494;
assign x_1579 = v_4248 | ~v_3495;
assign x_1580 = v_4248 | ~v_2109;
assign x_1581 = v_4248 | ~v_2110;
assign x_1582 = v_4248 | ~v_2111;
assign x_1583 = v_4248 | ~v_2112;
assign x_1584 = v_4248 | ~v_3496;
assign x_1585 = v_4248 | ~v_3499;
assign x_1586 = v_4248 | ~v_2075;
assign x_1587 = v_4248 | ~v_4216;
assign x_1588 = v_4248 | ~v_4217;
assign x_1589 = v_4248 | ~v_2078;
assign x_1590 = v_4248 | ~v_4218;
assign x_1591 = v_4248 | ~v_4219;
assign x_1592 = v_4248 | ~v_1225;
assign x_1593 = v_4248 | ~v_1226;
assign x_1594 = v_4248 | ~v_1227;
assign x_1595 = v_4248 | ~v_1228;
assign x_1596 = v_4248 | ~v_1193;
assign x_1597 = v_4248 | ~v_1194;
assign x_1598 = v_4248 | ~v_975;
assign x_1599 = v_4248 | ~v_976;
assign x_1600 = v_4248 | ~v_3502;
assign x_1601 = v_4248 | ~v_3503;
assign x_1602 = v_4248 | ~v_184;
assign x_1603 = v_4248 | ~v_171;
assign x_1604 = v_4248 | ~v_170;
assign x_1605 = v_4248 | ~v_169;
assign x_1606 = v_4248 | ~v_150;
assign x_1607 = v_4248 | ~v_149;
assign x_1608 = v_4248 | ~v_148;
assign x_1609 = v_4248 | ~v_103;
assign x_1610 = v_4248 | ~v_102;
assign x_1611 = v_4248 | ~v_101;
assign x_1612 = v_4248 | ~v_100;
assign x_1613 = v_4248 | ~v_95;
assign x_1614 = v_4247 | ~v_3511;
assign x_1615 = v_4247 | ~v_3512;
assign x_1616 = v_4247 | ~v_3513;
assign x_1617 = v_4247 | ~v_3514;
assign x_1618 = v_4247 | ~v_2156;
assign x_1619 = v_4247 | ~v_2157;
assign x_1620 = v_4247 | ~v_2158;
assign x_1621 = v_4247 | ~v_2159;
assign x_1622 = v_4247 | ~v_3479;
assign x_1623 = v_4247 | ~v_3480;
assign x_1624 = v_4247 | ~v_2104;
assign x_1625 = v_4247 | ~v_2105;
assign x_1626 = v_4247 | ~v_2106;
assign x_1627 = v_4247 | ~v_2107;
assign x_1628 = v_4247 | ~v_3481;
assign x_1629 = v_4247 | ~v_3484;
assign x_1630 = v_4247 | ~v_2060;
assign x_1631 = v_4247 | ~v_4211;
assign x_1632 = v_4247 | ~v_4212;
assign x_1633 = v_4247 | ~v_2063;
assign x_1634 = v_4247 | ~v_4213;
assign x_1635 = v_4247 | ~v_4214;
assign x_1636 = v_4247 | ~v_1220;
assign x_1637 = v_4247 | ~v_1221;
assign x_1638 = v_4247 | ~v_1222;
assign x_1639 = v_4247 | ~v_1223;
assign x_1640 = v_4247 | ~v_1178;
assign x_1641 = v_4247 | ~v_1179;
assign x_1642 = v_4247 | ~v_960;
assign x_1643 = v_4247 | ~v_961;
assign x_1644 = v_4247 | ~v_3487;
assign x_1645 = v_4247 | ~v_3488;
assign x_1646 = v_4247 | ~v_183;
assign x_1647 = v_4247 | ~v_167;
assign x_1648 = v_4247 | ~v_166;
assign x_1649 = v_4247 | ~v_165;
assign x_1650 = v_4247 | ~v_145;
assign x_1651 = v_4247 | ~v_144;
assign x_1652 = v_4247 | ~v_143;
assign x_1653 = v_4247 | ~v_61;
assign x_1654 = v_4247 | ~v_60;
assign x_1655 = v_4247 | ~v_59;
assign x_1656 = v_4247 | ~v_58;
assign x_1657 = v_4247 | ~v_53;
assign x_1658 = v_4246 | ~v_3506;
assign x_1659 = v_4246 | ~v_3507;
assign x_1660 = v_4246 | ~v_3508;
assign x_1661 = v_4246 | ~v_3509;
assign x_1662 = v_4246 | ~v_2151;
assign x_1663 = v_4246 | ~v_2152;
assign x_1664 = v_4246 | ~v_2153;
assign x_1665 = v_4246 | ~v_2154;
assign x_1666 = v_4246 | ~v_3464;
assign x_1667 = v_4246 | ~v_3465;
assign x_1668 = v_4246 | ~v_2099;
assign x_1669 = v_4246 | ~v_2100;
assign x_1670 = v_4246 | ~v_2101;
assign x_1671 = v_4246 | ~v_2102;
assign x_1672 = v_4246 | ~v_3466;
assign x_1673 = v_4246 | ~v_3469;
assign x_1674 = v_4246 | ~v_2045;
assign x_1675 = v_4246 | ~v_4206;
assign x_1676 = v_4246 | ~v_4207;
assign x_1677 = v_4246 | ~v_2048;
assign x_1678 = v_4246 | ~v_4208;
assign x_1679 = v_4246 | ~v_4209;
assign x_1680 = v_4246 | ~v_1215;
assign x_1681 = v_4246 | ~v_1216;
assign x_1682 = v_4246 | ~v_1217;
assign x_1683 = v_4246 | ~v_1218;
assign x_1684 = v_4246 | ~v_1163;
assign x_1685 = v_4246 | ~v_1164;
assign x_1686 = v_4246 | ~v_945;
assign x_1687 = v_4246 | ~v_946;
assign x_1688 = v_4246 | ~v_3471;
assign x_1689 = v_4246 | ~v_3472;
assign x_1690 = v_4246 | ~v_182;
assign x_1691 = v_4246 | ~v_163;
assign x_1692 = v_4246 | ~v_162;
assign x_1693 = v_4246 | ~v_161;
assign x_1694 = v_4246 | ~v_137;
assign x_1695 = v_4246 | ~v_136;
assign x_1696 = v_4246 | ~v_135;
assign x_1697 = v_4246 | ~v_18;
assign x_1698 = v_4246 | ~v_17;
assign x_1699 = v_4246 | ~v_16;
assign x_1700 = v_4246 | ~v_15;
assign x_1701 = v_4246 | ~v_10;
assign x_1702 = ~v_4244 | ~v_4243 | ~v_4242 | v_4245;
assign x_1703 = v_4244 | ~v_3516;
assign x_1704 = v_4244 | ~v_3517;
assign x_1705 = v_4244 | ~v_3518;
assign x_1706 = v_4244 | ~v_3519;
assign x_1707 = v_4244 | ~v_2161;
assign x_1708 = v_4244 | ~v_2162;
assign x_1709 = v_4244 | ~v_2163;
assign x_1710 = v_4244 | ~v_2164;
assign x_1711 = v_4244 | ~v_3548;
assign x_1712 = v_4244 | ~v_3549;
assign x_1713 = v_4244 | ~v_3550;
assign x_1714 = v_4244 | ~v_3551;
assign x_1715 = v_4244 | ~v_2071;
assign x_1716 = v_4244 | ~v_2072;
assign x_1717 = v_4244 | ~v_2073;
assign x_1718 = v_4244 | ~v_2074;
assign x_1719 = v_4244 | ~v_3496;
assign x_1720 = v_4244 | ~v_3499;
assign x_1721 = v_4244 | ~v_2075;
assign x_1722 = v_4244 | ~v_4216;
assign x_1723 = v_4244 | ~v_4217;
assign x_1724 = v_4244 | ~v_2078;
assign x_1725 = v_4244 | ~v_4218;
assign x_1726 = v_4244 | ~v_4219;
assign x_1727 = v_4244 | ~v_1191;
assign x_1728 = v_4244 | ~v_1192;
assign x_1729 = v_4244 | ~v_1193;
assign x_1730 = v_4244 | ~v_1194;
assign x_1731 = v_4244 | ~v_837;
assign x_1732 = v_4244 | ~v_838;
assign x_1733 = v_4244 | ~v_1195;
assign x_1734 = v_4244 | ~v_1196;
assign x_1735 = v_4244 | ~v_184;
assign x_1736 = v_4244 | ~v_171;
assign x_1737 = v_4244 | ~v_170;
assign x_1738 = v_4244 | ~v_169;
assign x_1739 = v_4244 | ~v_160;
assign x_1740 = v_4244 | ~v_151;
assign x_1741 = v_4244 | ~v_150;
assign x_1742 = v_4244 | ~v_149;
assign x_1743 = v_4244 | ~v_148;
assign x_1744 = v_4244 | ~v_147;
assign x_1745 = v_4244 | ~v_103;
assign x_1746 = v_4244 | ~v_100;
assign x_1747 = v_4243 | ~v_3511;
assign x_1748 = v_4243 | ~v_3512;
assign x_1749 = v_4243 | ~v_3513;
assign x_1750 = v_4243 | ~v_3514;
assign x_1751 = v_4243 | ~v_2156;
assign x_1752 = v_4243 | ~v_2157;
assign x_1753 = v_4243 | ~v_2158;
assign x_1754 = v_4243 | ~v_2159;
assign x_1755 = v_4243 | ~v_3543;
assign x_1756 = v_4243 | ~v_3544;
assign x_1757 = v_4243 | ~v_3545;
assign x_1758 = v_4243 | ~v_3546;
assign x_1759 = v_4243 | ~v_2056;
assign x_1760 = v_4243 | ~v_2057;
assign x_1761 = v_4243 | ~v_2058;
assign x_1762 = v_4243 | ~v_2059;
assign x_1763 = v_4243 | ~v_3481;
assign x_1764 = v_4243 | ~v_3484;
assign x_1765 = v_4243 | ~v_2060;
assign x_1766 = v_4243 | ~v_4211;
assign x_1767 = v_4243 | ~v_4212;
assign x_1768 = v_4243 | ~v_2063;
assign x_1769 = v_4243 | ~v_4213;
assign x_1770 = v_4243 | ~v_4214;
assign x_1771 = v_4243 | ~v_1176;
assign x_1772 = v_4243 | ~v_1177;
assign x_1773 = v_4243 | ~v_1178;
assign x_1774 = v_4243 | ~v_1179;
assign x_1775 = v_4243 | ~v_804;
assign x_1776 = v_4243 | ~v_805;
assign x_1777 = v_4243 | ~v_1180;
assign x_1778 = v_4243 | ~v_1181;
assign x_1779 = v_4243 | ~v_183;
assign x_1780 = v_4243 | ~v_167;
assign x_1781 = v_4243 | ~v_166;
assign x_1782 = v_4243 | ~v_165;
assign x_1783 = v_4243 | ~v_159;
assign x_1784 = v_4243 | ~v_146;
assign x_1785 = v_4243 | ~v_145;
assign x_1786 = v_4243 | ~v_144;
assign x_1787 = v_4243 | ~v_143;
assign x_1788 = v_4243 | ~v_142;
assign x_1789 = v_4243 | ~v_61;
assign x_1790 = v_4243 | ~v_58;
assign x_1791 = v_4242 | ~v_3506;
assign x_1792 = v_4242 | ~v_3507;
assign x_1793 = v_4242 | ~v_3508;
assign x_1794 = v_4242 | ~v_3509;
assign x_1795 = v_4242 | ~v_2151;
assign x_1796 = v_4242 | ~v_2152;
assign x_1797 = v_4242 | ~v_2153;
assign x_1798 = v_4242 | ~v_2154;
assign x_1799 = v_4242 | ~v_3538;
assign x_1800 = v_4242 | ~v_3539;
assign x_1801 = v_4242 | ~v_3540;
assign x_1802 = v_4242 | ~v_3541;
assign x_1803 = v_4242 | ~v_2041;
assign x_1804 = v_4242 | ~v_2042;
assign x_1805 = v_4242 | ~v_2043;
assign x_1806 = v_4242 | ~v_2044;
assign x_1807 = v_4242 | ~v_3466;
assign x_1808 = v_4242 | ~v_3469;
assign x_1809 = v_4242 | ~v_2045;
assign x_1810 = v_4242 | ~v_4206;
assign x_1811 = v_4242 | ~v_4207;
assign x_1812 = v_4242 | ~v_2048;
assign x_1813 = v_4242 | ~v_4208;
assign x_1814 = v_4242 | ~v_4209;
assign x_1815 = v_4242 | ~v_1161;
assign x_1816 = v_4242 | ~v_1162;
assign x_1817 = v_4242 | ~v_1163;
assign x_1818 = v_4242 | ~v_1164;
assign x_1819 = v_4242 | ~v_771;
assign x_1820 = v_4242 | ~v_772;
assign x_1821 = v_4242 | ~v_1165;
assign x_1822 = v_4242 | ~v_1166;
assign x_1823 = v_4242 | ~v_182;
assign x_1824 = v_4242 | ~v_163;
assign x_1825 = v_4242 | ~v_162;
assign x_1826 = v_4242 | ~v_161;
assign x_1827 = v_4242 | ~v_155;
assign x_1828 = v_4242 | ~v_138;
assign x_1829 = v_4242 | ~v_137;
assign x_1830 = v_4242 | ~v_136;
assign x_1831 = v_4242 | ~v_135;
assign x_1832 = v_4242 | ~v_134;
assign x_1833 = v_4242 | ~v_18;
assign x_1834 = v_4242 | ~v_15;
assign x_1835 = ~v_4240 | ~v_4239 | ~v_4238 | v_4241;
assign x_1836 = v_4240 | ~v_3494;
assign x_1837 = v_4240 | ~v_3495;
assign x_1838 = v_4240 | ~v_2109;
assign x_1839 = v_4240 | ~v_2110;
assign x_1840 = v_4240 | ~v_2111;
assign x_1841 = v_4240 | ~v_2112;
assign x_1842 = v_4240 | ~v_3496;
assign x_1843 = v_4240 | ~v_3497;
assign x_1844 = v_4240 | ~v_3498;
assign x_1845 = v_4240 | ~v_3499;
assign x_1846 = v_4240 | ~v_3500;
assign x_1847 = v_4240 | ~v_3501;
assign x_1848 = v_4240 | ~v_2075;
assign x_1849 = v_4240 | ~v_4216;
assign x_1850 = v_4240 | ~v_2076;
assign x_1851 = v_4240 | ~v_4217;
assign x_1852 = v_4240 | ~v_2077;
assign x_1853 = v_4240 | ~v_2078;
assign x_1854 = v_4240 | ~v_4218;
assign x_1855 = v_4240 | ~v_2079;
assign x_1856 = v_4240 | ~v_4219;
assign x_1857 = v_4240 | ~v_2080;
assign x_1858 = v_4240 | ~v_1147;
assign x_1859 = v_4240 | ~v_1148;
assign x_1860 = v_4240 | ~v_975;
assign x_1861 = v_4240 | ~v_976;
assign x_1862 = v_4240 | ~v_839;
assign x_1863 = v_4240 | ~v_840;
assign x_1864 = v_4240 | ~v_1149;
assign x_1865 = v_4240 | ~v_1150;
assign x_1866 = v_4240 | ~v_3502;
assign x_1867 = v_4240 | ~v_3503;
assign x_1868 = v_4240 | ~v_184;
assign x_1869 = v_4240 | ~v_169;
assign x_1870 = v_4240 | ~v_150;
assign x_1871 = v_4240 | ~v_149;
assign x_1872 = v_4240 | ~v_148;
assign x_1873 = v_4240 | ~v_147;
assign x_1874 = v_4240 | ~v_103;
assign x_1875 = v_4240 | ~v_102;
assign x_1876 = v_4240 | ~v_101;
assign x_1877 = v_4240 | ~v_100;
assign x_1878 = v_4240 | ~v_98;
assign x_1879 = v_4240 | ~v_94;
assign x_1880 = v_4239 | ~v_3479;
assign x_1881 = v_4239 | ~v_3480;
assign x_1882 = v_4239 | ~v_2104;
assign x_1883 = v_4239 | ~v_2105;
assign x_1884 = v_4239 | ~v_2106;
assign x_1885 = v_4239 | ~v_2107;
assign x_1886 = v_4239 | ~v_3481;
assign x_1887 = v_4239 | ~v_3482;
assign x_1888 = v_4239 | ~v_3483;
assign x_1889 = v_4239 | ~v_3484;
assign x_1890 = v_4239 | ~v_3485;
assign x_1891 = v_4239 | ~v_2060;
assign x_1892 = v_4239 | ~v_4211;
assign x_1893 = v_4239 | ~v_2061;
assign x_1894 = v_4239 | ~v_4212;
assign x_1895 = v_4239 | ~v_2062;
assign x_1896 = v_4239 | ~v_2063;
assign x_1897 = v_4239 | ~v_4213;
assign x_1898 = v_4239 | ~v_2064;
assign x_1899 = v_4239 | ~v_4214;
assign x_1900 = v_4239 | ~v_2065;
assign x_1901 = v_4239 | ~v_1142;
assign x_1902 = v_4239 | ~v_1143;
assign x_1903 = v_4239 | ~v_960;
assign x_1904 = v_4239 | ~v_961;
assign x_1905 = v_4239 | ~v_806;
assign x_1906 = v_4239 | ~v_807;
assign x_1907 = v_4239 | ~v_3486;
assign x_1908 = v_4239 | ~v_1144;
assign x_1909 = v_4239 | ~v_1145;
assign x_1910 = v_4239 | ~v_3487;
assign x_1911 = v_4239 | ~v_3488;
assign x_1912 = v_4239 | ~v_183;
assign x_1913 = v_4239 | ~v_165;
assign x_1914 = v_4239 | ~v_145;
assign x_1915 = v_4239 | ~v_144;
assign x_1916 = v_4239 | ~v_143;
assign x_1917 = v_4239 | ~v_142;
assign x_1918 = v_4239 | ~v_61;
assign x_1919 = v_4239 | ~v_60;
assign x_1920 = v_4239 | ~v_59;
assign x_1921 = v_4239 | ~v_58;
assign x_1922 = v_4239 | ~v_56;
assign x_1923 = v_4239 | ~v_52;
assign x_1924 = v_4238 | ~v_3464;
assign x_1925 = v_4238 | ~v_3465;
assign x_1926 = v_4238 | ~v_2099;
assign x_1927 = v_4238 | ~v_2100;
assign x_1928 = v_4238 | ~v_2101;
assign x_1929 = v_4238 | ~v_2102;
assign x_1930 = v_4238 | ~v_3466;
assign x_1931 = v_4238 | ~v_3467;
assign x_1932 = v_4238 | ~v_3468;
assign x_1933 = v_4238 | ~v_3469;
assign x_1934 = v_4238 | ~v_3470;
assign x_1935 = v_4238 | ~v_2045;
assign x_1936 = v_4238 | ~v_4206;
assign x_1937 = v_4238 | ~v_2046;
assign x_1938 = v_4238 | ~v_4207;
assign x_1939 = v_4238 | ~v_2047;
assign x_1940 = v_4238 | ~v_2048;
assign x_1941 = v_4238 | ~v_4208;
assign x_1942 = v_4238 | ~v_2049;
assign x_1943 = v_4238 | ~v_4209;
assign x_1944 = v_4238 | ~v_2050;
assign x_1945 = v_4238 | ~v_1137;
assign x_1946 = v_4238 | ~v_1138;
assign x_1947 = v_4238 | ~v_945;
assign x_1948 = v_4238 | ~v_946;
assign x_1949 = v_4238 | ~v_773;
assign x_1950 = v_4238 | ~v_774;
assign x_1951 = v_4238 | ~v_1139;
assign x_1952 = v_4238 | ~v_1140;
assign x_1953 = v_4238 | ~v_3471;
assign x_1954 = v_4238 | ~v_3472;
assign x_1955 = v_4238 | ~v_182;
assign x_1956 = v_4238 | ~v_161;
assign x_1957 = v_4238 | ~v_137;
assign x_1958 = v_4238 | ~v_3473;
assign x_1959 = v_4238 | ~v_136;
assign x_1960 = v_4238 | ~v_135;
assign x_1961 = v_4238 | ~v_134;
assign x_1962 = v_4238 | ~v_18;
assign x_1963 = v_4238 | ~v_17;
assign x_1964 = v_4238 | ~v_16;
assign x_1965 = v_4238 | ~v_15;
assign x_1966 = v_4238 | ~v_13;
assign x_1967 = v_4238 | ~v_9;
assign x_1968 = ~v_4236 | ~v_4235 | ~v_4234 | v_4237;
assign x_1969 = v_4236 | ~v_3616;
assign x_1970 = v_4236 | ~v_3617;
assign x_1971 = v_4236 | ~v_3618;
assign x_1972 = v_4236 | ~v_3619;
assign x_1973 = v_4236 | ~v_2093;
assign x_1974 = v_4236 | ~v_2094;
assign x_1975 = v_4236 | ~v_2095;
assign x_1976 = v_4236 | ~v_2096;
assign x_1977 = v_4236 | ~v_3496;
assign x_1978 = v_4236 | ~v_3564;
assign x_1979 = v_4236 | ~v_3565;
assign x_1980 = v_4236 | ~v_3499;
assign x_1981 = v_4236 | ~v_3566;
assign x_1982 = v_4236 | ~v_3567;
assign x_1983 = v_4236 | ~v_2075;
assign x_1984 = v_4236 | ~v_4216;
assign x_1985 = v_4236 | ~v_2141;
assign x_1986 = v_4236 | ~v_4217;
assign x_1987 = v_4236 | ~v_2142;
assign x_1988 = v_4236 | ~v_2078;
assign x_1989 = v_4236 | ~v_4218;
assign x_1990 = v_4236 | ~v_2143;
assign x_1991 = v_4236 | ~v_4219;
assign x_1992 = v_4236 | ~v_2144;
assign x_1993 = v_4236 | ~v_885;
assign x_1994 = v_4236 | ~v_1019;
assign x_1995 = v_4236 | ~v_1020;
assign x_1996 = v_4236 | ~v_886;
assign x_1997 = v_4236 | ~v_1021;
assign x_1998 = v_4236 | ~v_1022;
assign x_1999 = v_4236 | ~v_1023;
assign x_2000 = v_4236 | ~v_1024;
assign x_2001 = v_4236 | ~v_184;
assign x_2002 = v_4236 | ~v_181;
assign x_2003 = v_4236 | ~v_171;
assign x_2004 = v_4236 | ~v_170;
assign x_2005 = v_4236 | ~v_169;
assign x_2006 = v_4236 | ~v_148;
assign x_2007 = v_4236 | ~v_147;
assign x_2008 = v_4236 | ~v_103;
assign x_2009 = v_4236 | ~v_102;
assign x_2010 = v_4236 | ~v_101;
assign x_2011 = v_4236 | ~v_99;
assign x_2012 = v_4236 | ~v_97;
assign x_2013 = v_4235 | ~v_3611;
assign x_2014 = v_4235 | ~v_3612;
assign x_2015 = v_4235 | ~v_3613;
assign x_2016 = v_4235 | ~v_3614;
assign x_2017 = v_4235 | ~v_2088;
assign x_2018 = v_4235 | ~v_2089;
assign x_2019 = v_4235 | ~v_2090;
assign x_2020 = v_4235 | ~v_2091;
assign x_2021 = v_4235 | ~v_3481;
assign x_2022 = v_4235 | ~v_3559;
assign x_2023 = v_4235 | ~v_3560;
assign x_2024 = v_4235 | ~v_3484;
assign x_2025 = v_4235 | ~v_2060;
assign x_2026 = v_4235 | ~v_4211;
assign x_2027 = v_4235 | ~v_2136;
assign x_2028 = v_4235 | ~v_4212;
assign x_2029 = v_4235 | ~v_2137;
assign x_2030 = v_4235 | ~v_2063;
assign x_2031 = v_4235 | ~v_4213;
assign x_2032 = v_4235 | ~v_2138;
assign x_2033 = v_4235 | ~v_4214;
assign x_2034 = v_4235 | ~v_2139;
assign x_2035 = v_4235 | ~v_870;
assign x_2036 = v_4235 | ~v_1004;
assign x_2037 = v_4235 | ~v_1005;
assign x_2038 = v_4235 | ~v_871;
assign x_2039 = v_4235 | ~v_1006;
assign x_2040 = v_4235 | ~v_1007;
assign x_2041 = v_4235 | ~v_1008;
assign x_2042 = v_4235 | ~v_1009;
assign x_2043 = v_4235 | ~v_3561;
assign x_2044 = v_4235 | ~v_3562;
assign x_2045 = v_4235 | ~v_183;
assign x_2046 = v_4235 | ~v_180;
assign x_2047 = v_4235 | ~v_167;
assign x_2048 = v_4235 | ~v_166;
assign x_2049 = v_4235 | ~v_165;
assign x_2050 = v_4235 | ~v_143;
assign x_2051 = v_4235 | ~v_142;
assign x_2052 = v_4235 | ~v_61;
assign x_2053 = v_4235 | ~v_60;
assign x_2054 = v_4235 | ~v_59;
assign x_2055 = v_4235 | ~v_57;
assign x_2056 = v_4235 | ~v_55;
assign x_2057 = v_4234 | ~v_3606;
assign x_2058 = v_4234 | ~v_3607;
assign x_2059 = v_4234 | ~v_3608;
assign x_2060 = v_4234 | ~v_3609;
assign x_2061 = v_4234 | ~v_2083;
assign x_2062 = v_4234 | ~v_2084;
assign x_2063 = v_4234 | ~v_2085;
assign x_2064 = v_4234 | ~v_2086;
assign x_2065 = v_4234 | ~v_3466;
assign x_2066 = v_4234 | ~v_3554;
assign x_2067 = v_4234 | ~v_3555;
assign x_2068 = v_4234 | ~v_3469;
assign x_2069 = v_4234 | ~v_3556;
assign x_2070 = v_4234 | ~v_3557;
assign x_2071 = v_4234 | ~v_2045;
assign x_2072 = v_4234 | ~v_4206;
assign x_2073 = v_4234 | ~v_2131;
assign x_2074 = v_4234 | ~v_4207;
assign x_2075 = v_4234 | ~v_2132;
assign x_2076 = v_4234 | ~v_2048;
assign x_2077 = v_4234 | ~v_4208;
assign x_2078 = v_4234 | ~v_2133;
assign x_2079 = v_4234 | ~v_4209;
assign x_2080 = v_4234 | ~v_2134;
assign x_2081 = v_4234 | ~v_855;
assign x_2082 = v_4234 | ~v_989;
assign x_2083 = v_4234 | ~v_990;
assign x_2084 = v_4234 | ~v_856;
assign x_2085 = v_4234 | ~v_991;
assign x_2086 = v_4234 | ~v_992;
assign x_2087 = v_4234 | ~v_182;
assign x_2088 = v_4234 | ~v_179;
assign x_2089 = v_4234 | ~v_163;
assign x_2090 = v_4234 | ~v_162;
assign x_2091 = v_4234 | ~v_161;
assign x_2092 = v_4234 | ~v_135;
assign x_2093 = v_4234 | ~v_134;
assign x_2094 = v_4234 | ~v_993;
assign x_2095 = v_4234 | ~v_994;
assign x_2096 = v_4234 | ~v_18;
assign x_2097 = v_4234 | ~v_17;
assign x_2098 = v_4234 | ~v_16;
assign x_2099 = v_4234 | ~v_14;
assign x_2100 = v_4234 | ~v_12;
assign x_2101 = ~v_4232 | ~v_4231 | ~v_4230 | v_4233;
assign x_2102 = v_4232 | ~v_3616;
assign x_2103 = v_4232 | ~v_3617;
assign x_2104 = v_4232 | ~v_3618;
assign x_2105 = v_4232 | ~v_3619;
assign x_2106 = v_4232 | ~v_2093;
assign x_2107 = v_4232 | ~v_2094;
assign x_2108 = v_4232 | ~v_2095;
assign x_2109 = v_4232 | ~v_2096;
assign x_2110 = v_4232 | ~v_3532;
assign x_2111 = v_4232 | ~v_3533;
assign x_2112 = v_4232 | ~v_3534;
assign x_2113 = v_4232 | ~v_3535;
assign x_2114 = v_4232 | ~v_2125;
assign x_2115 = v_4232 | ~v_2126;
assign x_2116 = v_4232 | ~v_2127;
assign x_2117 = v_4232 | ~v_2128;
assign x_2118 = v_4232 | ~v_3496;
assign x_2119 = v_4232 | ~v_3499;
assign x_2120 = v_4232 | ~v_2075;
assign x_2121 = v_4232 | ~v_4216;
assign x_2122 = v_4232 | ~v_4217;
assign x_2123 = v_4232 | ~v_2078;
assign x_2124 = v_4232 | ~v_4218;
assign x_2125 = v_4232 | ~v_4219;
assign x_2126 = v_4232 | ~v_925;
assign x_2127 = v_4232 | ~v_926;
assign x_2128 = v_4232 | ~v_885;
assign x_2129 = v_4232 | ~v_886;
assign x_2130 = v_4232 | ~v_927;
assign x_2131 = v_4232 | ~v_928;
assign x_2132 = v_4232 | ~v_929;
assign x_2133 = v_4232 | ~v_930;
assign x_2134 = v_4232 | ~v_184;
assign x_2135 = v_4232 | ~v_181;
assign x_2136 = v_4232 | ~v_171;
assign x_2137 = v_4232 | ~v_170;
assign x_2138 = v_4232 | ~v_169;
assign x_2139 = v_4232 | ~v_150;
assign x_2140 = v_4232 | ~v_149;
assign x_2141 = v_4232 | ~v_147;
assign x_2142 = v_4232 | ~v_103;
assign x_2143 = v_4232 | ~v_102;
assign x_2144 = v_4232 | ~v_101;
assign x_2145 = v_4232 | ~v_96;
assign x_2146 = v_4231 | ~v_3611;
assign x_2147 = v_4231 | ~v_3612;
assign x_2148 = v_4231 | ~v_3613;
assign x_2149 = v_4231 | ~v_3614;
assign x_2150 = v_4231 | ~v_2088;
assign x_2151 = v_4231 | ~v_2089;
assign x_2152 = v_4231 | ~v_2090;
assign x_2153 = v_4231 | ~v_2091;
assign x_2154 = v_4231 | ~v_3527;
assign x_2155 = v_4231 | ~v_3528;
assign x_2156 = v_4231 | ~v_3529;
assign x_2157 = v_4231 | ~v_3530;
assign x_2158 = v_4231 | ~v_2120;
assign x_2159 = v_4231 | ~v_2121;
assign x_2160 = v_4231 | ~v_2122;
assign x_2161 = v_4231 | ~v_2123;
assign x_2162 = v_4231 | ~v_3481;
assign x_2163 = v_4231 | ~v_3484;
assign x_2164 = v_4231 | ~v_2060;
assign x_2165 = v_4231 | ~v_4211;
assign x_2166 = v_4231 | ~v_4212;
assign x_2167 = v_4231 | ~v_2063;
assign x_2168 = v_4231 | ~v_4213;
assign x_2169 = v_4231 | ~v_4214;
assign x_2170 = v_4231 | ~v_910;
assign x_2171 = v_4231 | ~v_911;
assign x_2172 = v_4231 | ~v_870;
assign x_2173 = v_4231 | ~v_871;
assign x_2174 = v_4231 | ~v_912;
assign x_2175 = v_4231 | ~v_913;
assign x_2176 = v_4231 | ~v_914;
assign x_2177 = v_4231 | ~v_915;
assign x_2178 = v_4231 | ~v_183;
assign x_2179 = v_4231 | ~v_180;
assign x_2180 = v_4231 | ~v_167;
assign x_2181 = v_4231 | ~v_166;
assign x_2182 = v_4231 | ~v_165;
assign x_2183 = v_4231 | ~v_145;
assign x_2184 = v_4231 | ~v_144;
assign x_2185 = v_4231 | ~v_142;
assign x_2186 = v_4231 | ~v_61;
assign x_2187 = v_4231 | ~v_60;
assign x_2188 = v_4231 | ~v_59;
assign x_2189 = v_4231 | ~v_54;
assign x_2190 = v_4230 | ~v_3606;
assign x_2191 = v_4230 | ~v_3607;
assign x_2192 = v_4230 | ~v_3608;
assign x_2193 = v_4230 | ~v_3609;
assign x_2194 = v_4230 | ~v_2083;
assign x_2195 = v_4230 | ~v_2084;
assign x_2196 = v_4230 | ~v_2085;
assign x_2197 = v_4230 | ~v_2086;
assign x_2198 = v_4230 | ~v_3522;
assign x_2199 = v_4230 | ~v_3523;
assign x_2200 = v_4230 | ~v_3524;
assign x_2201 = v_4230 | ~v_3525;
assign x_2202 = v_4230 | ~v_2115;
assign x_2203 = v_4230 | ~v_2116;
assign x_2204 = v_4230 | ~v_2117;
assign x_2205 = v_4230 | ~v_2118;
assign x_2206 = v_4230 | ~v_3466;
assign x_2207 = v_4230 | ~v_3469;
assign x_2208 = v_4230 | ~v_2045;
assign x_2209 = v_4230 | ~v_4206;
assign x_2210 = v_4230 | ~v_4207;
assign x_2211 = v_4230 | ~v_2048;
assign x_2212 = v_4230 | ~v_4208;
assign x_2213 = v_4230 | ~v_4209;
assign x_2214 = v_4230 | ~v_895;
assign x_2215 = v_4230 | ~v_896;
assign x_2216 = v_4230 | ~v_855;
assign x_2217 = v_4230 | ~v_856;
assign x_2218 = v_4230 | ~v_897;
assign x_2219 = v_4230 | ~v_898;
assign x_2220 = v_4230 | ~v_899;
assign x_2221 = v_4230 | ~v_900;
assign x_2222 = v_4230 | ~v_182;
assign x_2223 = v_4230 | ~v_179;
assign x_2224 = v_4230 | ~v_163;
assign x_2225 = v_4230 | ~v_162;
assign x_2226 = v_4230 | ~v_161;
assign x_2227 = v_4230 | ~v_137;
assign x_2228 = v_4230 | ~v_136;
assign x_2229 = v_4230 | ~v_134;
assign x_2230 = v_4230 | ~v_18;
assign x_2231 = v_4230 | ~v_17;
assign x_2232 = v_4230 | ~v_16;
assign x_2233 = v_4230 | ~v_11;
assign x_2234 = ~v_4228 | ~v_4227 | ~v_4226 | v_4229;
assign x_2235 = v_4228 | ~v_3616;
assign x_2236 = v_4228 | ~v_3617;
assign x_2237 = v_4228 | ~v_3618;
assign x_2238 = v_4228 | ~v_3619;
assign x_2239 = v_4228 | ~v_2093;
assign x_2240 = v_4228 | ~v_2094;
assign x_2241 = v_4228 | ~v_2095;
assign x_2242 = v_4228 | ~v_2096;
assign x_2243 = v_4228 | ~v_3494;
assign x_2244 = v_4228 | ~v_3495;
assign x_2245 = v_4228 | ~v_2109;
assign x_2246 = v_4228 | ~v_2110;
assign x_2247 = v_4228 | ~v_2111;
assign x_2248 = v_4228 | ~v_2112;
assign x_2249 = v_4228 | ~v_3496;
assign x_2250 = v_4228 | ~v_3499;
assign x_2251 = v_4228 | ~v_2075;
assign x_2252 = v_4228 | ~v_4216;
assign x_2253 = v_4228 | ~v_4217;
assign x_2254 = v_4228 | ~v_2078;
assign x_2255 = v_4228 | ~v_4218;
assign x_2256 = v_4228 | ~v_4219;
assign x_2257 = v_4228 | ~v_973;
assign x_2258 = v_4228 | ~v_974;
assign x_2259 = v_4228 | ~v_885;
assign x_2260 = v_4228 | ~v_886;
assign x_2261 = v_4228 | ~v_975;
assign x_2262 = v_4228 | ~v_976;
assign x_2263 = v_4228 | ~v_977;
assign x_2264 = v_4228 | ~v_978;
assign x_2265 = v_4228 | ~v_3502;
assign x_2266 = v_4228 | ~v_3503;
assign x_2267 = v_4228 | ~v_184;
assign x_2268 = v_4228 | ~v_181;
assign x_2269 = v_4228 | ~v_172;
assign x_2270 = v_4228 | ~v_171;
assign x_2271 = v_4228 | ~v_170;
assign x_2272 = v_4228 | ~v_169;
assign x_2273 = v_4228 | ~v_150;
assign x_2274 = v_4228 | ~v_149;
assign x_2275 = v_4228 | ~v_148;
assign x_2276 = v_4228 | ~v_147;
assign x_2277 = v_4228 | ~v_102;
assign x_2278 = v_4228 | ~v_101;
assign x_2279 = v_4227 | ~v_3611;
assign x_2280 = v_4227 | ~v_3612;
assign x_2281 = v_4227 | ~v_3613;
assign x_2282 = v_4227 | ~v_3614;
assign x_2283 = v_4227 | ~v_2088;
assign x_2284 = v_4227 | ~v_2089;
assign x_2285 = v_4227 | ~v_2090;
assign x_2286 = v_4227 | ~v_2091;
assign x_2287 = v_4227 | ~v_3479;
assign x_2288 = v_4227 | ~v_3480;
assign x_2289 = v_4227 | ~v_2104;
assign x_2290 = v_4227 | ~v_2105;
assign x_2291 = v_4227 | ~v_2106;
assign x_2292 = v_4227 | ~v_2107;
assign x_2293 = v_4227 | ~v_3481;
assign x_2294 = v_4227 | ~v_3484;
assign x_2295 = v_4227 | ~v_2060;
assign x_2296 = v_4227 | ~v_4211;
assign x_2297 = v_4227 | ~v_4212;
assign x_2298 = v_4227 | ~v_2063;
assign x_2299 = v_4227 | ~v_4213;
assign x_2300 = v_4227 | ~v_4214;
assign x_2301 = v_4227 | ~v_958;
assign x_2302 = v_4227 | ~v_959;
assign x_2303 = v_4227 | ~v_870;
assign x_2304 = v_4227 | ~v_871;
assign x_2305 = v_4227 | ~v_960;
assign x_2306 = v_4227 | ~v_961;
assign x_2307 = v_4227 | ~v_962;
assign x_2308 = v_4227 | ~v_963;
assign x_2309 = v_4227 | ~v_3487;
assign x_2310 = v_4227 | ~v_3488;
assign x_2311 = v_4227 | ~v_183;
assign x_2312 = v_4227 | ~v_180;
assign x_2313 = v_4227 | ~v_168;
assign x_2314 = v_4227 | ~v_167;
assign x_2315 = v_4227 | ~v_166;
assign x_2316 = v_4227 | ~v_165;
assign x_2317 = v_4227 | ~v_145;
assign x_2318 = v_4227 | ~v_144;
assign x_2319 = v_4227 | ~v_143;
assign x_2320 = v_4227 | ~v_142;
assign x_2321 = v_4227 | ~v_60;
assign x_2322 = v_4227 | ~v_59;
assign x_2323 = v_4226 | ~v_3606;
assign x_2324 = v_4226 | ~v_3607;
assign x_2325 = v_4226 | ~v_3608;
assign x_2326 = v_4226 | ~v_3609;
assign x_2327 = v_4226 | ~v_2083;
assign x_2328 = v_4226 | ~v_2084;
assign x_2329 = v_4226 | ~v_2085;
assign x_2330 = v_4226 | ~v_2086;
assign x_2331 = v_4226 | ~v_3464;
assign x_2332 = v_4226 | ~v_3465;
assign x_2333 = v_4226 | ~v_2099;
assign x_2334 = v_4226 | ~v_2100;
assign x_2335 = v_4226 | ~v_2101;
assign x_2336 = v_4226 | ~v_2102;
assign x_2337 = v_4226 | ~v_3466;
assign x_2338 = v_4226 | ~v_3469;
assign x_2339 = v_4226 | ~v_2045;
assign x_2340 = v_4226 | ~v_4206;
assign x_2341 = v_4226 | ~v_4207;
assign x_2342 = v_4226 | ~v_2048;
assign x_2343 = v_4226 | ~v_4208;
assign x_2344 = v_4226 | ~v_4209;
assign x_2345 = v_4226 | ~v_943;
assign x_2346 = v_4226 | ~v_944;
assign x_2347 = v_4226 | ~v_855;
assign x_2348 = v_4226 | ~v_856;
assign x_2349 = v_4226 | ~v_945;
assign x_2350 = v_4226 | ~v_946;
assign x_2351 = v_4226 | ~v_947;
assign x_2352 = v_4226 | ~v_948;
assign x_2353 = v_4226 | ~v_3471;
assign x_2354 = v_4226 | ~v_3472;
assign x_2355 = v_4226 | ~v_182;
assign x_2356 = v_4226 | ~v_179;
assign x_2357 = v_4226 | ~v_164;
assign x_2358 = v_4226 | ~v_163;
assign x_2359 = v_4226 | ~v_162;
assign x_2360 = v_4226 | ~v_161;
assign x_2361 = v_4226 | ~v_137;
assign x_2362 = v_4226 | ~v_136;
assign x_2363 = v_4226 | ~v_135;
assign x_2364 = v_4226 | ~v_134;
assign x_2365 = v_4226 | ~v_17;
assign x_2366 = v_4226 | ~v_16;
assign x_2367 = ~v_4224 | ~v_4223 | ~v_4222 | v_4225;
assign x_2368 = v_4224 | ~v_3616;
assign x_2369 = v_4224 | ~v_3617;
assign x_2370 = v_4224 | ~v_3618;
assign x_2371 = v_4224 | ~v_3619;
assign x_2372 = v_4224 | ~v_2093;
assign x_2373 = v_4224 | ~v_2094;
assign x_2374 = v_4224 | ~v_2095;
assign x_2375 = v_4224 | ~v_2096;
assign x_2376 = v_4224 | ~v_3548;
assign x_2377 = v_4224 | ~v_3549;
assign x_2378 = v_4224 | ~v_3550;
assign x_2379 = v_4224 | ~v_3551;
assign x_2380 = v_4224 | ~v_2071;
assign x_2381 = v_4224 | ~v_2072;
assign x_2382 = v_4224 | ~v_2073;
assign x_2383 = v_4224 | ~v_2074;
assign x_2384 = v_4224 | ~v_3496;
assign x_2385 = v_4224 | ~v_3499;
assign x_2386 = v_4224 | ~v_2075;
assign x_2387 = v_4224 | ~v_4216;
assign x_2388 = v_4224 | ~v_4217;
assign x_2389 = v_4224 | ~v_2078;
assign x_2390 = v_4224 | ~v_4218;
assign x_2391 = v_4224 | ~v_4219;
assign x_2392 = v_4224 | ~v_881;
assign x_2393 = v_4224 | ~v_882;
assign x_2394 = v_4224 | ~v_883;
assign x_2395 = v_4224 | ~v_884;
assign x_2396 = v_4224 | ~v_885;
assign x_2397 = v_4224 | ~v_886;
assign x_2398 = v_4224 | ~v_837;
assign x_2399 = v_4224 | ~v_838;
assign x_2400 = v_4224 | ~v_184;
assign x_2401 = v_4224 | ~v_181;
assign x_2402 = v_4224 | ~v_171;
assign x_2403 = v_4224 | ~v_170;
assign x_2404 = v_4224 | ~v_169;
assign x_2405 = v_4224 | ~v_160;
assign x_2406 = v_4224 | ~v_150;
assign x_2407 = v_4224 | ~v_149;
assign x_2408 = v_4224 | ~v_148;
assign x_2409 = v_4224 | ~v_103;
assign x_2410 = v_4224 | ~v_102;
assign x_2411 = v_4224 | ~v_95;
assign x_2412 = v_4223 | ~v_3611;
assign x_2413 = v_4223 | ~v_3612;
assign x_2414 = v_4223 | ~v_3613;
assign x_2415 = v_4223 | ~v_3614;
assign x_2416 = v_4223 | ~v_2088;
assign x_2417 = v_4223 | ~v_2089;
assign x_2418 = v_4223 | ~v_2090;
assign x_2419 = v_4223 | ~v_2091;
assign x_2420 = v_4223 | ~v_3543;
assign x_2421 = v_4223 | ~v_3544;
assign x_2422 = v_4223 | ~v_3545;
assign x_2423 = v_4223 | ~v_3546;
assign x_2424 = v_4223 | ~v_2056;
assign x_2425 = v_4223 | ~v_2057;
assign x_2426 = v_4223 | ~v_2058;
assign x_2427 = v_4223 | ~v_2059;
assign x_2428 = v_4223 | ~v_3481;
assign x_2429 = v_4223 | ~v_3484;
assign x_2430 = v_4223 | ~v_2060;
assign x_2431 = v_4223 | ~v_4211;
assign x_2432 = v_4223 | ~v_4212;
assign x_2433 = v_4223 | ~v_2063;
assign x_2434 = v_4223 | ~v_4213;
assign x_2435 = v_4223 | ~v_4214;
assign x_2436 = v_4223 | ~v_866;
assign x_2437 = v_4223 | ~v_867;
assign x_2438 = v_4223 | ~v_868;
assign x_2439 = v_4223 | ~v_869;
assign x_2440 = v_4223 | ~v_870;
assign x_2441 = v_4223 | ~v_871;
assign x_2442 = v_4223 | ~v_804;
assign x_2443 = v_4223 | ~v_805;
assign x_2444 = v_4223 | ~v_183;
assign x_2445 = v_4223 | ~v_180;
assign x_2446 = v_4223 | ~v_167;
assign x_2447 = v_4223 | ~v_166;
assign x_2448 = v_4223 | ~v_165;
assign x_2449 = v_4223 | ~v_159;
assign x_2450 = v_4223 | ~v_145;
assign x_2451 = v_4223 | ~v_144;
assign x_2452 = v_4223 | ~v_143;
assign x_2453 = v_4223 | ~v_61;
assign x_2454 = v_4223 | ~v_60;
assign x_2455 = v_4223 | ~v_53;
assign x_2456 = v_4222 | ~v_3606;
assign x_2457 = v_4222 | ~v_3607;
assign x_2458 = v_4222 | ~v_3608;
assign x_2459 = v_4222 | ~v_3609;
assign x_2460 = v_4222 | ~v_2083;
assign x_2461 = v_4222 | ~v_2084;
assign x_2462 = v_4222 | ~v_2085;
assign x_2463 = v_4222 | ~v_2086;
assign x_2464 = v_4222 | ~v_3538;
assign x_2465 = v_4222 | ~v_3539;
assign x_2466 = v_4222 | ~v_3540;
assign x_2467 = v_4222 | ~v_3541;
assign x_2468 = v_4222 | ~v_2041;
assign x_2469 = v_4222 | ~v_2042;
assign x_2470 = v_4222 | ~v_2043;
assign x_2471 = v_4222 | ~v_2044;
assign x_2472 = v_4222 | ~v_3466;
assign x_2473 = v_4222 | ~v_3469;
assign x_2474 = v_4222 | ~v_2045;
assign x_2475 = v_4222 | ~v_4206;
assign x_2476 = v_4222 | ~v_4207;
assign x_2477 = v_4222 | ~v_2048;
assign x_2478 = v_4222 | ~v_4208;
assign x_2479 = v_4222 | ~v_4209;
assign x_2480 = v_4222 | ~v_851;
assign x_2481 = v_4222 | ~v_852;
assign x_2482 = v_4222 | ~v_853;
assign x_2483 = v_4222 | ~v_854;
assign x_2484 = v_4222 | ~v_855;
assign x_2485 = v_4222 | ~v_856;
assign x_2486 = v_4222 | ~v_771;
assign x_2487 = v_4222 | ~v_772;
assign x_2488 = v_4222 | ~v_182;
assign x_2489 = v_4222 | ~v_179;
assign x_2490 = v_4222 | ~v_163;
assign x_2491 = v_4222 | ~v_162;
assign x_2492 = v_4222 | ~v_161;
assign x_2493 = v_4222 | ~v_155;
assign x_2494 = v_4222 | ~v_137;
assign x_2495 = v_4222 | ~v_136;
assign x_2496 = v_4222 | ~v_135;
assign x_2497 = v_4222 | ~v_18;
assign x_2498 = v_4222 | ~v_17;
assign x_2499 = v_4222 | ~v_10;
assign x_2500 = ~v_4220 | ~v_4215 | ~v_4210 | v_4221;
assign x_2501 = v_4220 | ~v_3548;
assign x_2502 = v_4220 | ~v_3549;
assign x_2503 = v_4220 | ~v_3550;
assign x_2504 = v_4220 | ~v_3551;
assign x_2505 = v_4220 | ~v_2071;
assign x_2506 = v_4220 | ~v_2072;
assign x_2507 = v_4220 | ~v_2073;
assign x_2508 = v_4220 | ~v_2074;
assign x_2509 = v_4220 | ~v_3496;
assign x_2510 = v_4220 | ~v_3497;
assign x_2511 = v_4220 | ~v_3498;
assign x_2512 = v_4220 | ~v_3499;
assign x_2513 = v_4220 | ~v_3500;
assign x_2514 = v_4220 | ~v_3501;
assign x_2515 = v_4220 | ~v_2075;
assign x_2516 = v_4220 | ~v_4216;
assign x_2517 = v_4220 | ~v_2076;
assign x_2518 = v_4220 | ~v_4217;
assign x_2519 = v_4220 | ~v_2077;
assign x_2520 = v_4220 | ~v_2078;
assign x_2521 = v_4220 | ~v_4218;
assign x_2522 = v_4220 | ~v_2079;
assign x_2523 = v_4220 | ~v_4219;
assign x_2524 = v_4220 | ~v_2080;
assign x_2525 = v_4220 | ~v_833;
assign x_2526 = v_4220 | ~v_834;
assign x_2527 = v_4220 | ~v_835;
assign x_2528 = v_4220 | ~v_836;
assign x_2529 = v_4220 | ~v_837;
assign x_2530 = v_4220 | ~v_838;
assign x_2531 = v_4220 | ~v_839;
assign x_2532 = v_4220 | ~v_840;
assign x_2533 = v_4220 | ~v_184;
assign x_2534 = v_4220 | ~v_169;
assign x_2535 = v_4220 | ~v_160;
assign x_2536 = v_4220 | ~v_150;
assign x_2537 = v_4220 | ~v_149;
assign x_2538 = v_4220 | ~v_148;
assign x_2539 = v_4220 | ~v_147;
assign x_2540 = v_4220 | ~v_103;
assign x_2541 = v_4220 | ~v_102;
assign x_2542 = v_4220 | ~v_100;
assign x_2543 = v_4220 | ~v_98;
assign x_2544 = v_4220 | ~v_94;
assign x_2545 = ~v_123 | ~v_139 | v_4219;
assign x_2546 = ~v_120 | ~v_140 | v_4218;
assign x_2547 = ~v_108 | v_139 | v_4217;
assign x_2548 = ~v_105 | v_140 | v_4216;
assign x_2549 = v_4215 | ~v_3543;
assign x_2550 = v_4215 | ~v_3544;
assign x_2551 = v_4215 | ~v_3545;
assign x_2552 = v_4215 | ~v_3546;
assign x_2553 = v_4215 | ~v_2056;
assign x_2554 = v_4215 | ~v_2057;
assign x_2555 = v_4215 | ~v_2058;
assign x_2556 = v_4215 | ~v_2059;
assign x_2557 = v_4215 | ~v_3481;
assign x_2558 = v_4215 | ~v_3482;
assign x_2559 = v_4215 | ~v_3483;
assign x_2560 = v_4215 | ~v_3484;
assign x_2561 = v_4215 | ~v_3485;
assign x_2562 = v_4215 | ~v_2060;
assign x_2563 = v_4215 | ~v_4211;
assign x_2564 = v_4215 | ~v_2061;
assign x_2565 = v_4215 | ~v_4212;
assign x_2566 = v_4215 | ~v_2062;
assign x_2567 = v_4215 | ~v_2063;
assign x_2568 = v_4215 | ~v_4213;
assign x_2569 = v_4215 | ~v_2064;
assign x_2570 = v_4215 | ~v_4214;
assign x_2571 = v_4215 | ~v_2065;
assign x_2572 = v_4215 | ~v_800;
assign x_2573 = v_4215 | ~v_801;
assign x_2574 = v_4215 | ~v_802;
assign x_2575 = v_4215 | ~v_803;
assign x_2576 = v_4215 | ~v_804;
assign x_2577 = v_4215 | ~v_805;
assign x_2578 = v_4215 | ~v_806;
assign x_2579 = v_4215 | ~v_807;
assign x_2580 = v_4215 | ~v_3486;
assign x_2581 = v_4215 | ~v_183;
assign x_2582 = v_4215 | ~v_165;
assign x_2583 = v_4215 | ~v_159;
assign x_2584 = v_4215 | ~v_145;
assign x_2585 = v_4215 | ~v_144;
assign x_2586 = v_4215 | ~v_143;
assign x_2587 = v_4215 | ~v_142;
assign x_2588 = v_4215 | ~v_61;
assign x_2589 = v_4215 | ~v_60;
assign x_2590 = v_4215 | ~v_58;
assign x_2591 = v_4215 | ~v_56;
assign x_2592 = v_4215 | ~v_52;
assign x_2593 = ~v_81 | ~v_139 | v_4214;
assign x_2594 = ~v_78 | ~v_140 | v_4213;
assign x_2595 = ~v_66 | v_139 | v_4212;
assign x_2596 = ~v_63 | v_140 | v_4211;
assign x_2597 = v_4210 | ~v_3538;
assign x_2598 = v_4210 | ~v_3539;
assign x_2599 = v_4210 | ~v_3540;
assign x_2600 = v_4210 | ~v_3541;
assign x_2601 = v_4210 | ~v_2041;
assign x_2602 = v_4210 | ~v_2042;
assign x_2603 = v_4210 | ~v_2043;
assign x_2604 = v_4210 | ~v_2044;
assign x_2605 = v_4210 | ~v_3466;
assign x_2606 = v_4210 | ~v_3467;
assign x_2607 = v_4210 | ~v_3468;
assign x_2608 = v_4210 | ~v_3469;
assign x_2609 = v_4210 | ~v_3470;
assign x_2610 = v_4210 | ~v_2045;
assign x_2611 = v_4210 | ~v_4206;
assign x_2612 = v_4210 | ~v_2046;
assign x_2613 = v_4210 | ~v_4207;
assign x_2614 = v_4210 | ~v_2047;
assign x_2615 = v_4210 | ~v_2048;
assign x_2616 = v_4210 | ~v_4208;
assign x_2617 = v_4210 | ~v_2049;
assign x_2618 = v_4210 | ~v_4209;
assign x_2619 = v_4210 | ~v_2050;
assign x_2620 = v_4210 | ~v_767;
assign x_2621 = v_4210 | ~v_768;
assign x_2622 = v_4210 | ~v_769;
assign x_2623 = v_4210 | ~v_770;
assign x_2624 = v_4210 | ~v_771;
assign x_2625 = v_4210 | ~v_772;
assign x_2626 = v_4210 | ~v_773;
assign x_2627 = v_4210 | ~v_774;
assign x_2628 = v_4210 | ~v_182;
assign x_2629 = v_4210 | ~v_161;
assign x_2630 = v_4210 | ~v_155;
assign x_2631 = v_4210 | ~v_137;
assign x_2632 = v_4210 | ~v_3473;
assign x_2633 = v_4210 | ~v_136;
assign x_2634 = v_4210 | ~v_135;
assign x_2635 = v_4210 | ~v_134;
assign x_2636 = v_4210 | ~v_18;
assign x_2637 = v_4210 | ~v_17;
assign x_2638 = v_4210 | ~v_15;
assign x_2639 = v_4210 | ~v_13;
assign x_2640 = v_4210 | ~v_9;
assign x_2641 = ~v_39 | ~v_139 | v_4209;
assign x_2642 = ~v_36 | ~v_140 | v_4208;
assign x_2643 = ~v_24 | v_139 | v_4207;
assign x_2644 = ~v_21 | v_140 | v_4206;
assign x_2645 = v_4205 | ~v_1566;
assign x_2646 = v_4205 | ~v_731;
assign x_2647 = v_4204 | ~v_739;
assign x_2648 = v_4204 | ~v_735;
assign x_2649 = ~v_725 | ~v_724 | ~v_723 | ~v_722 | ~v_4202 | ~v_4198 | ~v_4194 | ~v_4190 | ~v_4186 | ~v_4182 | ~v_4178 | ~v_4174 | ~v_4170 | ~v_4166 | ~v_4162 | ~v_4158 | ~v_4154 | ~v_4150 | ~v_4146 | ~v_4142 | ~v_4126 | v_4203;
assign x_2650 = v_4202 | ~v_4199;
assign x_2651 = v_4202 | ~v_4200;
assign x_2652 = v_4202 | ~v_4201;
assign x_2653 = v_98 | v_103 | v_101 | v_97 | v_100 | v_95 | v_94 | v_99 | v_102 | ~v_719 | ~v_718 | v_169 | v_148 | v_184 | ~v_483 | ~v_717 | ~v_299 | ~v_482 | ~v_716 | ~v_298 | ~v_1962 | ~v_1898 | ~v_4140 | ~v_1961 | ~v_1897 | ~v_4139 | ~v_1896 | ~v_1960 | ~v_1895 | ~v_4138 | ~v_1959 | ~v_1894 | ~v_4137 | ~v_1893 | ~v_3386 | ~v_3320 | ~v_3385 | ~v_3319 | ~v_3318 | ~v_3384 | ~v_3317 | ~v_3383 | ~v_3316 | ~v_3315 | v_4201;
assign x_2654 = v_53 | v_56 | v_55 | v_61 | v_52 | v_60 | v_59 | v_58 | v_57 | ~v_714 | ~v_713 | v_143 | v_165 | v_183 | ~v_3381 | ~v_3305 | ~v_266 | ~v_3380 | ~v_468 | ~v_712 | ~v_467 | ~v_711 | ~v_265 | ~v_1957 | ~v_1883 | ~v_4135 | ~v_1956 | ~v_1882 | ~v_4134 | ~v_1881 | ~v_1955 | ~v_1880 | ~v_4133 | ~v_1954 | ~v_1879 | ~v_4132 | ~v_1878 | ~v_3304 | ~v_3303 | ~v_3379 | ~v_3302 | ~v_3378 | ~v_3301 | ~v_3300 | v_4200;
assign x_2655 = v_13 | v_9 | v_18 | v_17 | v_16 | v_15 | v_14 | v_12 | v_10 | ~v_453 | ~v_709 | ~v_452 | ~v_708 | v_135 | ~v_707 | ~v_706 | ~v_3292 | v_161 | v_182 | ~v_233 | ~v_232 | ~v_1952 | ~v_1868 | ~v_4130 | ~v_1951 | ~v_1867 | ~v_4129 | ~v_1866 | ~v_1950 | ~v_1865 | ~v_4128 | ~v_1949 | ~v_1864 | ~v_4127 | ~v_1863 | ~v_3376 | ~v_3289 | ~v_3375 | ~v_3288 | ~v_3374 | ~v_3287 | ~v_3373 | ~v_3286 | ~v_3285 | v_4199;
assign x_2656 = v_4198 | ~v_4195;
assign x_2657 = v_4198 | ~v_4196;
assign x_2658 = v_4198 | ~v_4197;
assign x_2659 = v_101 | v_97 | v_100 | v_99 | v_93 | v_102 | v_172 | v_171 | v_170 | v_148 | v_147 | v_184 | ~v_483 | ~v_482 | ~v_593 | ~v_592 | ~v_545 | ~v_591 | ~v_590 | ~v_544 | ~v_1962 | ~v_4140 | ~v_1961 | ~v_4139 | ~v_1896 | ~v_1960 | ~v_4138 | ~v_1959 | ~v_4137 | ~v_1893 | ~v_3386 | ~v_3385 | ~v_3318 | ~v_3384 | ~v_3383 | ~v_3315 | ~v_2014 | ~v_2013 | ~v_2012 | ~v_2011 | ~v_3406 | ~v_3405 | ~v_3404 | ~v_3403 | v_4197;
assign x_2660 = v_55 | v_51 | v_60 | v_59 | v_58 | v_57 | v_143 | v_142 | v_168 | v_167 | v_166 | v_183 | ~v_3381 | ~v_3380 | ~v_468 | ~v_467 | ~v_588 | ~v_587 | ~v_530 | ~v_586 | ~v_585 | ~v_529 | ~v_1957 | ~v_4135 | ~v_1956 | ~v_4134 | ~v_1881 | ~v_1955 | ~v_4133 | ~v_1954 | ~v_4132 | ~v_1878 | ~v_3303 | ~v_3379 | ~v_3378 | ~v_3300 | ~v_2009 | ~v_2008 | ~v_2007 | ~v_2006 | ~v_3401 | ~v_3400 | ~v_3399 | ~v_3398 | v_4196;
assign x_2661 = v_17 | v_16 | v_8 | v_15 | v_14 | v_12 | ~v_453 | ~v_452 | v_135 | v_134 | v_164 | v_163 | v_162 | v_182 | ~v_583 | ~v_582 | ~v_515 | ~v_581 | ~v_580 | ~v_514 | ~v_1952 | ~v_4130 | ~v_1951 | ~v_4129 | ~v_1866 | ~v_1950 | ~v_4128 | ~v_1949 | ~v_4127 | ~v_1863 | ~v_3376 | ~v_3375 | ~v_3288 | ~v_3374 | ~v_3373 | ~v_3285 | ~v_2004 | ~v_2003 | ~v_2002 | ~v_2001 | ~v_3396 | ~v_3395 | ~v_3394 | ~v_3393 | v_4195;
assign x_2662 = v_4194 | ~v_4191;
assign x_2663 = v_4194 | ~v_4192;
assign x_2664 = v_4194 | ~v_4193;
assign x_2665 = v_103 | v_101 | v_96 | v_100 | v_95 | v_93 | v_102 | v_171 | v_170 | v_150 | v_149 | v_184 | ~v_545 | ~v_544 | ~v_561 | ~v_560 | ~v_559 | ~v_558 | ~v_387 | ~v_386 | ~v_4140 | ~v_4139 | ~v_1896 | ~v_4138 | ~v_4137 | ~v_1893 | ~v_3318 | ~v_3315 | ~v_2014 | ~v_2013 | ~v_2012 | ~v_2011 | ~v_3406 | ~v_3405 | ~v_3404 | ~v_3403 | ~v_1946 | ~v_1945 | ~v_1944 | ~v_1943 | ~v_3354 | ~v_3353 | ~v_3352 | ~v_3351 | v_4193;
assign x_2666 = v_54 | v_53 | v_61 | v_51 | v_60 | v_59 | v_58 | v_144 | v_145 | v_167 | v_166 | v_183 | ~v_530 | ~v_529 | ~v_556 | ~v_555 | ~v_554 | ~v_553 | ~v_372 | ~v_371 | ~v_4135 | ~v_4134 | ~v_1881 | ~v_4133 | ~v_4132 | ~v_1878 | ~v_3303 | ~v_3300 | ~v_2009 | ~v_2008 | ~v_2007 | ~v_2006 | ~v_3401 | ~v_3400 | ~v_3399 | ~v_3398 | ~v_1941 | ~v_1940 | ~v_1939 | ~v_1938 | ~v_3349 | ~v_3348 | ~v_3347 | ~v_3346 | v_4192;
assign x_2667 = v_18 | v_17 | v_16 | v_8 | v_15 | v_11 | v_10 | v_136 | v_137 | v_163 | v_162 | v_182 | ~v_515 | ~v_514 | ~v_551 | ~v_550 | ~v_549 | ~v_548 | ~v_357 | ~v_356 | ~v_4130 | ~v_4129 | ~v_1866 | ~v_4128 | ~v_4127 | ~v_1863 | ~v_3288 | ~v_3285 | ~v_2004 | ~v_2003 | ~v_2002 | ~v_2001 | ~v_3396 | ~v_3395 | ~v_3394 | ~v_3393 | ~v_1936 | ~v_1935 | ~v_1934 | ~v_1933 | ~v_3344 | ~v_3343 | ~v_3342 | ~v_3341 | v_4191;
assign x_2668 = v_4190 | ~v_4187;
assign x_2669 = v_4190 | ~v_4188;
assign x_2670 = v_4190 | ~v_4189;
assign x_2671 = v_103 | v_101 | v_100 | v_93 | v_151 | v_171 | v_170 | v_150 | v_149 | v_148 | v_147 | v_184 | ~v_3322 | ~v_3321 | ~v_577 | ~v_576 | ~v_545 | ~v_544 | ~v_575 | ~v_574 | ~v_435 | ~v_434 | ~v_4140 | ~v_4139 | ~v_1896 | ~v_4138 | ~v_4137 | ~v_1893 | ~v_3318 | ~v_3315 | ~v_2014 | ~v_2013 | ~v_2012 | ~v_2011 | ~v_3406 | ~v_3405 | ~v_3404 | ~v_3403 | ~v_1930 | ~v_1929 | ~v_1928 | ~v_1927 | ~v_3314 | ~v_3313 | v_4189;
assign x_2672 = v_61 | v_51 | v_59 | v_58 | v_144 | v_145 | v_143 | v_142 | v_167 | v_166 | v_146 | v_183 | ~v_3307 | ~v_3306 | ~v_572 | ~v_571 | ~v_530 | ~v_529 | ~v_570 | ~v_569 | ~v_420 | ~v_419 | ~v_4135 | ~v_4134 | ~v_1881 | ~v_4133 | ~v_4132 | ~v_1878 | ~v_3303 | ~v_3300 | ~v_2009 | ~v_2008 | ~v_2007 | ~v_2006 | ~v_3401 | ~v_3400 | ~v_3399 | ~v_3398 | ~v_1925 | ~v_1924 | ~v_1923 | ~v_1922 | ~v_3299 | ~v_3298 | v_4188;
assign x_2673 = v_18 | v_16 | v_8 | v_15 | v_136 | v_135 | v_134 | v_137 | v_138 | v_163 | v_162 | v_182 | ~v_3291 | ~v_3290 | ~v_567 | ~v_566 | ~v_515 | ~v_514 | ~v_565 | ~v_564 | ~v_405 | ~v_404 | ~v_4130 | ~v_4129 | ~v_1866 | ~v_4128 | ~v_4127 | ~v_1863 | ~v_3288 | ~v_3285 | ~v_2004 | ~v_2003 | ~v_2002 | ~v_2001 | ~v_3396 | ~v_3395 | ~v_3394 | ~v_3393 | ~v_1920 | ~v_1919 | ~v_1918 | ~v_1917 | ~v_3284 | ~v_3283 | v_4187;
assign x_2674 = v_4186 | ~v_4183;
assign x_2675 = v_4186 | ~v_4184;
assign x_2676 = v_4186 | ~v_4185;
assign x_2677 = v_103 | v_100 | v_93 | v_102 | v_171 | v_170 | v_160 | v_150 | v_149 | v_148 | v_147 | v_184 | ~v_545 | ~v_544 | ~v_543 | ~v_542 | ~v_541 | ~v_540 | ~v_297 | ~v_296 | ~v_4140 | ~v_4139 | ~v_1896 | ~v_4138 | ~v_4137 | ~v_1893 | ~v_3318 | ~v_3315 | ~v_2014 | ~v_2013 | ~v_2012 | ~v_2011 | ~v_3406 | ~v_3405 | ~v_3404 | ~v_3403 | ~v_1892 | ~v_1891 | ~v_1890 | ~v_1889 | ~v_3370 | ~v_3369 | ~v_3368 | ~v_3367 | v_4185;
assign x_2678 = v_61 | v_51 | v_60 | v_58 | v_144 | v_159 | v_145 | v_143 | v_142 | v_167 | v_166 | v_183 | ~v_530 | ~v_529 | ~v_528 | ~v_527 | ~v_526 | ~v_525 | ~v_264 | ~v_263 | ~v_4135 | ~v_4134 | ~v_1881 | ~v_4133 | ~v_4132 | ~v_1878 | ~v_3303 | ~v_3300 | ~v_2009 | ~v_2008 | ~v_2007 | ~v_2006 | ~v_3401 | ~v_3400 | ~v_3399 | ~v_3398 | ~v_1877 | ~v_1876 | ~v_1875 | ~v_1874 | ~v_3365 | ~v_3364 | ~v_3363 | ~v_3362 | v_4184;
assign x_2679 = v_18 | v_17 | v_8 | v_15 | v_136 | v_135 | v_134 | v_137 | v_163 | v_162 | v_155 | v_182 | ~v_515 | ~v_514 | ~v_513 | ~v_512 | ~v_511 | ~v_510 | ~v_231 | ~v_230 | ~v_4130 | ~v_4129 | ~v_1866 | ~v_4128 | ~v_4127 | ~v_1863 | ~v_3288 | ~v_3285 | ~v_2004 | ~v_2003 | ~v_2002 | ~v_2001 | ~v_3396 | ~v_3395 | ~v_3394 | ~v_3393 | ~v_1862 | ~v_1861 | ~v_1860 | ~v_1859 | ~v_3360 | ~v_3359 | ~v_3358 | ~v_3357 | v_4183;
assign x_2680 = v_4182 | ~v_4179;
assign x_2681 = v_4182 | ~v_4180;
assign x_2682 = v_4182 | ~v_4181;
assign x_2683 = v_98 | v_103 | v_101 | v_96 | v_100 | v_94 | v_151 | v_169 | v_150 | v_149 | v_147 | v_184 | ~v_299 | ~v_298 | ~v_387 | ~v_386 | ~v_499 | ~v_498 | ~v_497 | ~v_496 | ~v_1898 | ~v_4140 | ~v_1897 | ~v_4139 | ~v_1896 | ~v_1895 | ~v_4138 | ~v_1894 | ~v_4137 | ~v_1893 | ~v_3320 | ~v_3319 | ~v_3318 | ~v_3317 | ~v_3316 | ~v_3315 | ~v_1946 | ~v_1945 | ~v_1944 | ~v_1943 | ~v_3354 | ~v_3353 | ~v_3352 | ~v_3351 | v_4181;
assign x_2684 = v_54 | v_56 | v_61 | v_52 | v_59 | v_58 | v_144 | v_145 | v_142 | v_165 | v_146 | v_183 | ~v_3305 | ~v_266 | ~v_265 | ~v_372 | ~v_371 | ~v_494 | ~v_493 | ~v_492 | ~v_491 | ~v_1883 | ~v_4135 | ~v_1882 | ~v_4134 | ~v_1881 | ~v_1880 | ~v_4133 | ~v_1879 | ~v_4132 | ~v_1878 | ~v_3304 | ~v_3303 | ~v_3302 | ~v_3301 | ~v_3300 | ~v_1941 | ~v_1940 | ~v_1939 | ~v_1938 | ~v_3349 | ~v_3348 | ~v_3347 | ~v_3346 | v_4180;
assign x_2685 = v_13 | v_9 | v_18 | v_16 | v_15 | v_11 | v_136 | v_134 | ~v_3292 | v_137 | v_138 | v_161 | v_182 | ~v_233 | ~v_232 | ~v_357 | ~v_356 | ~v_489 | ~v_488 | ~v_487 | ~v_486 | ~v_1868 | ~v_4130 | ~v_1867 | ~v_4129 | ~v_1866 | ~v_1865 | ~v_4128 | ~v_1864 | ~v_4127 | ~v_1863 | ~v_3289 | ~v_3288 | ~v_3287 | ~v_3286 | ~v_3285 | ~v_1936 | ~v_1935 | ~v_1934 | ~v_1933 | ~v_3344 | ~v_3343 | ~v_3342 | ~v_3341 | v_4179;
assign x_2686 = v_4178 | ~v_4175;
assign x_2687 = v_4178 | ~v_4176;
assign x_2688 = v_4178 | ~v_4177;
assign x_2689 = v_103 | v_101 | v_97 | v_100 | v_99 | v_102 | v_171 | v_170 | v_169 | v_148 | v_147 | v_184 | ~v_703 | ~v_702 | ~v_483 | ~v_482 | ~v_701 | ~v_653 | ~v_700 | ~v_652 | ~v_1962 | ~v_4140 | ~v_1961 | ~v_4139 | ~v_1896 | ~v_1960 | ~v_4138 | ~v_1959 | ~v_4137 | ~v_1893 | ~v_3386 | ~v_3385 | ~v_3318 | ~v_3384 | ~v_3383 | ~v_3315 | ~v_1982 | ~v_1981 | ~v_1980 | ~v_1979 | ~v_3338 | ~v_3337 | ~v_3336 | ~v_3335 | v_4177;
assign x_2690 = v_55 | v_61 | v_60 | v_59 | v_58 | v_57 | v_143 | v_142 | v_167 | v_166 | v_165 | v_183 | ~v_698 | ~v_697 | ~v_3381 | ~v_3380 | ~v_468 | ~v_467 | ~v_696 | ~v_638 | ~v_695 | ~v_637 | ~v_1957 | ~v_4135 | ~v_1956 | ~v_4134 | ~v_1881 | ~v_1955 | ~v_4133 | ~v_1954 | ~v_4132 | ~v_1878 | ~v_3303 | ~v_3379 | ~v_3378 | ~v_3300 | ~v_1977 | ~v_1976 | ~v_1975 | ~v_1974 | ~v_3333 | ~v_3332 | ~v_3331 | ~v_3330 | v_4176;
assign x_2691 = v_18 | v_17 | v_16 | v_15 | v_14 | v_12 | ~v_453 | ~v_452 | v_135 | v_134 | v_163 | v_162 | v_161 | v_182 | ~v_693 | ~v_692 | ~v_691 | ~v_623 | ~v_690 | ~v_622 | ~v_1952 | ~v_4130 | ~v_1951 | ~v_4129 | ~v_1866 | ~v_1950 | ~v_4128 | ~v_1949 | ~v_4127 | ~v_1863 | ~v_3376 | ~v_3375 | ~v_3288 | ~v_3374 | ~v_3373 | ~v_3285 | ~v_1972 | ~v_1971 | ~v_1970 | ~v_1969 | ~v_3328 | ~v_3327 | ~v_3326 | ~v_3325 | v_4175;
assign x_2692 = v_4174 | ~v_4171;
assign x_2693 = v_4174 | ~v_4172;
assign x_2694 = v_4174 | ~v_4173;
assign x_2695 = v_101 | v_96 | v_100 | v_102 | v_172 | v_171 | v_170 | v_169 | v_150 | v_149 | v_147 | v_184 | ~v_671 | ~v_670 | ~v_387 | ~v_386 | ~v_653 | ~v_652 | ~v_669 | ~v_668 | ~v_4140 | ~v_4139 | ~v_1896 | ~v_4138 | ~v_4137 | ~v_1893 | ~v_3318 | ~v_3315 | ~v_1946 | ~v_1945 | ~v_1944 | ~v_1943 | ~v_3354 | ~v_3353 | ~v_3352 | ~v_3351 | ~v_1982 | ~v_1981 | ~v_1980 | ~v_1979 | ~v_3338 | ~v_3337 | ~v_3336 | ~v_3335 | v_4173;
assign x_2696 = v_54 | v_60 | v_59 | v_58 | v_144 | v_145 | v_142 | v_168 | v_167 | v_166 | v_165 | v_183 | ~v_666 | ~v_665 | ~v_372 | ~v_371 | ~v_638 | ~v_637 | ~v_664 | ~v_663 | ~v_4135 | ~v_4134 | ~v_1881 | ~v_4133 | ~v_4132 | ~v_1878 | ~v_3303 | ~v_3300 | ~v_1941 | ~v_1940 | ~v_1939 | ~v_1938 | ~v_3349 | ~v_3348 | ~v_3347 | ~v_3346 | ~v_1977 | ~v_1976 | ~v_1975 | ~v_1974 | ~v_3333 | ~v_3332 | ~v_3331 | ~v_3330 | v_4172;
assign x_2697 = v_17 | v_16 | v_15 | v_11 | v_136 | v_134 | v_137 | v_164 | v_163 | v_162 | v_161 | v_182 | ~v_661 | ~v_660 | ~v_357 | ~v_356 | ~v_623 | ~v_622 | ~v_659 | ~v_658 | ~v_4130 | ~v_4129 | ~v_1866 | ~v_4128 | ~v_4127 | ~v_1863 | ~v_3288 | ~v_3285 | ~v_1936 | ~v_1935 | ~v_1934 | ~v_1933 | ~v_3344 | ~v_3343 | ~v_3342 | ~v_3341 | ~v_1972 | ~v_1971 | ~v_1970 | ~v_1969 | ~v_3328 | ~v_3327 | ~v_3326 | ~v_3325 | v_4171;
assign x_2698 = v_4170 | ~v_4167;
assign x_2699 = v_4170 | ~v_4168;
assign x_2700 = v_4170 | ~v_4169;
assign x_2701 = v_103 | v_101 | v_100 | v_95 | v_102 | v_171 | v_170 | v_169 | v_150 | v_149 | v_148 | v_184 | ~v_3322 | ~v_3321 | ~v_435 | ~v_434 | ~v_653 | ~v_652 | ~v_687 | ~v_686 | ~v_685 | ~v_684 | ~v_4140 | ~v_4139 | ~v_1896 | ~v_4138 | ~v_4137 | ~v_1893 | ~v_3318 | ~v_3315 | ~v_1930 | ~v_1929 | ~v_1928 | ~v_1927 | ~v_3314 | ~v_3313 | ~v_1982 | ~v_1981 | ~v_1980 | ~v_1979 | ~v_3338 | ~v_3337 | ~v_3336 | ~v_3335 | v_4169;
assign x_2702 = v_53 | v_61 | v_60 | v_59 | v_58 | v_144 | v_145 | v_143 | v_167 | v_166 | v_165 | v_183 | ~v_3307 | ~v_3306 | ~v_420 | ~v_419 | ~v_638 | ~v_637 | ~v_682 | ~v_681 | ~v_680 | ~v_679 | ~v_4135 | ~v_4134 | ~v_1881 | ~v_4133 | ~v_4132 | ~v_1878 | ~v_3303 | ~v_3300 | ~v_1925 | ~v_1924 | ~v_1923 | ~v_1922 | ~v_3299 | ~v_3298 | ~v_1977 | ~v_1976 | ~v_1975 | ~v_1974 | ~v_3333 | ~v_3332 | ~v_3331 | ~v_3330 | v_4168;
assign x_2703 = v_18 | v_17 | v_16 | v_15 | v_10 | v_136 | v_135 | v_137 | v_163 | v_162 | v_161 | v_182 | ~v_3291 | ~v_3290 | ~v_405 | ~v_404 | ~v_623 | ~v_622 | ~v_677 | ~v_676 | ~v_675 | ~v_674 | ~v_4130 | ~v_4129 | ~v_1866 | ~v_4128 | ~v_4127 | ~v_1863 | ~v_3288 | ~v_3285 | ~v_1920 | ~v_1919 | ~v_1918 | ~v_1917 | ~v_3284 | ~v_3283 | ~v_1972 | ~v_1971 | ~v_1970 | ~v_1969 | ~v_3328 | ~v_3327 | ~v_3326 | ~v_3325 | v_4167;
assign x_2704 = v_4166 | ~v_4163;
assign x_2705 = v_4166 | ~v_4164;
assign x_2706 = v_4166 | ~v_4165;
assign x_2707 = v_103 | v_100 | v_151 | v_171 | v_170 | v_169 | v_160 | v_150 | v_149 | v_148 | v_147 | v_184 | ~v_655 | ~v_654 | ~v_297 | ~v_296 | ~v_653 | ~v_652 | ~v_651 | ~v_650 | ~v_4140 | ~v_4139 | ~v_1896 | ~v_4138 | ~v_4137 | ~v_1893 | ~v_3318 | ~v_3315 | ~v_1892 | ~v_1891 | ~v_1890 | ~v_1889 | ~v_3370 | ~v_3369 | ~v_3368 | ~v_3367 | ~v_1982 | ~v_1981 | ~v_1980 | ~v_1979 | ~v_3338 | ~v_3337 | ~v_3336 | ~v_3335 | v_4165;
assign x_2708 = v_61 | v_58 | v_144 | v_159 | v_145 | v_143 | v_142 | v_167 | v_166 | v_165 | v_146 | v_183 | ~v_640 | ~v_639 | ~v_264 | ~v_263 | ~v_638 | ~v_637 | ~v_636 | ~v_635 | ~v_4135 | ~v_4134 | ~v_1881 | ~v_4133 | ~v_4132 | ~v_1878 | ~v_3303 | ~v_3300 | ~v_1877 | ~v_1876 | ~v_1875 | ~v_1874 | ~v_3365 | ~v_3364 | ~v_3363 | ~v_3362 | ~v_1977 | ~v_1976 | ~v_1975 | ~v_1974 | ~v_3333 | ~v_3332 | ~v_3331 | ~v_3330 | v_4164;
assign x_2709 = v_18 | v_15 | v_136 | v_135 | v_134 | v_137 | v_138 | v_163 | v_162 | v_161 | v_155 | v_182 | ~v_625 | ~v_624 | ~v_231 | ~v_230 | ~v_623 | ~v_622 | ~v_621 | ~v_620 | ~v_4130 | ~v_4129 | ~v_1866 | ~v_4128 | ~v_4127 | ~v_1863 | ~v_3288 | ~v_3285 | ~v_1862 | ~v_1861 | ~v_1860 | ~v_1859 | ~v_3360 | ~v_3359 | ~v_3358 | ~v_3357 | ~v_1972 | ~v_1971 | ~v_1970 | ~v_1969 | ~v_3328 | ~v_3327 | ~v_3326 | ~v_3325 | v_4163;
assign x_2710 = v_4162 | ~v_4159;
assign x_2711 = v_4162 | ~v_4160;
assign x_2712 = v_4162 | ~v_4161;
assign x_2713 = v_98 | v_103 | v_101 | v_100 | v_94 | v_102 | v_169 | v_150 | v_149 | v_148 | v_147 | v_184 | ~v_609 | ~v_608 | ~v_3322 | ~v_3321 | ~v_299 | ~v_298 | ~v_435 | ~v_434 | ~v_607 | ~v_606 | ~v_1898 | ~v_4140 | ~v_1897 | ~v_4139 | ~v_1896 | ~v_1895 | ~v_4138 | ~v_1894 | ~v_4137 | ~v_1893 | ~v_3320 | ~v_3319 | ~v_3318 | ~v_3317 | ~v_3316 | ~v_3315 | ~v_1930 | ~v_1929 | ~v_1928 | ~v_1927 | ~v_3314 | ~v_3313 | v_4161;
assign x_2714 = v_56 | v_61 | v_52 | v_60 | v_59 | v_58 | v_144 | v_145 | v_143 | v_142 | v_165 | v_183 | ~v_604 | ~v_603 | ~v_3307 | ~v_3306 | ~v_3305 | ~v_266 | ~v_265 | ~v_420 | ~v_419 | ~v_602 | ~v_601 | ~v_1883 | ~v_4135 | ~v_1882 | ~v_4134 | ~v_1881 | ~v_1880 | ~v_4133 | ~v_1879 | ~v_4132 | ~v_1878 | ~v_3304 | ~v_3303 | ~v_3302 | ~v_3301 | ~v_3300 | ~v_1925 | ~v_1924 | ~v_1923 | ~v_1922 | ~v_3299 | ~v_3298 | v_4160;
assign x_2715 = v_13 | v_9 | v_18 | v_17 | v_16 | v_15 | v_136 | v_135 | v_134 | ~v_3292 | v_137 | v_161 | v_182 | ~v_599 | ~v_598 | ~v_3291 | ~v_3290 | ~v_233 | ~v_232 | ~v_405 | ~v_404 | ~v_597 | ~v_596 | ~v_1868 | ~v_4130 | ~v_1867 | ~v_4129 | ~v_1866 | ~v_1865 | ~v_4128 | ~v_1864 | ~v_4127 | ~v_1863 | ~v_3289 | ~v_3288 | ~v_3287 | ~v_3286 | ~v_3285 | ~v_1920 | ~v_1919 | ~v_1918 | ~v_1917 | ~v_3284 | ~v_3283 | v_4159;
assign x_2716 = v_4158 | ~v_4155;
assign x_2717 = v_4158 | ~v_4156;
assign x_2718 = v_4158 | ~v_4157;
assign x_2719 = v_103 | v_101 | v_97 | v_99 | v_102 | v_171 | v_170 | v_169 | v_148 | v_147 | v_184 | v_181 | ~v_483 | ~v_482 | ~v_481 | ~v_480 | ~v_345 | ~v_479 | ~v_478 | ~v_344 | ~v_1962 | ~v_4140 | ~v_1961 | ~v_4139 | ~v_1896 | ~v_1960 | ~v_4138 | ~v_1959 | ~v_4137 | ~v_1893 | ~v_3386 | ~v_3385 | ~v_3318 | ~v_3384 | ~v_3383 | ~v_3315 | ~v_1914 | ~v_1913 | ~v_1912 | ~v_1911 | ~v_3438 | ~v_3437 | ~v_3436 | ~v_3435 | v_4157;
assign x_2720 = v_55 | v_61 | v_60 | v_59 | v_57 | v_180 | v_143 | v_142 | v_167 | v_166 | v_165 | v_183 | ~v_3381 | ~v_3380 | ~v_468 | ~v_467 | ~v_466 | ~v_465 | ~v_330 | ~v_464 | ~v_463 | ~v_329 | ~v_1957 | ~v_4135 | ~v_1956 | ~v_4134 | ~v_1881 | ~v_1955 | ~v_4133 | ~v_1954 | ~v_4132 | ~v_1878 | ~v_3303 | ~v_3379 | ~v_3378 | ~v_3300 | ~v_1909 | ~v_1908 | ~v_1907 | ~v_1906 | ~v_3433 | ~v_3432 | ~v_3431 | ~v_3430 | v_4156;
assign x_2721 = v_18 | v_17 | v_16 | v_14 | v_12 | ~v_453 | ~v_452 | v_135 | v_134 | v_179 | v_163 | v_162 | v_161 | v_182 | ~v_451 | ~v_450 | ~v_315 | ~v_449 | ~v_448 | ~v_314 | ~v_1952 | ~v_4130 | ~v_1951 | ~v_4129 | ~v_1866 | ~v_1950 | ~v_4128 | ~v_1949 | ~v_4127 | ~v_1863 | ~v_3376 | ~v_3375 | ~v_3288 | ~v_3374 | ~v_3373 | ~v_3285 | ~v_1904 | ~v_1903 | ~v_1902 | ~v_1901 | ~v_3428 | ~v_3427 | ~v_3426 | ~v_3425 | v_4155;
assign x_2722 = v_4154 | ~v_4151;
assign x_2723 = v_4154 | ~v_4152;
assign x_2724 = v_4154 | ~v_4153;
assign x_2725 = v_103 | v_101 | v_96 | v_102 | v_171 | v_170 | v_169 | v_150 | v_149 | v_147 | v_184 | v_181 | ~v_391 | ~v_390 | ~v_387 | ~v_386 | ~v_345 | ~v_344 | ~v_385 | ~v_384 | ~v_4140 | ~v_4139 | ~v_1896 | ~v_4138 | ~v_4137 | ~v_1893 | ~v_3318 | ~v_3315 | ~v_1946 | ~v_1945 | ~v_1944 | ~v_1943 | ~v_3354 | ~v_3353 | ~v_3352 | ~v_3351 | ~v_1914 | ~v_1913 | ~v_1912 | ~v_1911 | ~v_3438 | ~v_3437 | ~v_3436 | ~v_3435 | v_4153;
assign x_2726 = v_54 | v_61 | v_60 | v_59 | v_144 | v_180 | v_145 | v_142 | v_167 | v_166 | v_165 | v_183 | ~v_376 | ~v_375 | ~v_372 | ~v_371 | ~v_330 | ~v_329 | ~v_370 | ~v_369 | ~v_4135 | ~v_4134 | ~v_1881 | ~v_4133 | ~v_4132 | ~v_1878 | ~v_3303 | ~v_3300 | ~v_1941 | ~v_1940 | ~v_1939 | ~v_1938 | ~v_3349 | ~v_3348 | ~v_3347 | ~v_3346 | ~v_1909 | ~v_1908 | ~v_1907 | ~v_1906 | ~v_3433 | ~v_3432 | ~v_3431 | ~v_3430 | v_4152;
assign x_2727 = v_18 | v_17 | v_16 | v_11 | v_136 | v_134 | v_137 | v_179 | v_163 | v_162 | v_161 | v_182 | ~v_361 | ~v_360 | ~v_357 | ~v_356 | ~v_315 | ~v_314 | ~v_355 | ~v_354 | ~v_4130 | ~v_4129 | ~v_1866 | ~v_4128 | ~v_4127 | ~v_1863 | ~v_3288 | ~v_3285 | ~v_1936 | ~v_1935 | ~v_1934 | ~v_1933 | ~v_3344 | ~v_3343 | ~v_3342 | ~v_3341 | ~v_1904 | ~v_1903 | ~v_1902 | ~v_1901 | ~v_3428 | ~v_3427 | ~v_3426 | ~v_3425 | v_4151;
assign x_2728 = v_4150 | ~v_4147;
assign x_2729 = v_4150 | ~v_4148;
assign x_2730 = v_4150 | ~v_4149;
assign x_2731 = v_101 | v_102 | v_172 | v_171 | v_170 | v_169 | v_150 | v_149 | v_148 | v_147 | v_184 | v_181 | ~v_3322 | ~v_3321 | ~v_437 | ~v_436 | ~v_435 | ~v_434 | ~v_345 | ~v_344 | ~v_433 | ~v_432 | ~v_4140 | ~v_4139 | ~v_1896 | ~v_4138 | ~v_4137 | ~v_1893 | ~v_3318 | ~v_3315 | ~v_1930 | ~v_1929 | ~v_1928 | ~v_1927 | ~v_3314 | ~v_3313 | ~v_1914 | ~v_1913 | ~v_1912 | ~v_1911 | ~v_3438 | ~v_3437 | ~v_3436 | ~v_3435 | v_4149;
assign x_2732 = v_60 | v_59 | v_144 | v_180 | v_145 | v_143 | v_142 | v_168 | v_167 | v_166 | v_165 | v_183 | ~v_3307 | ~v_3306 | ~v_422 | ~v_421 | ~v_420 | ~v_419 | ~v_330 | ~v_329 | ~v_418 | ~v_417 | ~v_4135 | ~v_4134 | ~v_1881 | ~v_4133 | ~v_4132 | ~v_1878 | ~v_3303 | ~v_3300 | ~v_1925 | ~v_1924 | ~v_1923 | ~v_1922 | ~v_3299 | ~v_3298 | ~v_1909 | ~v_1908 | ~v_1907 | ~v_1906 | ~v_3433 | ~v_3432 | ~v_3431 | ~v_3430 | v_4148;
assign x_2733 = v_17 | v_16 | v_136 | v_135 | v_134 | v_137 | v_179 | v_164 | v_163 | v_162 | v_161 | v_182 | ~v_3291 | ~v_3290 | ~v_407 | ~v_406 | ~v_405 | ~v_404 | ~v_315 | ~v_314 | ~v_403 | ~v_402 | ~v_4130 | ~v_4129 | ~v_1866 | ~v_4128 | ~v_4127 | ~v_1863 | ~v_3288 | ~v_3285 | ~v_1920 | ~v_1919 | ~v_1918 | ~v_1917 | ~v_3284 | ~v_3283 | ~v_1904 | ~v_1903 | ~v_1902 | ~v_1901 | ~v_3428 | ~v_3427 | ~v_3426 | ~v_3425 | v_4147;
assign x_2734 = v_4146 | ~v_4143;
assign x_2735 = v_4146 | ~v_4144;
assign x_2736 = v_4146 | ~v_4145;
assign x_2737 = v_103 | v_95 | v_102 | v_171 | v_170 | v_169 | v_160 | v_150 | v_149 | v_148 | v_184 | v_181 | ~v_297 | ~v_296 | ~v_345 | ~v_344 | ~v_343 | ~v_342 | ~v_341 | ~v_340 | ~v_4140 | ~v_4139 | ~v_1896 | ~v_4138 | ~v_4137 | ~v_1893 | ~v_3318 | ~v_3315 | ~v_1892 | ~v_1891 | ~v_1890 | ~v_1889 | ~v_3370 | ~v_3369 | ~v_3368 | ~v_3367 | ~v_1914 | ~v_1913 | ~v_1912 | ~v_1911 | ~v_3438 | ~v_3437 | ~v_3436 | ~v_3435 | v_4145;
assign x_2738 = v_53 | v_61 | v_60 | v_144 | v_180 | v_159 | v_145 | v_143 | v_167 | v_166 | v_165 | v_183 | ~v_264 | ~v_263 | ~v_330 | ~v_329 | ~v_328 | ~v_327 | ~v_326 | ~v_325 | ~v_4135 | ~v_4134 | ~v_1881 | ~v_4133 | ~v_4132 | ~v_1878 | ~v_3303 | ~v_3300 | ~v_1877 | ~v_1876 | ~v_1875 | ~v_1874 | ~v_3365 | ~v_3364 | ~v_3363 | ~v_3362 | ~v_1909 | ~v_1908 | ~v_1907 | ~v_1906 | ~v_3433 | ~v_3432 | ~v_3431 | ~v_3430 | v_4144;
assign x_2739 = v_18 | v_17 | v_10 | v_136 | v_135 | v_137 | v_179 | v_163 | v_162 | v_161 | v_155 | v_182 | ~v_231 | ~v_230 | ~v_315 | ~v_314 | ~v_313 | ~v_312 | ~v_311 | ~v_310 | ~v_4130 | ~v_4129 | ~v_1866 | ~v_4128 | ~v_4127 | ~v_1863 | ~v_3288 | ~v_3285 | ~v_1862 | ~v_1861 | ~v_1860 | ~v_1859 | ~v_3360 | ~v_3359 | ~v_3358 | ~v_3357 | ~v_1904 | ~v_1903 | ~v_1902 | ~v_1901 | ~v_3428 | ~v_3427 | ~v_3426 | ~v_3425 | v_4143;
assign x_2740 = v_4142 | ~v_4131;
assign x_2741 = v_4142 | ~v_4136;
assign x_2742 = v_4142 | ~v_4141;
assign x_2743 = v_98 | v_103 | v_100 | v_94 | v_102 | v_169 | v_160 | v_150 | v_149 | v_148 | v_147 | v_184 | ~v_299 | ~v_298 | ~v_297 | ~v_296 | ~v_295 | ~v_294 | ~v_293 | ~v_292 | ~v_1898 | ~v_4140 | ~v_1897 | ~v_4139 | ~v_1896 | ~v_1895 | ~v_4138 | ~v_1894 | ~v_4137 | ~v_1893 | ~v_3320 | ~v_3319 | ~v_3318 | ~v_3317 | ~v_3316 | ~v_3315 | ~v_1892 | ~v_1891 | ~v_1890 | ~v_1889 | ~v_3370 | ~v_3369 | ~v_3368 | ~v_3367 | v_4141;
assign x_2744 = v_4140 | v_139;
assign x_2745 = v_4140 | v_123;
assign x_2746 = v_4139 | v_140;
assign x_2747 = v_4139 | v_120;
assign x_2748 = v_4138 | ~v_139;
assign x_2749 = v_4138 | v_108;
assign x_2750 = v_4137 | ~v_140;
assign x_2751 = v_4137 | v_105;
assign x_2752 = v_56 | v_61 | v_52 | v_60 | v_58 | v_144 | v_159 | v_145 | v_143 | v_142 | v_165 | v_183 | ~v_3305 | ~v_266 | ~v_265 | ~v_264 | ~v_263 | ~v_262 | ~v_261 | ~v_260 | ~v_259 | ~v_1883 | ~v_4135 | ~v_1882 | ~v_4134 | ~v_1881 | ~v_1880 | ~v_4133 | ~v_1879 | ~v_4132 | ~v_1878 | ~v_3304 | ~v_3303 | ~v_3302 | ~v_3301 | ~v_3300 | ~v_1877 | ~v_1876 | ~v_1875 | ~v_1874 | ~v_3365 | ~v_3364 | ~v_3363 | ~v_3362 | v_4136;
assign x_2753 = v_4135 | v_139;
assign x_2754 = v_4135 | v_81;
assign x_2755 = v_4134 | v_140;
assign x_2756 = v_4134 | v_78;
assign x_2757 = v_4133 | ~v_139;
assign x_2758 = v_4133 | v_66;
assign x_2759 = v_4132 | ~v_140;
assign x_2760 = v_4132 | v_63;
assign x_2761 = v_13 | v_9 | v_18 | v_17 | v_15 | v_136 | v_135 | v_134 | ~v_3292 | v_137 | v_161 | v_155 | v_182 | ~v_233 | ~v_232 | ~v_231 | ~v_230 | ~v_229 | ~v_228 | ~v_227 | ~v_226 | ~v_1868 | ~v_4130 | ~v_1867 | ~v_4129 | ~v_1866 | ~v_1865 | ~v_4128 | ~v_1864 | ~v_4127 | ~v_1863 | ~v_3289 | ~v_3288 | ~v_3287 | ~v_3286 | ~v_3285 | ~v_1862 | ~v_1861 | ~v_1860 | ~v_1859 | ~v_3360 | ~v_3359 | ~v_3358 | ~v_3357 | v_4131;
assign x_2762 = v_4130 | v_139;
assign x_2763 = v_4130 | v_39;
assign x_2764 = v_4129 | v_140;
assign x_2765 = v_4129 | v_36;
assign x_2766 = v_4128 | ~v_139;
assign x_2767 = v_4128 | v_24;
assign x_2768 = v_4127 | ~v_140;
assign x_2769 = v_4127 | v_21;
assign x_2770 = v_4126 | ~v_4124;
assign x_2771 = v_4126 | ~v_4125;
assign x_2772 = v_4126 | ~v_2219;
assign x_2773 = v_4126 | ~v_2220;
assign x_2774 = v_4126 | ~v_140;
assign x_2775 = v_4126 | ~v_139;
assign x_2776 = ~v_189 | ~v_1276 | v_4125;
assign x_2777 = ~v_195 | ~v_197 | v_4124;
assign x_2778 = v_4123 | ~v_4042;
assign x_2779 = v_4123 | ~v_4122;
assign x_2780 = v_140 | v_139 | ~v_4121 | ~v_2405 | ~v_2404 | ~v_4044 | ~v_4043 | v_4122;
assign x_2781 = v_4121 | ~v_4060;
assign x_2782 = v_4121 | ~v_4064;
assign x_2783 = v_4121 | ~v_4068;
assign x_2784 = v_4121 | ~v_4072;
assign x_2785 = v_4121 | ~v_4076;
assign x_2786 = v_4121 | ~v_4080;
assign x_2787 = v_4121 | ~v_4084;
assign x_2788 = v_4121 | ~v_4088;
assign x_2789 = v_4121 | ~v_4092;
assign x_2790 = v_4121 | ~v_4096;
assign x_2791 = v_4121 | ~v_4100;
assign x_2792 = v_4121 | ~v_4104;
assign x_2793 = v_4121 | ~v_4108;
assign x_2794 = v_4121 | ~v_4112;
assign x_2795 = v_4121 | ~v_4116;
assign x_2796 = v_4121 | ~v_4120;
assign x_2797 = v_4121 | ~v_1263;
assign x_2798 = v_4121 | ~v_1264;
assign x_2799 = v_4121 | ~v_1265;
assign x_2800 = v_4121 | ~v_1266;
assign x_2801 = ~v_4119 | ~v_4118 | ~v_4117 | v_4120;
assign x_2802 = v_4119 | ~v_3133;
assign x_2803 = v_4119 | ~v_3134;
assign x_2804 = v_4119 | ~v_3199;
assign x_2805 = v_4119 | ~v_3135;
assign x_2806 = v_4119 | ~v_839;
assign x_2807 = v_4119 | ~v_3200;
assign x_2808 = v_4119 | ~v_1257;
assign x_2809 = v_4119 | ~v_1023;
assign x_2810 = v_4119 | ~v_3136;
assign x_2811 = v_4119 | ~v_3137;
assign x_2812 = v_4119 | ~v_3201;
assign x_2813 = v_4119 | ~v_3138;
assign x_2814 = v_4119 | ~v_840;
assign x_2815 = v_4119 | ~v_3202;
assign x_2816 = v_4119 | ~v_1258;
assign x_2817 = v_4119 | ~v_1024;
assign x_2818 = v_4119 | ~v_4055;
assign x_2819 = v_4119 | ~v_4056;
assign x_2820 = v_4119 | ~v_2446;
assign x_2821 = v_4119 | ~v_2447;
assign x_2822 = v_4119 | ~v_2512;
assign x_2823 = v_4119 | ~v_2448;
assign x_2824 = v_4119 | ~v_2513;
assign x_2825 = v_4119 | ~v_4057;
assign x_2826 = v_4119 | ~v_4058;
assign x_2827 = v_4119 | ~v_2449;
assign x_2828 = v_4119 | ~v_2450;
assign x_2829 = v_4119 | ~v_2514;
assign x_2830 = v_4119 | ~v_2451;
assign x_2831 = v_4119 | ~v_2515;
assign x_2832 = v_4119 | ~v_184;
assign x_2833 = v_4119 | ~v_170;
assign x_2834 = v_4119 | ~v_149;
assign x_2835 = v_4119 | ~v_1259;
assign x_2836 = v_4119 | ~v_1260;
assign x_2837 = v_4119 | ~v_103;
assign x_2838 = v_4119 | ~v_102;
assign x_2839 = v_4119 | ~v_101;
assign x_2840 = v_4119 | ~v_100;
assign x_2841 = v_4119 | ~v_99;
assign x_2842 = v_4119 | ~v_98;
assign x_2843 = v_4119 | ~v_96;
assign x_2844 = v_4119 | ~v_95;
assign x_2845 = v_4119 | ~v_93;
assign x_2846 = v_4118 | ~v_3118;
assign x_2847 = v_4118 | ~v_3119;
assign x_2848 = v_4118 | ~v_3194;
assign x_2849 = v_4118 | ~v_3120;
assign x_2850 = v_4118 | ~v_806;
assign x_2851 = v_4118 | ~v_3195;
assign x_2852 = v_4118 | ~v_1252;
assign x_2853 = v_4118 | ~v_1008;
assign x_2854 = v_4118 | ~v_3121;
assign x_2855 = v_4118 | ~v_3122;
assign x_2856 = v_4118 | ~v_1253;
assign x_2857 = v_4118 | ~v_1009;
assign x_2858 = v_4118 | ~v_4050;
assign x_2859 = v_4118 | ~v_4051;
assign x_2860 = v_4118 | ~v_2431;
assign x_2861 = v_4118 | ~v_2432;
assign x_2862 = v_4118 | ~v_2507;
assign x_2863 = v_4118 | ~v_2433;
assign x_2864 = v_4118 | ~v_2508;
assign x_2865 = v_4118 | ~v_4052;
assign x_2866 = v_4118 | ~v_4053;
assign x_2867 = v_4118 | ~v_2434;
assign x_2868 = v_4118 | ~v_2435;
assign x_2869 = v_4118 | ~v_2509;
assign x_2870 = v_4118 | ~v_2436;
assign x_2871 = v_4118 | ~v_2510;
assign x_2872 = v_4118 | ~v_3123;
assign x_2873 = v_4118 | ~v_807;
assign x_2874 = v_4118 | ~v_3196;
assign x_2875 = v_4118 | ~v_183;
assign x_2876 = v_4118 | ~v_166;
assign x_2877 = v_4118 | ~v_144;
assign x_2878 = v_4118 | ~v_3197;
assign x_2879 = v_4118 | ~v_1254;
assign x_2880 = v_4118 | ~v_1255;
assign x_2881 = v_4118 | ~v_61;
assign x_2882 = v_4118 | ~v_60;
assign x_2883 = v_4118 | ~v_59;
assign x_2884 = v_4118 | ~v_58;
assign x_2885 = v_4118 | ~v_57;
assign x_2886 = v_4118 | ~v_56;
assign x_2887 = v_4118 | ~v_54;
assign x_2888 = v_4118 | ~v_53;
assign x_2889 = v_4118 | ~v_51;
assign x_2890 = v_4117 | ~v_3103;
assign x_2891 = v_4117 | ~v_3189;
assign x_2892 = v_4117 | ~v_3104;
assign x_2893 = v_4117 | ~v_773;
assign x_2894 = v_4117 | ~v_3190;
assign x_2895 = v_4117 | ~v_3105;
assign x_2896 = v_4117 | ~v_3191;
assign x_2897 = v_4117 | ~v_3106;
assign x_2898 = v_4117 | ~v_774;
assign x_2899 = v_4117 | ~v_3192;
assign x_2900 = v_4117 | ~v_4045;
assign x_2901 = v_4117 | ~v_4046;
assign x_2902 = v_4117 | ~v_2416;
assign x_2903 = v_4117 | ~v_2417;
assign x_2904 = v_4117 | ~v_2502;
assign x_2905 = v_4117 | ~v_2418;
assign x_2906 = v_4117 | ~v_2503;
assign x_2907 = v_4117 | ~v_4047;
assign x_2908 = v_4117 | ~v_4048;
assign x_2909 = v_4117 | ~v_2419;
assign x_2910 = v_4117 | ~v_2420;
assign x_2911 = v_4117 | ~v_2504;
assign x_2912 = v_4117 | ~v_2421;
assign x_2913 = v_4117 | ~v_2505;
assign x_2914 = v_4117 | ~v_182;
assign x_2915 = v_4117 | ~v_162;
assign x_2916 = v_4117 | ~v_1247;
assign x_2917 = v_4117 | ~v_1248;
assign x_2918 = v_4117 | ~v_136;
assign x_2919 = v_4117 | ~v_3107;
assign x_2920 = v_4117 | ~v_1249;
assign x_2921 = v_4117 | ~v_993;
assign x_2922 = v_4117 | ~v_3108;
assign x_2923 = v_4117 | ~v_1250;
assign x_2924 = v_4117 | ~v_994;
assign x_2925 = v_4117 | ~v_18;
assign x_2926 = v_4117 | ~v_17;
assign x_2927 = v_4117 | ~v_16;
assign x_2928 = v_4117 | ~v_15;
assign x_2929 = v_4117 | ~v_14;
assign x_2930 = v_4117 | ~v_13;
assign x_2931 = v_4117 | ~v_11;
assign x_2932 = v_4117 | ~v_10;
assign x_2933 = v_4117 | ~v_8;
assign x_2934 = ~v_4115 | ~v_4114 | ~v_4113 | v_4116;
assign x_2935 = v_4115 | ~v_3219;
assign x_2936 = v_4115 | ~v_3220;
assign x_2937 = v_4115 | ~v_1085;
assign x_2938 = v_4115 | ~v_1131;
assign x_2939 = v_4115 | ~v_1132;
assign x_2940 = v_4115 | ~v_3221;
assign x_2941 = v_4115 | ~v_3222;
assign x_2942 = v_4115 | ~v_1086;
assign x_2943 = v_4115 | ~v_1133;
assign x_2944 = v_4115 | ~v_1134;
assign x_2945 = v_4115 | ~v_2532;
assign x_2946 = v_4115 | ~v_2533;
assign x_2947 = v_4115 | ~v_2534;
assign x_2948 = v_4115 | ~v_2535;
assign x_2949 = v_4115 | ~v_3133;
assign x_2950 = v_4115 | ~v_3199;
assign x_2951 = v_4115 | ~v_3200;
assign x_2952 = v_4115 | ~v_1023;
assign x_2953 = v_4115 | ~v_3136;
assign x_2954 = v_4115 | ~v_3201;
assign x_2955 = v_4115 | ~v_3202;
assign x_2956 = v_4115 | ~v_1024;
assign x_2957 = v_4115 | ~v_4055;
assign x_2958 = v_4115 | ~v_4056;
assign x_2959 = v_4115 | ~v_2446;
assign x_2960 = v_4115 | ~v_2512;
assign x_2961 = v_4115 | ~v_2513;
assign x_2962 = v_4115 | ~v_4057;
assign x_2963 = v_4115 | ~v_4058;
assign x_2964 = v_4115 | ~v_2449;
assign x_2965 = v_4115 | ~v_2514;
assign x_2966 = v_4115 | ~v_2515;
assign x_2967 = v_4115 | ~v_184;
assign x_2968 = v_4115 | ~v_172;
assign x_2969 = v_4115 | ~v_171;
assign x_2970 = v_4115 | ~v_169;
assign x_2971 = v_4115 | ~v_149;
assign x_2972 = v_4115 | ~v_147;
assign x_2973 = v_4115 | ~v_102;
assign x_2974 = v_4115 | ~v_101;
assign x_2975 = v_4115 | ~v_100;
assign x_2976 = v_4115 | ~v_99;
assign x_2977 = v_4115 | ~v_96;
assign x_2978 = v_4115 | ~v_94;
assign x_2979 = v_4114 | ~v_3214;
assign x_2980 = v_4114 | ~v_3215;
assign x_2981 = v_4114 | ~v_1070;
assign x_2982 = v_4114 | ~v_1126;
assign x_2983 = v_4114 | ~v_1127;
assign x_2984 = v_4114 | ~v_3216;
assign x_2985 = v_4114 | ~v_3217;
assign x_2986 = v_4114 | ~v_1071;
assign x_2987 = v_4114 | ~v_1128;
assign x_2988 = v_4114 | ~v_1129;
assign x_2989 = v_4114 | ~v_2527;
assign x_2990 = v_4114 | ~v_2528;
assign x_2991 = v_4114 | ~v_2529;
assign x_2992 = v_4114 | ~v_2530;
assign x_2993 = v_4114 | ~v_3118;
assign x_2994 = v_4114 | ~v_3194;
assign x_2995 = v_4114 | ~v_3195;
assign x_2996 = v_4114 | ~v_1008;
assign x_2997 = v_4114 | ~v_3121;
assign x_2998 = v_4114 | ~v_1009;
assign x_2999 = v_4114 | ~v_4050;
assign x_3000 = v_4114 | ~v_4051;
assign x_3001 = v_4114 | ~v_2431;
assign x_3002 = v_4114 | ~v_2507;
assign x_3003 = v_4114 | ~v_2508;
assign x_3004 = v_4114 | ~v_4052;
assign x_3005 = v_4114 | ~v_4053;
assign x_3006 = v_4114 | ~v_2434;
assign x_3007 = v_4114 | ~v_2509;
assign x_3008 = v_4114 | ~v_2510;
assign x_3009 = v_4114 | ~v_3196;
assign x_3010 = v_4114 | ~v_183;
assign x_3011 = v_4114 | ~v_168;
assign x_3012 = v_4114 | ~v_167;
assign x_3013 = v_4114 | ~v_165;
assign x_3014 = v_4114 | ~v_144;
assign x_3015 = v_4114 | ~v_142;
assign x_3016 = v_4114 | ~v_3197;
assign x_3017 = v_4114 | ~v_60;
assign x_3018 = v_4114 | ~v_59;
assign x_3019 = v_4114 | ~v_58;
assign x_3020 = v_4114 | ~v_57;
assign x_3021 = v_4114 | ~v_54;
assign x_3022 = v_4114 | ~v_52;
assign x_3023 = v_4113 | ~v_3209;
assign x_3024 = v_4113 | ~v_3210;
assign x_3025 = v_4113 | ~v_1055;
assign x_3026 = v_4113 | ~v_1121;
assign x_3027 = v_4113 | ~v_1122;
assign x_3028 = v_4113 | ~v_3211;
assign x_3029 = v_4113 | ~v_3212;
assign x_3030 = v_4113 | ~v_1056;
assign x_3031 = v_4113 | ~v_1123;
assign x_3032 = v_4113 | ~v_1124;
assign x_3033 = v_4113 | ~v_2522;
assign x_3034 = v_4113 | ~v_2523;
assign x_3035 = v_4113 | ~v_2524;
assign x_3036 = v_4113 | ~v_2525;
assign x_3037 = v_4113 | ~v_3189;
assign x_3038 = v_4113 | ~v_3190;
assign x_3039 = v_4113 | ~v_3191;
assign x_3040 = v_4113 | ~v_3192;
assign x_3041 = v_4113 | ~v_4045;
assign x_3042 = v_4113 | ~v_4046;
assign x_3043 = v_4113 | ~v_2416;
assign x_3044 = v_4113 | ~v_2502;
assign x_3045 = v_4113 | ~v_2503;
assign x_3046 = v_4113 | ~v_4047;
assign x_3047 = v_4113 | ~v_4048;
assign x_3048 = v_4113 | ~v_2419;
assign x_3049 = v_4113 | ~v_2504;
assign x_3050 = v_4113 | ~v_2505;
assign x_3051 = v_4113 | ~v_182;
assign x_3052 = v_4113 | ~v_164;
assign x_3053 = v_4113 | ~v_163;
assign x_3054 = v_4113 | ~v_161;
assign x_3055 = v_4113 | ~v_136;
assign x_3056 = v_4113 | ~v_134;
assign x_3057 = v_4113 | ~v_3107;
assign x_3058 = v_4113 | ~v_993;
assign x_3059 = v_4113 | ~v_3108;
assign x_3060 = v_4113 | ~v_994;
assign x_3061 = v_4113 | ~v_17;
assign x_3062 = v_4113 | ~v_16;
assign x_3063 = v_4113 | ~v_15;
assign x_3064 = v_4113 | ~v_14;
assign x_3065 = v_4113 | ~v_11;
assign x_3066 = v_4113 | ~v_9;
assign x_3067 = ~v_4111 | ~v_4110 | ~v_4109 | v_4112;
assign x_3068 = v_4111 | ~v_3167;
assign x_3069 = v_4111 | ~v_3168;
assign x_3070 = v_4111 | ~v_927;
assign x_3071 = v_4111 | ~v_3169;
assign x_3072 = v_4111 | ~v_3170;
assign x_3073 = v_4111 | ~v_928;
assign x_3074 = v_4111 | ~v_1099;
assign x_3075 = v_4111 | ~v_1100;
assign x_3076 = v_4111 | ~v_1101;
assign x_3077 = v_4111 | ~v_1102;
assign x_3078 = v_4111 | ~v_2480;
assign x_3079 = v_4111 | ~v_2481;
assign x_3080 = v_4111 | ~v_2482;
assign x_3081 = v_4111 | ~v_2483;
assign x_3082 = v_4111 | ~v_3219;
assign x_3083 = v_4111 | ~v_3220;
assign x_3084 = v_4111 | ~v_1085;
assign x_3085 = v_4111 | ~v_3221;
assign x_3086 = v_4111 | ~v_3222;
assign x_3087 = v_4111 | ~v_1086;
assign x_3088 = v_4111 | ~v_2532;
assign x_3089 = v_4111 | ~v_2533;
assign x_3090 = v_4111 | ~v_2534;
assign x_3091 = v_4111 | ~v_2535;
assign x_3092 = v_4111 | ~v_3133;
assign x_3093 = v_4111 | ~v_3136;
assign x_3094 = v_4111 | ~v_4055;
assign x_3095 = v_4111 | ~v_4056;
assign x_3096 = v_4111 | ~v_2446;
assign x_3097 = v_4111 | ~v_4057;
assign x_3098 = v_4111 | ~v_4058;
assign x_3099 = v_4111 | ~v_2449;
assign x_3100 = v_4111 | ~v_184;
assign x_3101 = v_4111 | ~v_171;
assign x_3102 = v_4111 | ~v_169;
assign x_3103 = v_4111 | ~v_150;
assign x_3104 = v_4111 | ~v_148;
assign x_3105 = v_4111 | ~v_103;
assign x_3106 = v_4111 | ~v_102;
assign x_3107 = v_4111 | ~v_101;
assign x_3108 = v_4111 | ~v_100;
assign x_3109 = v_4111 | ~v_97;
assign x_3110 = v_4111 | ~v_95;
assign x_3111 = v_4111 | ~v_94;
assign x_3112 = v_4110 | ~v_3162;
assign x_3113 = v_4110 | ~v_3163;
assign x_3114 = v_4110 | ~v_912;
assign x_3115 = v_4110 | ~v_3164;
assign x_3116 = v_4110 | ~v_3165;
assign x_3117 = v_4110 | ~v_913;
assign x_3118 = v_4110 | ~v_1094;
assign x_3119 = v_4110 | ~v_1095;
assign x_3120 = v_4110 | ~v_1096;
assign x_3121 = v_4110 | ~v_1097;
assign x_3122 = v_4110 | ~v_2475;
assign x_3123 = v_4110 | ~v_2476;
assign x_3124 = v_4110 | ~v_2477;
assign x_3125 = v_4110 | ~v_2478;
assign x_3126 = v_4110 | ~v_3214;
assign x_3127 = v_4110 | ~v_3215;
assign x_3128 = v_4110 | ~v_1070;
assign x_3129 = v_4110 | ~v_3216;
assign x_3130 = v_4110 | ~v_3217;
assign x_3131 = v_4110 | ~v_1071;
assign x_3132 = v_4110 | ~v_2527;
assign x_3133 = v_4110 | ~v_2528;
assign x_3134 = v_4110 | ~v_2529;
assign x_3135 = v_4110 | ~v_2530;
assign x_3136 = v_4110 | ~v_3118;
assign x_3137 = v_4110 | ~v_3121;
assign x_3138 = v_4110 | ~v_4050;
assign x_3139 = v_4110 | ~v_4051;
assign x_3140 = v_4110 | ~v_2431;
assign x_3141 = v_4110 | ~v_4052;
assign x_3142 = v_4110 | ~v_4053;
assign x_3143 = v_4110 | ~v_2434;
assign x_3144 = v_4110 | ~v_183;
assign x_3145 = v_4110 | ~v_167;
assign x_3146 = v_4110 | ~v_165;
assign x_3147 = v_4110 | ~v_145;
assign x_3148 = v_4110 | ~v_143;
assign x_3149 = v_4110 | ~v_61;
assign x_3150 = v_4110 | ~v_60;
assign x_3151 = v_4110 | ~v_59;
assign x_3152 = v_4110 | ~v_58;
assign x_3153 = v_4110 | ~v_55;
assign x_3154 = v_4110 | ~v_53;
assign x_3155 = v_4110 | ~v_52;
assign x_3156 = v_4109 | ~v_3157;
assign x_3157 = v_4109 | ~v_3158;
assign x_3158 = v_4109 | ~v_897;
assign x_3159 = v_4109 | ~v_3159;
assign x_3160 = v_4109 | ~v_3160;
assign x_3161 = v_4109 | ~v_898;
assign x_3162 = v_4109 | ~v_1089;
assign x_3163 = v_4109 | ~v_1090;
assign x_3164 = v_4109 | ~v_1091;
assign x_3165 = v_4109 | ~v_1092;
assign x_3166 = v_4109 | ~v_2470;
assign x_3167 = v_4109 | ~v_2471;
assign x_3168 = v_4109 | ~v_2472;
assign x_3169 = v_4109 | ~v_2473;
assign x_3170 = v_4109 | ~v_3209;
assign x_3171 = v_4109 | ~v_3210;
assign x_3172 = v_4109 | ~v_1055;
assign x_3173 = v_4109 | ~v_3211;
assign x_3174 = v_4109 | ~v_3212;
assign x_3175 = v_4109 | ~v_1056;
assign x_3176 = v_4109 | ~v_2522;
assign x_3177 = v_4109 | ~v_2523;
assign x_3178 = v_4109 | ~v_2524;
assign x_3179 = v_4109 | ~v_2525;
assign x_3180 = v_4109 | ~v_4045;
assign x_3181 = v_4109 | ~v_4046;
assign x_3182 = v_4109 | ~v_2416;
assign x_3183 = v_4109 | ~v_4047;
assign x_3184 = v_4109 | ~v_4048;
assign x_3185 = v_4109 | ~v_2419;
assign x_3186 = v_4109 | ~v_182;
assign x_3187 = v_4109 | ~v_163;
assign x_3188 = v_4109 | ~v_161;
assign x_3189 = v_4109 | ~v_137;
assign x_3190 = v_4109 | ~v_135;
assign x_3191 = v_4109 | ~v_3107;
assign x_3192 = v_4109 | ~v_3108;
assign x_3193 = v_4109 | ~v_18;
assign x_3194 = v_4109 | ~v_17;
assign x_3195 = v_4109 | ~v_16;
assign x_3196 = v_4109 | ~v_15;
assign x_3197 = v_4109 | ~v_12;
assign x_3198 = v_4109 | ~v_10;
assign x_3199 = v_4109 | ~v_9;
assign x_3200 = ~v_4107 | ~v_4106 | ~v_4105 | v_4108;
assign x_3201 = v_4107 | ~v_3129;
assign x_3202 = v_4107 | ~v_3130;
assign x_3203 = v_4107 | ~v_975;
assign x_3204 = v_4107 | ~v_3131;
assign x_3205 = v_4107 | ~v_3132;
assign x_3206 = v_4107 | ~v_976;
assign x_3207 = v_4107 | ~v_1115;
assign x_3208 = v_4107 | ~v_1116;
assign x_3209 = v_4107 | ~v_2442;
assign x_3210 = v_4107 | ~v_2443;
assign x_3211 = v_4107 | ~v_2444;
assign x_3212 = v_4107 | ~v_2445;
assign x_3213 = v_4107 | ~v_3219;
assign x_3214 = v_4107 | ~v_3220;
assign x_3215 = v_4107 | ~v_1085;
assign x_3216 = v_4107 | ~v_3221;
assign x_3217 = v_4107 | ~v_3222;
assign x_3218 = v_4107 | ~v_1086;
assign x_3219 = v_4107 | ~v_2532;
assign x_3220 = v_4107 | ~v_2533;
assign x_3221 = v_4107 | ~v_2534;
assign x_3222 = v_4107 | ~v_2535;
assign x_3223 = v_4107 | ~v_3133;
assign x_3224 = v_4107 | ~v_3136;
assign x_3225 = v_4107 | ~v_4055;
assign x_3226 = v_4107 | ~v_4056;
assign x_3227 = v_4107 | ~v_2446;
assign x_3228 = v_4107 | ~v_4057;
assign x_3229 = v_4107 | ~v_4058;
assign x_3230 = v_4107 | ~v_2449;
assign x_3231 = v_4107 | ~v_1117;
assign x_3232 = v_4107 | ~v_1118;
assign x_3233 = v_4107 | ~v_184;
assign x_3234 = v_4107 | ~v_171;
assign x_3235 = v_4107 | ~v_169;
assign x_3236 = v_4107 | ~v_151;
assign x_3237 = v_4107 | ~v_150;
assign x_3238 = v_4107 | ~v_149;
assign x_3239 = v_4107 | ~v_148;
assign x_3240 = v_4107 | ~v_147;
assign x_3241 = v_4107 | ~v_103;
assign x_3242 = v_4107 | ~v_101;
assign x_3243 = v_4107 | ~v_100;
assign x_3244 = v_4107 | ~v_94;
assign x_3245 = v_4106 | ~v_3114;
assign x_3246 = v_4106 | ~v_3115;
assign x_3247 = v_4106 | ~v_960;
assign x_3248 = v_4106 | ~v_3116;
assign x_3249 = v_4106 | ~v_3117;
assign x_3250 = v_4106 | ~v_961;
assign x_3251 = v_4106 | ~v_1110;
assign x_3252 = v_4106 | ~v_1111;
assign x_3253 = v_4106 | ~v_2427;
assign x_3254 = v_4106 | ~v_2428;
assign x_3255 = v_4106 | ~v_2429;
assign x_3256 = v_4106 | ~v_2430;
assign x_3257 = v_4106 | ~v_3214;
assign x_3258 = v_4106 | ~v_3215;
assign x_3259 = v_4106 | ~v_1070;
assign x_3260 = v_4106 | ~v_3216;
assign x_3261 = v_4106 | ~v_3217;
assign x_3262 = v_4106 | ~v_1071;
assign x_3263 = v_4106 | ~v_2527;
assign x_3264 = v_4106 | ~v_2528;
assign x_3265 = v_4106 | ~v_2529;
assign x_3266 = v_4106 | ~v_2530;
assign x_3267 = v_4106 | ~v_3118;
assign x_3268 = v_4106 | ~v_3121;
assign x_3269 = v_4106 | ~v_4050;
assign x_3270 = v_4106 | ~v_4051;
assign x_3271 = v_4106 | ~v_2431;
assign x_3272 = v_4106 | ~v_4052;
assign x_3273 = v_4106 | ~v_4053;
assign x_3274 = v_4106 | ~v_2434;
assign x_3275 = v_4106 | ~v_1112;
assign x_3276 = v_4106 | ~v_1113;
assign x_3277 = v_4106 | ~v_183;
assign x_3278 = v_4106 | ~v_167;
assign x_3279 = v_4106 | ~v_165;
assign x_3280 = v_4106 | ~v_146;
assign x_3281 = v_4106 | ~v_145;
assign x_3282 = v_4106 | ~v_144;
assign x_3283 = v_4106 | ~v_143;
assign x_3284 = v_4106 | ~v_142;
assign x_3285 = v_4106 | ~v_61;
assign x_3286 = v_4106 | ~v_59;
assign x_3287 = v_4106 | ~v_58;
assign x_3288 = v_4106 | ~v_52;
assign x_3289 = v_4105 | ~v_3099;
assign x_3290 = v_4105 | ~v_3100;
assign x_3291 = v_4105 | ~v_945;
assign x_3292 = v_4105 | ~v_3101;
assign x_3293 = v_4105 | ~v_3102;
assign x_3294 = v_4105 | ~v_946;
assign x_3295 = v_4105 | ~v_1105;
assign x_3296 = v_4105 | ~v_1106;
assign x_3297 = v_4105 | ~v_2412;
assign x_3298 = v_4105 | ~v_2413;
assign x_3299 = v_4105 | ~v_2414;
assign x_3300 = v_4105 | ~v_2415;
assign x_3301 = v_4105 | ~v_3209;
assign x_3302 = v_4105 | ~v_3210;
assign x_3303 = v_4105 | ~v_1055;
assign x_3304 = v_4105 | ~v_3211;
assign x_3305 = v_4105 | ~v_3212;
assign x_3306 = v_4105 | ~v_1056;
assign x_3307 = v_4105 | ~v_2522;
assign x_3308 = v_4105 | ~v_2523;
assign x_3309 = v_4105 | ~v_2524;
assign x_3310 = v_4105 | ~v_2525;
assign x_3311 = v_4105 | ~v_4045;
assign x_3312 = v_4105 | ~v_4046;
assign x_3313 = v_4105 | ~v_2416;
assign x_3314 = v_4105 | ~v_4047;
assign x_3315 = v_4105 | ~v_4048;
assign x_3316 = v_4105 | ~v_2419;
assign x_3317 = v_4105 | ~v_1107;
assign x_3318 = v_4105 | ~v_1108;
assign x_3319 = v_4105 | ~v_182;
assign x_3320 = v_4105 | ~v_163;
assign x_3321 = v_4105 | ~v_161;
assign x_3322 = v_4105 | ~v_138;
assign x_3323 = v_4105 | ~v_137;
assign x_3324 = v_4105 | ~v_136;
assign x_3325 = v_4105 | ~v_135;
assign x_3326 = v_4105 | ~v_134;
assign x_3327 = v_4105 | ~v_3107;
assign x_3328 = v_4105 | ~v_3108;
assign x_3329 = v_4105 | ~v_18;
assign x_3330 = v_4105 | ~v_16;
assign x_3331 = v_4105 | ~v_15;
assign x_3332 = v_4105 | ~v_9;
assign x_3333 = ~v_4103 | ~v_4102 | ~v_4101 | v_4104;
assign x_3334 = v_4103 | ~v_3183;
assign x_3335 = v_4103 | ~v_3184;
assign x_3336 = v_4103 | ~v_837;
assign x_3337 = v_4103 | ~v_3185;
assign x_3338 = v_4103 | ~v_3186;
assign x_3339 = v_4103 | ~v_838;
assign x_3340 = v_4103 | ~v_1081;
assign x_3341 = v_4103 | ~v_1082;
assign x_3342 = v_4103 | ~v_1083;
assign x_3343 = v_4103 | ~v_1084;
assign x_3344 = v_4103 | ~v_2496;
assign x_3345 = v_4103 | ~v_2497;
assign x_3346 = v_4103 | ~v_2498;
assign x_3347 = v_4103 | ~v_2499;
assign x_3348 = v_4103 | ~v_3219;
assign x_3349 = v_4103 | ~v_3220;
assign x_3350 = v_4103 | ~v_1085;
assign x_3351 = v_4103 | ~v_3221;
assign x_3352 = v_4103 | ~v_3222;
assign x_3353 = v_4103 | ~v_1086;
assign x_3354 = v_4103 | ~v_2532;
assign x_3355 = v_4103 | ~v_2533;
assign x_3356 = v_4103 | ~v_2534;
assign x_3357 = v_4103 | ~v_2535;
assign x_3358 = v_4103 | ~v_3133;
assign x_3359 = v_4103 | ~v_3136;
assign x_3360 = v_4103 | ~v_4055;
assign x_3361 = v_4103 | ~v_4056;
assign x_3362 = v_4103 | ~v_2446;
assign x_3363 = v_4103 | ~v_4057;
assign x_3364 = v_4103 | ~v_4058;
assign x_3365 = v_4103 | ~v_2449;
assign x_3366 = v_4103 | ~v_184;
assign x_3367 = v_4103 | ~v_171;
assign x_3368 = v_4103 | ~v_169;
assign x_3369 = v_4103 | ~v_160;
assign x_3370 = v_4103 | ~v_150;
assign x_3371 = v_4103 | ~v_149;
assign x_3372 = v_4103 | ~v_148;
assign x_3373 = v_4103 | ~v_147;
assign x_3374 = v_4103 | ~v_103;
assign x_3375 = v_4103 | ~v_102;
assign x_3376 = v_4103 | ~v_100;
assign x_3377 = v_4103 | ~v_94;
assign x_3378 = v_4102 | ~v_3178;
assign x_3379 = v_4102 | ~v_3179;
assign x_3380 = v_4102 | ~v_804;
assign x_3381 = v_4102 | ~v_3180;
assign x_3382 = v_4102 | ~v_3181;
assign x_3383 = v_4102 | ~v_805;
assign x_3384 = v_4102 | ~v_1066;
assign x_3385 = v_4102 | ~v_1067;
assign x_3386 = v_4102 | ~v_1068;
assign x_3387 = v_4102 | ~v_1069;
assign x_3388 = v_4102 | ~v_2491;
assign x_3389 = v_4102 | ~v_2492;
assign x_3390 = v_4102 | ~v_2493;
assign x_3391 = v_4102 | ~v_2494;
assign x_3392 = v_4102 | ~v_3214;
assign x_3393 = v_4102 | ~v_3215;
assign x_3394 = v_4102 | ~v_1070;
assign x_3395 = v_4102 | ~v_3216;
assign x_3396 = v_4102 | ~v_3217;
assign x_3397 = v_4102 | ~v_1071;
assign x_3398 = v_4102 | ~v_2527;
assign x_3399 = v_4102 | ~v_2528;
assign x_3400 = v_4102 | ~v_2529;
assign x_3401 = v_4102 | ~v_2530;
assign x_3402 = v_4102 | ~v_3118;
assign x_3403 = v_4102 | ~v_3121;
assign x_3404 = v_4102 | ~v_4050;
assign x_3405 = v_4102 | ~v_4051;
assign x_3406 = v_4102 | ~v_2431;
assign x_3407 = v_4102 | ~v_4052;
assign x_3408 = v_4102 | ~v_4053;
assign x_3409 = v_4102 | ~v_2434;
assign x_3410 = v_4102 | ~v_183;
assign x_3411 = v_4102 | ~v_167;
assign x_3412 = v_4102 | ~v_165;
assign x_3413 = v_4102 | ~v_159;
assign x_3414 = v_4102 | ~v_145;
assign x_3415 = v_4102 | ~v_144;
assign x_3416 = v_4102 | ~v_143;
assign x_3417 = v_4102 | ~v_142;
assign x_3418 = v_4102 | ~v_61;
assign x_3419 = v_4102 | ~v_60;
assign x_3420 = v_4102 | ~v_58;
assign x_3421 = v_4102 | ~v_52;
assign x_3422 = v_4101 | ~v_3173;
assign x_3423 = v_4101 | ~v_3174;
assign x_3424 = v_4101 | ~v_771;
assign x_3425 = v_4101 | ~v_3175;
assign x_3426 = v_4101 | ~v_3176;
assign x_3427 = v_4101 | ~v_772;
assign x_3428 = v_4101 | ~v_1051;
assign x_3429 = v_4101 | ~v_1052;
assign x_3430 = v_4101 | ~v_1053;
assign x_3431 = v_4101 | ~v_1054;
assign x_3432 = v_4101 | ~v_2486;
assign x_3433 = v_4101 | ~v_2487;
assign x_3434 = v_4101 | ~v_2488;
assign x_3435 = v_4101 | ~v_2489;
assign x_3436 = v_4101 | ~v_3209;
assign x_3437 = v_4101 | ~v_3210;
assign x_3438 = v_4101 | ~v_1055;
assign x_3439 = v_4101 | ~v_3211;
assign x_3440 = v_4101 | ~v_3212;
assign x_3441 = v_4101 | ~v_1056;
assign x_3442 = v_4101 | ~v_2522;
assign x_3443 = v_4101 | ~v_2523;
assign x_3444 = v_4101 | ~v_2524;
assign x_3445 = v_4101 | ~v_2525;
assign x_3446 = v_4101 | ~v_4045;
assign x_3447 = v_4101 | ~v_4046;
assign x_3448 = v_4101 | ~v_2416;
assign x_3449 = v_4101 | ~v_4047;
assign x_3450 = v_4101 | ~v_4048;
assign x_3451 = v_4101 | ~v_2419;
assign x_3452 = v_4101 | ~v_182;
assign x_3453 = v_4101 | ~v_163;
assign x_3454 = v_4101 | ~v_161;
assign x_3455 = v_4101 | ~v_155;
assign x_3456 = v_4101 | ~v_137;
assign x_3457 = v_4101 | ~v_136;
assign x_3458 = v_4101 | ~v_135;
assign x_3459 = v_4101 | ~v_134;
assign x_3460 = v_4101 | ~v_3107;
assign x_3461 = v_4101 | ~v_3108;
assign x_3462 = v_4101 | ~v_18;
assign x_3463 = v_4101 | ~v_17;
assign x_3464 = v_4101 | ~v_15;
assign x_3465 = v_4101 | ~v_9;
assign x_3466 = ~v_4099 | ~v_4098 | ~v_4097 | v_4100;
assign x_3467 = v_4099 | ~v_1037;
assign x_3468 = v_4099 | ~v_1038;
assign x_3469 = v_4099 | ~v_1039;
assign x_3470 = v_4099 | ~v_1040;
assign x_3471 = v_4099 | ~v_3167;
assign x_3472 = v_4099 | ~v_3168;
assign x_3473 = v_4099 | ~v_927;
assign x_3474 = v_4099 | ~v_3169;
assign x_3475 = v_4099 | ~v_3170;
assign x_3476 = v_4099 | ~v_928;
assign x_3477 = v_4099 | ~v_2480;
assign x_3478 = v_4099 | ~v_2481;
assign x_3479 = v_4099 | ~v_2482;
assign x_3480 = v_4099 | ~v_2483;
assign x_3481 = v_4099 | ~v_3133;
assign x_3482 = v_4099 | ~v_3134;
assign x_3483 = v_4099 | ~v_3135;
assign x_3484 = v_4099 | ~v_839;
assign x_3485 = v_4099 | ~v_3136;
assign x_3486 = v_4099 | ~v_3137;
assign x_3487 = v_4099 | ~v_3138;
assign x_3488 = v_4099 | ~v_840;
assign x_3489 = v_4099 | ~v_4055;
assign x_3490 = v_4099 | ~v_4056;
assign x_3491 = v_4099 | ~v_2446;
assign x_3492 = v_4099 | ~v_2447;
assign x_3493 = v_4099 | ~v_2448;
assign x_3494 = v_4099 | ~v_4057;
assign x_3495 = v_4099 | ~v_4058;
assign x_3496 = v_4099 | ~v_2449;
assign x_3497 = v_4099 | ~v_2450;
assign x_3498 = v_4099 | ~v_2451;
assign x_3499 = v_4099 | ~v_184;
assign x_3500 = v_4099 | ~v_170;
assign x_3501 = v_4099 | ~v_151;
assign x_3502 = v_4099 | ~v_150;
assign x_3503 = v_4099 | ~v_148;
assign x_3504 = v_4099 | ~v_147;
assign x_3505 = v_4099 | ~v_103;
assign x_3506 = v_4099 | ~v_101;
assign x_3507 = v_4099 | ~v_100;
assign x_3508 = v_4099 | ~v_98;
assign x_3509 = v_4099 | ~v_97;
assign x_3510 = v_4099 | ~v_93;
assign x_3511 = v_4098 | ~v_1032;
assign x_3512 = v_4098 | ~v_1033;
assign x_3513 = v_4098 | ~v_1034;
assign x_3514 = v_4098 | ~v_1035;
assign x_3515 = v_4098 | ~v_3162;
assign x_3516 = v_4098 | ~v_3163;
assign x_3517 = v_4098 | ~v_912;
assign x_3518 = v_4098 | ~v_3164;
assign x_3519 = v_4098 | ~v_3165;
assign x_3520 = v_4098 | ~v_913;
assign x_3521 = v_4098 | ~v_2475;
assign x_3522 = v_4098 | ~v_2476;
assign x_3523 = v_4098 | ~v_2477;
assign x_3524 = v_4098 | ~v_2478;
assign x_3525 = v_4098 | ~v_3118;
assign x_3526 = v_4098 | ~v_3119;
assign x_3527 = v_4098 | ~v_3120;
assign x_3528 = v_4098 | ~v_806;
assign x_3529 = v_4098 | ~v_3121;
assign x_3530 = v_4098 | ~v_3122;
assign x_3531 = v_4098 | ~v_4050;
assign x_3532 = v_4098 | ~v_4051;
assign x_3533 = v_4098 | ~v_2431;
assign x_3534 = v_4098 | ~v_2432;
assign x_3535 = v_4098 | ~v_2433;
assign x_3536 = v_4098 | ~v_4052;
assign x_3537 = v_4098 | ~v_4053;
assign x_3538 = v_4098 | ~v_2434;
assign x_3539 = v_4098 | ~v_2435;
assign x_3540 = v_4098 | ~v_2436;
assign x_3541 = v_4098 | ~v_3123;
assign x_3542 = v_4098 | ~v_807;
assign x_3543 = v_4098 | ~v_183;
assign x_3544 = v_4098 | ~v_166;
assign x_3545 = v_4098 | ~v_146;
assign x_3546 = v_4098 | ~v_145;
assign x_3547 = v_4098 | ~v_143;
assign x_3548 = v_4098 | ~v_142;
assign x_3549 = v_4098 | ~v_61;
assign x_3550 = v_4098 | ~v_59;
assign x_3551 = v_4098 | ~v_58;
assign x_3552 = v_4098 | ~v_56;
assign x_3553 = v_4098 | ~v_55;
assign x_3554 = v_4098 | ~v_51;
assign x_3555 = v_4097 | ~v_1027;
assign x_3556 = v_4097 | ~v_1028;
assign x_3557 = v_4097 | ~v_1029;
assign x_3558 = v_4097 | ~v_1030;
assign x_3559 = v_4097 | ~v_3157;
assign x_3560 = v_4097 | ~v_3158;
assign x_3561 = v_4097 | ~v_897;
assign x_3562 = v_4097 | ~v_3159;
assign x_3563 = v_4097 | ~v_3160;
assign x_3564 = v_4097 | ~v_898;
assign x_3565 = v_4097 | ~v_2470;
assign x_3566 = v_4097 | ~v_2471;
assign x_3567 = v_4097 | ~v_2472;
assign x_3568 = v_4097 | ~v_2473;
assign x_3569 = v_4097 | ~v_3103;
assign x_3570 = v_4097 | ~v_3104;
assign x_3571 = v_4097 | ~v_773;
assign x_3572 = v_4097 | ~v_3105;
assign x_3573 = v_4097 | ~v_3106;
assign x_3574 = v_4097 | ~v_774;
assign x_3575 = v_4097 | ~v_4045;
assign x_3576 = v_4097 | ~v_4046;
assign x_3577 = v_4097 | ~v_2416;
assign x_3578 = v_4097 | ~v_2417;
assign x_3579 = v_4097 | ~v_2418;
assign x_3580 = v_4097 | ~v_4047;
assign x_3581 = v_4097 | ~v_4048;
assign x_3582 = v_4097 | ~v_2419;
assign x_3583 = v_4097 | ~v_2420;
assign x_3584 = v_4097 | ~v_2421;
assign x_3585 = v_4097 | ~v_182;
assign x_3586 = v_4097 | ~v_162;
assign x_3587 = v_4097 | ~v_138;
assign x_3588 = v_4097 | ~v_137;
assign x_3589 = v_4097 | ~v_135;
assign x_3590 = v_4097 | ~v_134;
assign x_3591 = v_4097 | ~v_3107;
assign x_3592 = v_4097 | ~v_3108;
assign x_3593 = v_4097 | ~v_18;
assign x_3594 = v_4097 | ~v_16;
assign x_3595 = v_4097 | ~v_15;
assign x_3596 = v_4097 | ~v_13;
assign x_3597 = v_4097 | ~v_12;
assign x_3598 = v_4097 | ~v_8;
assign x_3599 = ~v_4095 | ~v_4094 | ~v_4093 | v_4096;
assign x_3600 = v_4095 | ~v_3151;
assign x_3601 = v_4095 | ~v_3152;
assign x_3602 = v_4095 | ~v_1193;
assign x_3603 = v_4095 | ~v_1241;
assign x_3604 = v_4095 | ~v_3153;
assign x_3605 = v_4095 | ~v_3154;
assign x_3606 = v_4095 | ~v_1194;
assign x_3607 = v_4095 | ~v_1242;
assign x_3608 = v_4095 | ~v_2464;
assign x_3609 = v_4095 | ~v_2465;
assign x_3610 = v_4095 | ~v_2466;
assign x_3611 = v_4095 | ~v_2467;
assign x_3612 = v_4095 | ~v_3133;
assign x_3613 = v_4095 | ~v_3199;
assign x_3614 = v_4095 | ~v_3200;
assign x_3615 = v_4095 | ~v_1023;
assign x_3616 = v_4095 | ~v_3136;
assign x_3617 = v_4095 | ~v_3201;
assign x_3618 = v_4095 | ~v_3202;
assign x_3619 = v_4095 | ~v_1024;
assign x_3620 = v_4095 | ~v_4055;
assign x_3621 = v_4095 | ~v_4056;
assign x_3622 = v_4095 | ~v_2446;
assign x_3623 = v_4095 | ~v_2512;
assign x_3624 = v_4095 | ~v_2513;
assign x_3625 = v_4095 | ~v_4057;
assign x_3626 = v_4095 | ~v_4058;
assign x_3627 = v_4095 | ~v_2449;
assign x_3628 = v_4095 | ~v_2514;
assign x_3629 = v_4095 | ~v_2515;
assign x_3630 = v_4095 | ~v_1243;
assign x_3631 = v_4095 | ~v_1244;
assign x_3632 = v_4095 | ~v_184;
assign x_3633 = v_4095 | ~v_171;
assign x_3634 = v_4095 | ~v_170;
assign x_3635 = v_4095 | ~v_169;
assign x_3636 = v_4095 | ~v_149;
assign x_3637 = v_4095 | ~v_147;
assign x_3638 = v_4095 | ~v_103;
assign x_3639 = v_4095 | ~v_102;
assign x_3640 = v_4095 | ~v_101;
assign x_3641 = v_4095 | ~v_100;
assign x_3642 = v_4095 | ~v_99;
assign x_3643 = v_4095 | ~v_96;
assign x_3644 = v_4094 | ~v_3146;
assign x_3645 = v_4094 | ~v_3147;
assign x_3646 = v_4094 | ~v_1178;
assign x_3647 = v_4094 | ~v_1236;
assign x_3648 = v_4094 | ~v_3148;
assign x_3649 = v_4094 | ~v_3149;
assign x_3650 = v_4094 | ~v_1179;
assign x_3651 = v_4094 | ~v_1237;
assign x_3652 = v_4094 | ~v_2459;
assign x_3653 = v_4094 | ~v_2460;
assign x_3654 = v_4094 | ~v_2461;
assign x_3655 = v_4094 | ~v_2462;
assign x_3656 = v_4094 | ~v_3118;
assign x_3657 = v_4094 | ~v_3194;
assign x_3658 = v_4094 | ~v_3195;
assign x_3659 = v_4094 | ~v_1008;
assign x_3660 = v_4094 | ~v_3121;
assign x_3661 = v_4094 | ~v_1009;
assign x_3662 = v_4094 | ~v_4050;
assign x_3663 = v_4094 | ~v_4051;
assign x_3664 = v_4094 | ~v_2431;
assign x_3665 = v_4094 | ~v_2507;
assign x_3666 = v_4094 | ~v_2508;
assign x_3667 = v_4094 | ~v_4052;
assign x_3668 = v_4094 | ~v_4053;
assign x_3669 = v_4094 | ~v_2434;
assign x_3670 = v_4094 | ~v_2509;
assign x_3671 = v_4094 | ~v_2510;
assign x_3672 = v_4094 | ~v_3196;
assign x_3673 = v_4094 | ~v_1238;
assign x_3674 = v_4094 | ~v_1239;
assign x_3675 = v_4094 | ~v_183;
assign x_3676 = v_4094 | ~v_167;
assign x_3677 = v_4094 | ~v_166;
assign x_3678 = v_4094 | ~v_165;
assign x_3679 = v_4094 | ~v_144;
assign x_3680 = v_4094 | ~v_142;
assign x_3681 = v_4094 | ~v_3197;
assign x_3682 = v_4094 | ~v_61;
assign x_3683 = v_4094 | ~v_60;
assign x_3684 = v_4094 | ~v_59;
assign x_3685 = v_4094 | ~v_58;
assign x_3686 = v_4094 | ~v_57;
assign x_3687 = v_4094 | ~v_54;
assign x_3688 = v_4093 | ~v_3141;
assign x_3689 = v_4093 | ~v_3142;
assign x_3690 = v_4093 | ~v_1163;
assign x_3691 = v_4093 | ~v_1231;
assign x_3692 = v_4093 | ~v_3143;
assign x_3693 = v_4093 | ~v_3144;
assign x_3694 = v_4093 | ~v_1164;
assign x_3695 = v_4093 | ~v_1232;
assign x_3696 = v_4093 | ~v_2454;
assign x_3697 = v_4093 | ~v_2455;
assign x_3698 = v_4093 | ~v_2456;
assign x_3699 = v_4093 | ~v_2457;
assign x_3700 = v_4093 | ~v_3189;
assign x_3701 = v_4093 | ~v_3190;
assign x_3702 = v_4093 | ~v_3191;
assign x_3703 = v_4093 | ~v_3192;
assign x_3704 = v_4093 | ~v_4045;
assign x_3705 = v_4093 | ~v_4046;
assign x_3706 = v_4093 | ~v_2416;
assign x_3707 = v_4093 | ~v_2502;
assign x_3708 = v_4093 | ~v_2503;
assign x_3709 = v_4093 | ~v_4047;
assign x_3710 = v_4093 | ~v_4048;
assign x_3711 = v_4093 | ~v_2419;
assign x_3712 = v_4093 | ~v_2504;
assign x_3713 = v_4093 | ~v_2505;
assign x_3714 = v_4093 | ~v_1233;
assign x_3715 = v_4093 | ~v_1234;
assign x_3716 = v_4093 | ~v_182;
assign x_3717 = v_4093 | ~v_163;
assign x_3718 = v_4093 | ~v_162;
assign x_3719 = v_4093 | ~v_161;
assign x_3720 = v_4093 | ~v_136;
assign x_3721 = v_4093 | ~v_134;
assign x_3722 = v_4093 | ~v_3107;
assign x_3723 = v_4093 | ~v_993;
assign x_3724 = v_4093 | ~v_3108;
assign x_3725 = v_4093 | ~v_994;
assign x_3726 = v_4093 | ~v_18;
assign x_3727 = v_4093 | ~v_17;
assign x_3728 = v_4093 | ~v_16;
assign x_3729 = v_4093 | ~v_15;
assign x_3730 = v_4093 | ~v_14;
assign x_3731 = v_4093 | ~v_11;
assign x_3732 = ~v_4091 | ~v_4090 | ~v_4089 | v_4092;
assign x_3733 = v_4091 | ~v_1209;
assign x_3734 = v_4091 | ~v_1210;
assign x_3735 = v_4091 | ~v_3151;
assign x_3736 = v_4091 | ~v_3152;
assign x_3737 = v_4091 | ~v_1193;
assign x_3738 = v_4091 | ~v_3153;
assign x_3739 = v_4091 | ~v_3154;
assign x_3740 = v_4091 | ~v_1194;
assign x_3741 = v_4091 | ~v_2464;
assign x_3742 = v_4091 | ~v_2465;
assign x_3743 = v_4091 | ~v_2466;
assign x_3744 = v_4091 | ~v_2467;
assign x_3745 = v_4091 | ~v_3167;
assign x_3746 = v_4091 | ~v_3168;
assign x_3747 = v_4091 | ~v_927;
assign x_3748 = v_4091 | ~v_3169;
assign x_3749 = v_4091 | ~v_3170;
assign x_3750 = v_4091 | ~v_928;
assign x_3751 = v_4091 | ~v_2480;
assign x_3752 = v_4091 | ~v_2481;
assign x_3753 = v_4091 | ~v_2482;
assign x_3754 = v_4091 | ~v_2483;
assign x_3755 = v_4091 | ~v_3133;
assign x_3756 = v_4091 | ~v_3136;
assign x_3757 = v_4091 | ~v_4055;
assign x_3758 = v_4091 | ~v_4056;
assign x_3759 = v_4091 | ~v_2446;
assign x_3760 = v_4091 | ~v_4057;
assign x_3761 = v_4091 | ~v_4058;
assign x_3762 = v_4091 | ~v_2449;
assign x_3763 = v_4091 | ~v_1211;
assign x_3764 = v_4091 | ~v_1212;
assign x_3765 = v_4091 | ~v_184;
assign x_3766 = v_4091 | ~v_172;
assign x_3767 = v_4091 | ~v_171;
assign x_3768 = v_4091 | ~v_170;
assign x_3769 = v_4091 | ~v_169;
assign x_3770 = v_4091 | ~v_150;
assign x_3771 = v_4091 | ~v_148;
assign x_3772 = v_4091 | ~v_147;
assign x_3773 = v_4091 | ~v_102;
assign x_3774 = v_4091 | ~v_101;
assign x_3775 = v_4091 | ~v_100;
assign x_3776 = v_4091 | ~v_97;
assign x_3777 = v_4090 | ~v_1204;
assign x_3778 = v_4090 | ~v_1205;
assign x_3779 = v_4090 | ~v_3146;
assign x_3780 = v_4090 | ~v_3147;
assign x_3781 = v_4090 | ~v_1178;
assign x_3782 = v_4090 | ~v_3148;
assign x_3783 = v_4090 | ~v_3149;
assign x_3784 = v_4090 | ~v_1179;
assign x_3785 = v_4090 | ~v_2459;
assign x_3786 = v_4090 | ~v_2460;
assign x_3787 = v_4090 | ~v_2461;
assign x_3788 = v_4090 | ~v_2462;
assign x_3789 = v_4090 | ~v_3162;
assign x_3790 = v_4090 | ~v_3163;
assign x_3791 = v_4090 | ~v_912;
assign x_3792 = v_4090 | ~v_3164;
assign x_3793 = v_4090 | ~v_3165;
assign x_3794 = v_4090 | ~v_913;
assign x_3795 = v_4090 | ~v_2475;
assign x_3796 = v_4090 | ~v_2476;
assign x_3797 = v_4090 | ~v_2477;
assign x_3798 = v_4090 | ~v_2478;
assign x_3799 = v_4090 | ~v_3118;
assign x_3800 = v_4090 | ~v_3121;
assign x_3801 = v_4090 | ~v_4050;
assign x_3802 = v_4090 | ~v_4051;
assign x_3803 = v_4090 | ~v_2431;
assign x_3804 = v_4090 | ~v_4052;
assign x_3805 = v_4090 | ~v_4053;
assign x_3806 = v_4090 | ~v_2434;
assign x_3807 = v_4090 | ~v_1206;
assign x_3808 = v_4090 | ~v_1207;
assign x_3809 = v_4090 | ~v_183;
assign x_3810 = v_4090 | ~v_168;
assign x_3811 = v_4090 | ~v_167;
assign x_3812 = v_4090 | ~v_166;
assign x_3813 = v_4090 | ~v_165;
assign x_3814 = v_4090 | ~v_145;
assign x_3815 = v_4090 | ~v_143;
assign x_3816 = v_4090 | ~v_142;
assign x_3817 = v_4090 | ~v_60;
assign x_3818 = v_4090 | ~v_59;
assign x_3819 = v_4090 | ~v_58;
assign x_3820 = v_4090 | ~v_55;
assign x_3821 = v_4089 | ~v_1199;
assign x_3822 = v_4089 | ~v_1200;
assign x_3823 = v_4089 | ~v_3141;
assign x_3824 = v_4089 | ~v_3142;
assign x_3825 = v_4089 | ~v_1163;
assign x_3826 = v_4089 | ~v_3143;
assign x_3827 = v_4089 | ~v_3144;
assign x_3828 = v_4089 | ~v_1164;
assign x_3829 = v_4089 | ~v_2454;
assign x_3830 = v_4089 | ~v_2455;
assign x_3831 = v_4089 | ~v_2456;
assign x_3832 = v_4089 | ~v_2457;
assign x_3833 = v_4089 | ~v_3157;
assign x_3834 = v_4089 | ~v_3158;
assign x_3835 = v_4089 | ~v_897;
assign x_3836 = v_4089 | ~v_3159;
assign x_3837 = v_4089 | ~v_3160;
assign x_3838 = v_4089 | ~v_898;
assign x_3839 = v_4089 | ~v_2470;
assign x_3840 = v_4089 | ~v_2471;
assign x_3841 = v_4089 | ~v_2472;
assign x_3842 = v_4089 | ~v_2473;
assign x_3843 = v_4089 | ~v_4045;
assign x_3844 = v_4089 | ~v_4046;
assign x_3845 = v_4089 | ~v_2416;
assign x_3846 = v_4089 | ~v_4047;
assign x_3847 = v_4089 | ~v_4048;
assign x_3848 = v_4089 | ~v_2419;
assign x_3849 = v_4089 | ~v_1201;
assign x_3850 = v_4089 | ~v_1202;
assign x_3851 = v_4089 | ~v_182;
assign x_3852 = v_4089 | ~v_164;
assign x_3853 = v_4089 | ~v_163;
assign x_3854 = v_4089 | ~v_162;
assign x_3855 = v_4089 | ~v_161;
assign x_3856 = v_4089 | ~v_137;
assign x_3857 = v_4089 | ~v_135;
assign x_3858 = v_4089 | ~v_134;
assign x_3859 = v_4089 | ~v_3107;
assign x_3860 = v_4089 | ~v_3108;
assign x_3861 = v_4089 | ~v_17;
assign x_3862 = v_4089 | ~v_16;
assign x_3863 = v_4089 | ~v_15;
assign x_3864 = v_4089 | ~v_12;
assign x_3865 = ~v_4087 | ~v_4086 | ~v_4085 | v_4088;
assign x_3866 = v_4087 | ~v_1225;
assign x_3867 = v_4087 | ~v_1226;
assign x_3868 = v_4087 | ~v_1227;
assign x_3869 = v_4087 | ~v_1228;
assign x_3870 = v_4087 | ~v_3151;
assign x_3871 = v_4087 | ~v_3152;
assign x_3872 = v_4087 | ~v_1193;
assign x_3873 = v_4087 | ~v_3153;
assign x_3874 = v_4087 | ~v_3154;
assign x_3875 = v_4087 | ~v_1194;
assign x_3876 = v_4087 | ~v_2464;
assign x_3877 = v_4087 | ~v_2465;
assign x_3878 = v_4087 | ~v_2466;
assign x_3879 = v_4087 | ~v_2467;
assign x_3880 = v_4087 | ~v_3129;
assign x_3881 = v_4087 | ~v_3130;
assign x_3882 = v_4087 | ~v_975;
assign x_3883 = v_4087 | ~v_3131;
assign x_3884 = v_4087 | ~v_3132;
assign x_3885 = v_4087 | ~v_976;
assign x_3886 = v_4087 | ~v_2442;
assign x_3887 = v_4087 | ~v_2443;
assign x_3888 = v_4087 | ~v_2444;
assign x_3889 = v_4087 | ~v_2445;
assign x_3890 = v_4087 | ~v_3133;
assign x_3891 = v_4087 | ~v_3136;
assign x_3892 = v_4087 | ~v_4055;
assign x_3893 = v_4087 | ~v_4056;
assign x_3894 = v_4087 | ~v_2446;
assign x_3895 = v_4087 | ~v_4057;
assign x_3896 = v_4087 | ~v_4058;
assign x_3897 = v_4087 | ~v_2449;
assign x_3898 = v_4087 | ~v_184;
assign x_3899 = v_4087 | ~v_171;
assign x_3900 = v_4087 | ~v_170;
assign x_3901 = v_4087 | ~v_169;
assign x_3902 = v_4087 | ~v_150;
assign x_3903 = v_4087 | ~v_149;
assign x_3904 = v_4087 | ~v_148;
assign x_3905 = v_4087 | ~v_103;
assign x_3906 = v_4087 | ~v_102;
assign x_3907 = v_4087 | ~v_101;
assign x_3908 = v_4087 | ~v_100;
assign x_3909 = v_4087 | ~v_95;
assign x_3910 = v_4086 | ~v_1220;
assign x_3911 = v_4086 | ~v_1221;
assign x_3912 = v_4086 | ~v_1222;
assign x_3913 = v_4086 | ~v_1223;
assign x_3914 = v_4086 | ~v_3146;
assign x_3915 = v_4086 | ~v_3147;
assign x_3916 = v_4086 | ~v_1178;
assign x_3917 = v_4086 | ~v_3148;
assign x_3918 = v_4086 | ~v_3149;
assign x_3919 = v_4086 | ~v_1179;
assign x_3920 = v_4086 | ~v_2459;
assign x_3921 = v_4086 | ~v_2460;
assign x_3922 = v_4086 | ~v_2461;
assign x_3923 = v_4086 | ~v_2462;
assign x_3924 = v_4086 | ~v_3114;
assign x_3925 = v_4086 | ~v_3115;
assign x_3926 = v_4086 | ~v_960;
assign x_3927 = v_4086 | ~v_3116;
assign x_3928 = v_4086 | ~v_3117;
assign x_3929 = v_4086 | ~v_961;
assign x_3930 = v_4086 | ~v_2427;
assign x_3931 = v_4086 | ~v_2428;
assign x_3932 = v_4086 | ~v_2429;
assign x_3933 = v_4086 | ~v_2430;
assign x_3934 = v_4086 | ~v_3118;
assign x_3935 = v_4086 | ~v_3121;
assign x_3936 = v_4086 | ~v_4050;
assign x_3937 = v_4086 | ~v_4051;
assign x_3938 = v_4086 | ~v_2431;
assign x_3939 = v_4086 | ~v_4052;
assign x_3940 = v_4086 | ~v_4053;
assign x_3941 = v_4086 | ~v_2434;
assign x_3942 = v_4086 | ~v_183;
assign x_3943 = v_4086 | ~v_167;
assign x_3944 = v_4086 | ~v_166;
assign x_3945 = v_4086 | ~v_165;
assign x_3946 = v_4086 | ~v_145;
assign x_3947 = v_4086 | ~v_144;
assign x_3948 = v_4086 | ~v_143;
assign x_3949 = v_4086 | ~v_61;
assign x_3950 = v_4086 | ~v_60;
assign x_3951 = v_4086 | ~v_59;
assign x_3952 = v_4086 | ~v_58;
assign x_3953 = v_4086 | ~v_53;
assign x_3954 = v_4085 | ~v_1215;
assign x_3955 = v_4085 | ~v_1216;
assign x_3956 = v_4085 | ~v_1217;
assign x_3957 = v_4085 | ~v_1218;
assign x_3958 = v_4085 | ~v_3141;
assign x_3959 = v_4085 | ~v_3142;
assign x_3960 = v_4085 | ~v_1163;
assign x_3961 = v_4085 | ~v_3143;
assign x_3962 = v_4085 | ~v_3144;
assign x_3963 = v_4085 | ~v_1164;
assign x_3964 = v_4085 | ~v_2454;
assign x_3965 = v_4085 | ~v_2455;
assign x_3966 = v_4085 | ~v_2456;
assign x_3967 = v_4085 | ~v_2457;
assign x_3968 = v_4085 | ~v_3099;
assign x_3969 = v_4085 | ~v_3100;
assign x_3970 = v_4085 | ~v_945;
assign x_3971 = v_4085 | ~v_3101;
assign x_3972 = v_4085 | ~v_3102;
assign x_3973 = v_4085 | ~v_946;
assign x_3974 = v_4085 | ~v_2412;
assign x_3975 = v_4085 | ~v_2413;
assign x_3976 = v_4085 | ~v_2414;
assign x_3977 = v_4085 | ~v_2415;
assign x_3978 = v_4085 | ~v_4045;
assign x_3979 = v_4085 | ~v_4046;
assign x_3980 = v_4085 | ~v_2416;
assign x_3981 = v_4085 | ~v_4047;
assign x_3982 = v_4085 | ~v_4048;
assign x_3983 = v_4085 | ~v_2419;
assign x_3984 = v_4085 | ~v_182;
assign x_3985 = v_4085 | ~v_163;
assign x_3986 = v_4085 | ~v_162;
assign x_3987 = v_4085 | ~v_161;
assign x_3988 = v_4085 | ~v_137;
assign x_3989 = v_4085 | ~v_136;
assign x_3990 = v_4085 | ~v_135;
assign x_3991 = v_4085 | ~v_3107;
assign x_3992 = v_4085 | ~v_3108;
assign x_3993 = v_4085 | ~v_18;
assign x_3994 = v_4085 | ~v_17;
assign x_3995 = v_4085 | ~v_16;
assign x_3996 = v_4085 | ~v_15;
assign x_3997 = v_4085 | ~v_10;
assign x_3998 = ~v_4083 | ~v_4082 | ~v_4081 | v_4084;
assign x_3999 = v_4083 | ~v_1191;
assign x_4000 = v_4083 | ~v_1192;
assign x_4001 = v_4083 | ~v_3151;
assign x_4002 = v_4083 | ~v_3152;
assign x_4003 = v_4083 | ~v_1193;
assign x_4004 = v_4083 | ~v_3153;
assign x_4005 = v_4083 | ~v_3154;
assign x_4006 = v_4083 | ~v_1194;
assign x_4007 = v_4083 | ~v_2464;
assign x_4008 = v_4083 | ~v_2465;
assign x_4009 = v_4083 | ~v_2466;
assign x_4010 = v_4083 | ~v_2467;
assign x_4011 = v_4083 | ~v_3183;
assign x_4012 = v_4083 | ~v_3184;
assign x_4013 = v_4083 | ~v_837;
assign x_4014 = v_4083 | ~v_3185;
assign x_4015 = v_4083 | ~v_3186;
assign x_4016 = v_4083 | ~v_838;
assign x_4017 = v_4083 | ~v_2496;
assign x_4018 = v_4083 | ~v_2497;
assign x_4019 = v_4083 | ~v_2498;
assign x_4020 = v_4083 | ~v_2499;
assign x_4021 = v_4083 | ~v_3133;
assign x_4022 = v_4083 | ~v_3136;
assign x_4023 = v_4083 | ~v_4055;
assign x_4024 = v_4083 | ~v_4056;
assign x_4025 = v_4083 | ~v_2446;
assign x_4026 = v_4083 | ~v_4057;
assign x_4027 = v_4083 | ~v_4058;
assign x_4028 = v_4083 | ~v_2449;
assign x_4029 = v_4083 | ~v_1195;
assign x_4030 = v_4083 | ~v_1196;
assign x_4031 = v_4083 | ~v_184;
assign x_4032 = v_4083 | ~v_171;
assign x_4033 = v_4083 | ~v_170;
assign x_4034 = v_4083 | ~v_169;
assign x_4035 = v_4083 | ~v_160;
assign x_4036 = v_4083 | ~v_151;
assign x_4037 = v_4083 | ~v_150;
assign x_4038 = v_4083 | ~v_149;
assign x_4039 = v_4083 | ~v_148;
assign x_4040 = v_4083 | ~v_147;
assign x_4041 = v_4083 | ~v_103;
assign x_4042 = v_4083 | ~v_100;
assign x_4043 = v_4082 | ~v_1176;
assign x_4044 = v_4082 | ~v_1177;
assign x_4045 = v_4082 | ~v_3146;
assign x_4046 = v_4082 | ~v_3147;
assign x_4047 = v_4082 | ~v_1178;
assign x_4048 = v_4082 | ~v_3148;
assign x_4049 = v_4082 | ~v_3149;
assign x_4050 = v_4082 | ~v_1179;
assign x_4051 = v_4082 | ~v_2459;
assign x_4052 = v_4082 | ~v_2460;
assign x_4053 = v_4082 | ~v_2461;
assign x_4054 = v_4082 | ~v_2462;
assign x_4055 = v_4082 | ~v_3178;
assign x_4056 = v_4082 | ~v_3179;
assign x_4057 = v_4082 | ~v_804;
assign x_4058 = v_4082 | ~v_3180;
assign x_4059 = v_4082 | ~v_3181;
assign x_4060 = v_4082 | ~v_805;
assign x_4061 = v_4082 | ~v_2491;
assign x_4062 = v_4082 | ~v_2492;
assign x_4063 = v_4082 | ~v_2493;
assign x_4064 = v_4082 | ~v_2494;
assign x_4065 = v_4082 | ~v_3118;
assign x_4066 = v_4082 | ~v_3121;
assign x_4067 = v_4082 | ~v_4050;
assign x_4068 = v_4082 | ~v_4051;
assign x_4069 = v_4082 | ~v_2431;
assign x_4070 = v_4082 | ~v_4052;
assign x_4071 = v_4082 | ~v_4053;
assign x_4072 = v_4082 | ~v_2434;
assign x_4073 = v_4082 | ~v_1180;
assign x_4074 = v_4082 | ~v_1181;
assign x_4075 = v_4082 | ~v_183;
assign x_4076 = v_4082 | ~v_167;
assign x_4077 = v_4082 | ~v_166;
assign x_4078 = v_4082 | ~v_165;
assign x_4079 = v_4082 | ~v_159;
assign x_4080 = v_4082 | ~v_146;
assign x_4081 = v_4082 | ~v_145;
assign x_4082 = v_4082 | ~v_144;
assign x_4083 = v_4082 | ~v_143;
assign x_4084 = v_4082 | ~v_142;
assign x_4085 = v_4082 | ~v_61;
assign x_4086 = v_4082 | ~v_58;
assign x_4087 = v_4081 | ~v_1161;
assign x_4088 = v_4081 | ~v_1162;
assign x_4089 = v_4081 | ~v_3141;
assign x_4090 = v_4081 | ~v_3142;
assign x_4091 = v_4081 | ~v_1163;
assign x_4092 = v_4081 | ~v_3143;
assign x_4093 = v_4081 | ~v_3144;
assign x_4094 = v_4081 | ~v_1164;
assign x_4095 = v_4081 | ~v_2454;
assign x_4096 = v_4081 | ~v_2455;
assign x_4097 = v_4081 | ~v_2456;
assign x_4098 = v_4081 | ~v_2457;
assign x_4099 = v_4081 | ~v_3173;
assign x_4100 = v_4081 | ~v_3174;
assign x_4101 = v_4081 | ~v_771;
assign x_4102 = v_4081 | ~v_3175;
assign x_4103 = v_4081 | ~v_3176;
assign x_4104 = v_4081 | ~v_772;
assign x_4105 = v_4081 | ~v_2486;
assign x_4106 = v_4081 | ~v_2487;
assign x_4107 = v_4081 | ~v_2488;
assign x_4108 = v_4081 | ~v_2489;
assign x_4109 = v_4081 | ~v_4045;
assign x_4110 = v_4081 | ~v_4046;
assign x_4111 = v_4081 | ~v_2416;
assign x_4112 = v_4081 | ~v_4047;
assign x_4113 = v_4081 | ~v_4048;
assign x_4114 = v_4081 | ~v_2419;
assign x_4115 = v_4081 | ~v_1165;
assign x_4116 = v_4081 | ~v_1166;
assign x_4117 = v_4081 | ~v_182;
assign x_4118 = v_4081 | ~v_163;
assign x_4119 = v_4081 | ~v_162;
assign x_4120 = v_4081 | ~v_161;
assign x_4121 = v_4081 | ~v_155;
assign x_4122 = v_4081 | ~v_138;
assign x_4123 = v_4081 | ~v_137;
assign x_4124 = v_4081 | ~v_136;
assign x_4125 = v_4081 | ~v_135;
assign x_4126 = v_4081 | ~v_134;
assign x_4127 = v_4081 | ~v_3107;
assign x_4128 = v_4081 | ~v_3108;
assign x_4129 = v_4081 | ~v_18;
assign x_4130 = v_4081 | ~v_15;
assign x_4131 = ~v_4079 | ~v_4078 | ~v_4077 | v_4080;
assign x_4132 = v_4079 | ~v_1147;
assign x_4133 = v_4079 | ~v_1148;
assign x_4134 = v_4079 | ~v_3129;
assign x_4135 = v_4079 | ~v_3130;
assign x_4136 = v_4079 | ~v_975;
assign x_4137 = v_4079 | ~v_3131;
assign x_4138 = v_4079 | ~v_3132;
assign x_4139 = v_4079 | ~v_976;
assign x_4140 = v_4079 | ~v_2442;
assign x_4141 = v_4079 | ~v_2443;
assign x_4142 = v_4079 | ~v_2444;
assign x_4143 = v_4079 | ~v_2445;
assign x_4144 = v_4079 | ~v_3133;
assign x_4145 = v_4079 | ~v_3134;
assign x_4146 = v_4079 | ~v_3135;
assign x_4147 = v_4079 | ~v_839;
assign x_4148 = v_4079 | ~v_3136;
assign x_4149 = v_4079 | ~v_3137;
assign x_4150 = v_4079 | ~v_3138;
assign x_4151 = v_4079 | ~v_840;
assign x_4152 = v_4079 | ~v_4055;
assign x_4153 = v_4079 | ~v_4056;
assign x_4154 = v_4079 | ~v_2446;
assign x_4155 = v_4079 | ~v_2447;
assign x_4156 = v_4079 | ~v_2448;
assign x_4157 = v_4079 | ~v_4057;
assign x_4158 = v_4079 | ~v_4058;
assign x_4159 = v_4079 | ~v_2449;
assign x_4160 = v_4079 | ~v_2450;
assign x_4161 = v_4079 | ~v_2451;
assign x_4162 = v_4079 | ~v_1149;
assign x_4163 = v_4079 | ~v_1150;
assign x_4164 = v_4079 | ~v_184;
assign x_4165 = v_4079 | ~v_170;
assign x_4166 = v_4079 | ~v_150;
assign x_4167 = v_4079 | ~v_149;
assign x_4168 = v_4079 | ~v_148;
assign x_4169 = v_4079 | ~v_147;
assign x_4170 = v_4079 | ~v_103;
assign x_4171 = v_4079 | ~v_102;
assign x_4172 = v_4079 | ~v_101;
assign x_4173 = v_4079 | ~v_100;
assign x_4174 = v_4079 | ~v_98;
assign x_4175 = v_4079 | ~v_93;
assign x_4176 = v_4078 | ~v_1142;
assign x_4177 = v_4078 | ~v_1143;
assign x_4178 = v_4078 | ~v_3114;
assign x_4179 = v_4078 | ~v_3115;
assign x_4180 = v_4078 | ~v_960;
assign x_4181 = v_4078 | ~v_3116;
assign x_4182 = v_4078 | ~v_3117;
assign x_4183 = v_4078 | ~v_961;
assign x_4184 = v_4078 | ~v_2427;
assign x_4185 = v_4078 | ~v_2428;
assign x_4186 = v_4078 | ~v_2429;
assign x_4187 = v_4078 | ~v_2430;
assign x_4188 = v_4078 | ~v_3118;
assign x_4189 = v_4078 | ~v_3119;
assign x_4190 = v_4078 | ~v_3120;
assign x_4191 = v_4078 | ~v_806;
assign x_4192 = v_4078 | ~v_3121;
assign x_4193 = v_4078 | ~v_3122;
assign x_4194 = v_4078 | ~v_4050;
assign x_4195 = v_4078 | ~v_4051;
assign x_4196 = v_4078 | ~v_2431;
assign x_4197 = v_4078 | ~v_2432;
assign x_4198 = v_4078 | ~v_2433;
assign x_4199 = v_4078 | ~v_4052;
assign x_4200 = v_4078 | ~v_4053;
assign x_4201 = v_4078 | ~v_2434;
assign x_4202 = v_4078 | ~v_2435;
assign x_4203 = v_4078 | ~v_2436;
assign x_4204 = v_4078 | ~v_3123;
assign x_4205 = v_4078 | ~v_807;
assign x_4206 = v_4078 | ~v_1144;
assign x_4207 = v_4078 | ~v_1145;
assign x_4208 = v_4078 | ~v_183;
assign x_4209 = v_4078 | ~v_166;
assign x_4210 = v_4078 | ~v_145;
assign x_4211 = v_4078 | ~v_144;
assign x_4212 = v_4078 | ~v_143;
assign x_4213 = v_4078 | ~v_142;
assign x_4214 = v_4078 | ~v_61;
assign x_4215 = v_4078 | ~v_60;
assign x_4216 = v_4078 | ~v_59;
assign x_4217 = v_4078 | ~v_58;
assign x_4218 = v_4078 | ~v_56;
assign x_4219 = v_4078 | ~v_51;
assign x_4220 = v_4077 | ~v_1137;
assign x_4221 = v_4077 | ~v_1138;
assign x_4222 = v_4077 | ~v_3099;
assign x_4223 = v_4077 | ~v_3100;
assign x_4224 = v_4077 | ~v_945;
assign x_4225 = v_4077 | ~v_3101;
assign x_4226 = v_4077 | ~v_3102;
assign x_4227 = v_4077 | ~v_946;
assign x_4228 = v_4077 | ~v_2412;
assign x_4229 = v_4077 | ~v_2413;
assign x_4230 = v_4077 | ~v_2414;
assign x_4231 = v_4077 | ~v_2415;
assign x_4232 = v_4077 | ~v_3103;
assign x_4233 = v_4077 | ~v_3104;
assign x_4234 = v_4077 | ~v_773;
assign x_4235 = v_4077 | ~v_3105;
assign x_4236 = v_4077 | ~v_3106;
assign x_4237 = v_4077 | ~v_774;
assign x_4238 = v_4077 | ~v_4045;
assign x_4239 = v_4077 | ~v_4046;
assign x_4240 = v_4077 | ~v_2416;
assign x_4241 = v_4077 | ~v_2417;
assign x_4242 = v_4077 | ~v_2418;
assign x_4243 = v_4077 | ~v_4047;
assign x_4244 = v_4077 | ~v_4048;
assign x_4245 = v_4077 | ~v_2419;
assign x_4246 = v_4077 | ~v_2420;
assign x_4247 = v_4077 | ~v_2421;
assign x_4248 = v_4077 | ~v_1139;
assign x_4249 = v_4077 | ~v_1140;
assign x_4250 = v_4077 | ~v_182;
assign x_4251 = v_4077 | ~v_162;
assign x_4252 = v_4077 | ~v_137;
assign x_4253 = v_4077 | ~v_136;
assign x_4254 = v_4077 | ~v_135;
assign x_4255 = v_4077 | ~v_134;
assign x_4256 = v_4077 | ~v_3107;
assign x_4257 = v_4077 | ~v_3108;
assign x_4258 = v_4077 | ~v_18;
assign x_4259 = v_4077 | ~v_17;
assign x_4260 = v_4077 | ~v_16;
assign x_4261 = v_4077 | ~v_15;
assign x_4262 = v_4077 | ~v_13;
assign x_4263 = v_4077 | ~v_8;
assign x_4264 = ~v_4075 | ~v_4074 | ~v_4073 | v_4076;
assign x_4265 = v_4075 | ~v_3251;
assign x_4266 = v_4075 | ~v_3252;
assign x_4267 = v_4075 | ~v_885;
assign x_4268 = v_4075 | ~v_1019;
assign x_4269 = v_4075 | ~v_1020;
assign x_4270 = v_4075 | ~v_3253;
assign x_4271 = v_4075 | ~v_3254;
assign x_4272 = v_4075 | ~v_886;
assign x_4273 = v_4075 | ~v_1021;
assign x_4274 = v_4075 | ~v_1022;
assign x_4275 = v_4075 | ~v_2564;
assign x_4276 = v_4075 | ~v_2565;
assign x_4277 = v_4075 | ~v_2566;
assign x_4278 = v_4075 | ~v_2567;
assign x_4279 = v_4075 | ~v_3133;
assign x_4280 = v_4075 | ~v_3199;
assign x_4281 = v_4075 | ~v_3200;
assign x_4282 = v_4075 | ~v_1023;
assign x_4283 = v_4075 | ~v_3136;
assign x_4284 = v_4075 | ~v_3201;
assign x_4285 = v_4075 | ~v_3202;
assign x_4286 = v_4075 | ~v_1024;
assign x_4287 = v_4075 | ~v_4055;
assign x_4288 = v_4075 | ~v_4056;
assign x_4289 = v_4075 | ~v_2446;
assign x_4290 = v_4075 | ~v_2512;
assign x_4291 = v_4075 | ~v_2513;
assign x_4292 = v_4075 | ~v_4057;
assign x_4293 = v_4075 | ~v_4058;
assign x_4294 = v_4075 | ~v_2449;
assign x_4295 = v_4075 | ~v_2514;
assign x_4296 = v_4075 | ~v_2515;
assign x_4297 = v_4075 | ~v_184;
assign x_4298 = v_4075 | ~v_181;
assign x_4299 = v_4075 | ~v_171;
assign x_4300 = v_4075 | ~v_170;
assign x_4301 = v_4075 | ~v_169;
assign x_4302 = v_4075 | ~v_149;
assign x_4303 = v_4075 | ~v_147;
assign x_4304 = v_4075 | ~v_103;
assign x_4305 = v_4075 | ~v_102;
assign x_4306 = v_4075 | ~v_101;
assign x_4307 = v_4075 | ~v_99;
assign x_4308 = v_4075 | ~v_96;
assign x_4309 = v_4074 | ~v_3246;
assign x_4310 = v_4074 | ~v_3247;
assign x_4311 = v_4074 | ~v_870;
assign x_4312 = v_4074 | ~v_1004;
assign x_4313 = v_4074 | ~v_1005;
assign x_4314 = v_4074 | ~v_3248;
assign x_4315 = v_4074 | ~v_3249;
assign x_4316 = v_4074 | ~v_871;
assign x_4317 = v_4074 | ~v_1006;
assign x_4318 = v_4074 | ~v_1007;
assign x_4319 = v_4074 | ~v_2559;
assign x_4320 = v_4074 | ~v_2560;
assign x_4321 = v_4074 | ~v_2561;
assign x_4322 = v_4074 | ~v_2562;
assign x_4323 = v_4074 | ~v_3118;
assign x_4324 = v_4074 | ~v_3194;
assign x_4325 = v_4074 | ~v_3195;
assign x_4326 = v_4074 | ~v_1008;
assign x_4327 = v_4074 | ~v_3121;
assign x_4328 = v_4074 | ~v_1009;
assign x_4329 = v_4074 | ~v_4050;
assign x_4330 = v_4074 | ~v_4051;
assign x_4331 = v_4074 | ~v_2431;
assign x_4332 = v_4074 | ~v_2507;
assign x_4333 = v_4074 | ~v_2508;
assign x_4334 = v_4074 | ~v_4052;
assign x_4335 = v_4074 | ~v_4053;
assign x_4336 = v_4074 | ~v_2434;
assign x_4337 = v_4074 | ~v_2509;
assign x_4338 = v_4074 | ~v_2510;
assign x_4339 = v_4074 | ~v_3196;
assign x_4340 = v_4074 | ~v_183;
assign x_4341 = v_4074 | ~v_180;
assign x_4342 = v_4074 | ~v_167;
assign x_4343 = v_4074 | ~v_166;
assign x_4344 = v_4074 | ~v_165;
assign x_4345 = v_4074 | ~v_144;
assign x_4346 = v_4074 | ~v_142;
assign x_4347 = v_4074 | ~v_3197;
assign x_4348 = v_4074 | ~v_61;
assign x_4349 = v_4074 | ~v_60;
assign x_4350 = v_4074 | ~v_59;
assign x_4351 = v_4074 | ~v_57;
assign x_4352 = v_4074 | ~v_54;
assign x_4353 = v_4073 | ~v_3241;
assign x_4354 = v_4073 | ~v_3242;
assign x_4355 = v_4073 | ~v_855;
assign x_4356 = v_4073 | ~v_989;
assign x_4357 = v_4073 | ~v_990;
assign x_4358 = v_4073 | ~v_3243;
assign x_4359 = v_4073 | ~v_3244;
assign x_4360 = v_4073 | ~v_856;
assign x_4361 = v_4073 | ~v_991;
assign x_4362 = v_4073 | ~v_992;
assign x_4363 = v_4073 | ~v_2554;
assign x_4364 = v_4073 | ~v_2555;
assign x_4365 = v_4073 | ~v_2556;
assign x_4366 = v_4073 | ~v_2557;
assign x_4367 = v_4073 | ~v_3189;
assign x_4368 = v_4073 | ~v_3190;
assign x_4369 = v_4073 | ~v_3191;
assign x_4370 = v_4073 | ~v_3192;
assign x_4371 = v_4073 | ~v_4045;
assign x_4372 = v_4073 | ~v_4046;
assign x_4373 = v_4073 | ~v_2416;
assign x_4374 = v_4073 | ~v_2502;
assign x_4375 = v_4073 | ~v_2503;
assign x_4376 = v_4073 | ~v_4047;
assign x_4377 = v_4073 | ~v_4048;
assign x_4378 = v_4073 | ~v_2419;
assign x_4379 = v_4073 | ~v_2504;
assign x_4380 = v_4073 | ~v_2505;
assign x_4381 = v_4073 | ~v_182;
assign x_4382 = v_4073 | ~v_179;
assign x_4383 = v_4073 | ~v_163;
assign x_4384 = v_4073 | ~v_162;
assign x_4385 = v_4073 | ~v_161;
assign x_4386 = v_4073 | ~v_136;
assign x_4387 = v_4073 | ~v_134;
assign x_4388 = v_4073 | ~v_3107;
assign x_4389 = v_4073 | ~v_993;
assign x_4390 = v_4073 | ~v_3108;
assign x_4391 = v_4073 | ~v_994;
assign x_4392 = v_4073 | ~v_18;
assign x_4393 = v_4073 | ~v_17;
assign x_4394 = v_4073 | ~v_16;
assign x_4395 = v_4073 | ~v_14;
assign x_4396 = v_4073 | ~v_11;
assign x_4397 = ~v_4071 | ~v_4070 | ~v_4069 | v_4072;
assign x_4398 = v_4071 | ~v_925;
assign x_4399 = v_4071 | ~v_926;
assign x_4400 = v_4071 | ~v_3251;
assign x_4401 = v_4071 | ~v_3252;
assign x_4402 = v_4071 | ~v_885;
assign x_4403 = v_4071 | ~v_3253;
assign x_4404 = v_4071 | ~v_3254;
assign x_4405 = v_4071 | ~v_886;
assign x_4406 = v_4071 | ~v_2564;
assign x_4407 = v_4071 | ~v_2565;
assign x_4408 = v_4071 | ~v_2566;
assign x_4409 = v_4071 | ~v_2567;
assign x_4410 = v_4071 | ~v_3167;
assign x_4411 = v_4071 | ~v_3168;
assign x_4412 = v_4071 | ~v_927;
assign x_4413 = v_4071 | ~v_3169;
assign x_4414 = v_4071 | ~v_3170;
assign x_4415 = v_4071 | ~v_928;
assign x_4416 = v_4071 | ~v_2480;
assign x_4417 = v_4071 | ~v_2481;
assign x_4418 = v_4071 | ~v_2482;
assign x_4419 = v_4071 | ~v_2483;
assign x_4420 = v_4071 | ~v_3133;
assign x_4421 = v_4071 | ~v_3136;
assign x_4422 = v_4071 | ~v_4055;
assign x_4423 = v_4071 | ~v_4056;
assign x_4424 = v_4071 | ~v_2446;
assign x_4425 = v_4071 | ~v_4057;
assign x_4426 = v_4071 | ~v_4058;
assign x_4427 = v_4071 | ~v_2449;
assign x_4428 = v_4071 | ~v_929;
assign x_4429 = v_4071 | ~v_930;
assign x_4430 = v_4071 | ~v_184;
assign x_4431 = v_4071 | ~v_181;
assign x_4432 = v_4071 | ~v_171;
assign x_4433 = v_4071 | ~v_170;
assign x_4434 = v_4071 | ~v_169;
assign x_4435 = v_4071 | ~v_150;
assign x_4436 = v_4071 | ~v_148;
assign x_4437 = v_4071 | ~v_147;
assign x_4438 = v_4071 | ~v_103;
assign x_4439 = v_4071 | ~v_102;
assign x_4440 = v_4071 | ~v_101;
assign x_4441 = v_4071 | ~v_97;
assign x_4442 = v_4070 | ~v_910;
assign x_4443 = v_4070 | ~v_911;
assign x_4444 = v_4070 | ~v_3246;
assign x_4445 = v_4070 | ~v_3247;
assign x_4446 = v_4070 | ~v_870;
assign x_4447 = v_4070 | ~v_3248;
assign x_4448 = v_4070 | ~v_3249;
assign x_4449 = v_4070 | ~v_871;
assign x_4450 = v_4070 | ~v_2559;
assign x_4451 = v_4070 | ~v_2560;
assign x_4452 = v_4070 | ~v_2561;
assign x_4453 = v_4070 | ~v_2562;
assign x_4454 = v_4070 | ~v_3162;
assign x_4455 = v_4070 | ~v_3163;
assign x_4456 = v_4070 | ~v_912;
assign x_4457 = v_4070 | ~v_3164;
assign x_4458 = v_4070 | ~v_3165;
assign x_4459 = v_4070 | ~v_913;
assign x_4460 = v_4070 | ~v_2475;
assign x_4461 = v_4070 | ~v_2476;
assign x_4462 = v_4070 | ~v_2477;
assign x_4463 = v_4070 | ~v_2478;
assign x_4464 = v_4070 | ~v_3118;
assign x_4465 = v_4070 | ~v_3121;
assign x_4466 = v_4070 | ~v_4050;
assign x_4467 = v_4070 | ~v_4051;
assign x_4468 = v_4070 | ~v_2431;
assign x_4469 = v_4070 | ~v_4052;
assign x_4470 = v_4070 | ~v_4053;
assign x_4471 = v_4070 | ~v_2434;
assign x_4472 = v_4070 | ~v_914;
assign x_4473 = v_4070 | ~v_915;
assign x_4474 = v_4070 | ~v_183;
assign x_4475 = v_4070 | ~v_180;
assign x_4476 = v_4070 | ~v_167;
assign x_4477 = v_4070 | ~v_166;
assign x_4478 = v_4070 | ~v_165;
assign x_4479 = v_4070 | ~v_145;
assign x_4480 = v_4070 | ~v_143;
assign x_4481 = v_4070 | ~v_142;
assign x_4482 = v_4070 | ~v_61;
assign x_4483 = v_4070 | ~v_60;
assign x_4484 = v_4070 | ~v_59;
assign x_4485 = v_4070 | ~v_55;
assign x_4486 = v_4069 | ~v_895;
assign x_4487 = v_4069 | ~v_896;
assign x_4488 = v_4069 | ~v_3241;
assign x_4489 = v_4069 | ~v_3242;
assign x_4490 = v_4069 | ~v_855;
assign x_4491 = v_4069 | ~v_3243;
assign x_4492 = v_4069 | ~v_3244;
assign x_4493 = v_4069 | ~v_856;
assign x_4494 = v_4069 | ~v_2554;
assign x_4495 = v_4069 | ~v_2555;
assign x_4496 = v_4069 | ~v_2556;
assign x_4497 = v_4069 | ~v_2557;
assign x_4498 = v_4069 | ~v_3157;
assign x_4499 = v_4069 | ~v_3158;
assign x_4500 = v_4069 | ~v_897;
assign x_4501 = v_4069 | ~v_3159;
assign x_4502 = v_4069 | ~v_3160;
assign x_4503 = v_4069 | ~v_898;
assign x_4504 = v_4069 | ~v_2470;
assign x_4505 = v_4069 | ~v_2471;
assign x_4506 = v_4069 | ~v_2472;
assign x_4507 = v_4069 | ~v_2473;
assign x_4508 = v_4069 | ~v_4045;
assign x_4509 = v_4069 | ~v_4046;
assign x_4510 = v_4069 | ~v_2416;
assign x_4511 = v_4069 | ~v_4047;
assign x_4512 = v_4069 | ~v_4048;
assign x_4513 = v_4069 | ~v_2419;
assign x_4514 = v_4069 | ~v_899;
assign x_4515 = v_4069 | ~v_900;
assign x_4516 = v_4069 | ~v_182;
assign x_4517 = v_4069 | ~v_179;
assign x_4518 = v_4069 | ~v_163;
assign x_4519 = v_4069 | ~v_162;
assign x_4520 = v_4069 | ~v_161;
assign x_4521 = v_4069 | ~v_137;
assign x_4522 = v_4069 | ~v_135;
assign x_4523 = v_4069 | ~v_134;
assign x_4524 = v_4069 | ~v_3107;
assign x_4525 = v_4069 | ~v_3108;
assign x_4526 = v_4069 | ~v_18;
assign x_4527 = v_4069 | ~v_17;
assign x_4528 = v_4069 | ~v_16;
assign x_4529 = v_4069 | ~v_12;
assign x_4530 = ~v_4067 | ~v_4066 | ~v_4065 | v_4068;
assign x_4531 = v_4067 | ~v_973;
assign x_4532 = v_4067 | ~v_974;
assign x_4533 = v_4067 | ~v_3251;
assign x_4534 = v_4067 | ~v_3252;
assign x_4535 = v_4067 | ~v_885;
assign x_4536 = v_4067 | ~v_3253;
assign x_4537 = v_4067 | ~v_3254;
assign x_4538 = v_4067 | ~v_886;
assign x_4539 = v_4067 | ~v_2564;
assign x_4540 = v_4067 | ~v_2565;
assign x_4541 = v_4067 | ~v_2566;
assign x_4542 = v_4067 | ~v_2567;
assign x_4543 = v_4067 | ~v_3129;
assign x_4544 = v_4067 | ~v_3130;
assign x_4545 = v_4067 | ~v_975;
assign x_4546 = v_4067 | ~v_3131;
assign x_4547 = v_4067 | ~v_3132;
assign x_4548 = v_4067 | ~v_976;
assign x_4549 = v_4067 | ~v_2442;
assign x_4550 = v_4067 | ~v_2443;
assign x_4551 = v_4067 | ~v_2444;
assign x_4552 = v_4067 | ~v_2445;
assign x_4553 = v_4067 | ~v_3133;
assign x_4554 = v_4067 | ~v_3136;
assign x_4555 = v_4067 | ~v_4055;
assign x_4556 = v_4067 | ~v_4056;
assign x_4557 = v_4067 | ~v_2446;
assign x_4558 = v_4067 | ~v_4057;
assign x_4559 = v_4067 | ~v_4058;
assign x_4560 = v_4067 | ~v_2449;
assign x_4561 = v_4067 | ~v_977;
assign x_4562 = v_4067 | ~v_978;
assign x_4563 = v_4067 | ~v_184;
assign x_4564 = v_4067 | ~v_181;
assign x_4565 = v_4067 | ~v_172;
assign x_4566 = v_4067 | ~v_171;
assign x_4567 = v_4067 | ~v_170;
assign x_4568 = v_4067 | ~v_169;
assign x_4569 = v_4067 | ~v_150;
assign x_4570 = v_4067 | ~v_149;
assign x_4571 = v_4067 | ~v_148;
assign x_4572 = v_4067 | ~v_147;
assign x_4573 = v_4067 | ~v_102;
assign x_4574 = v_4067 | ~v_101;
assign x_4575 = v_4066 | ~v_958;
assign x_4576 = v_4066 | ~v_959;
assign x_4577 = v_4066 | ~v_3246;
assign x_4578 = v_4066 | ~v_3247;
assign x_4579 = v_4066 | ~v_870;
assign x_4580 = v_4066 | ~v_3248;
assign x_4581 = v_4066 | ~v_3249;
assign x_4582 = v_4066 | ~v_871;
assign x_4583 = v_4066 | ~v_2559;
assign x_4584 = v_4066 | ~v_2560;
assign x_4585 = v_4066 | ~v_2561;
assign x_4586 = v_4066 | ~v_2562;
assign x_4587 = v_4066 | ~v_3114;
assign x_4588 = v_4066 | ~v_3115;
assign x_4589 = v_4066 | ~v_960;
assign x_4590 = v_4066 | ~v_3116;
assign x_4591 = v_4066 | ~v_3117;
assign x_4592 = v_4066 | ~v_961;
assign x_4593 = v_4066 | ~v_2427;
assign x_4594 = v_4066 | ~v_2428;
assign x_4595 = v_4066 | ~v_2429;
assign x_4596 = v_4066 | ~v_2430;
assign x_4597 = v_4066 | ~v_3118;
assign x_4598 = v_4066 | ~v_3121;
assign x_4599 = v_4066 | ~v_4050;
assign x_4600 = v_4066 | ~v_4051;
assign x_4601 = v_4066 | ~v_2431;
assign x_4602 = v_4066 | ~v_4052;
assign x_4603 = v_4066 | ~v_4053;
assign x_4604 = v_4066 | ~v_2434;
assign x_4605 = v_4066 | ~v_962;
assign x_4606 = v_4066 | ~v_963;
assign x_4607 = v_4066 | ~v_183;
assign x_4608 = v_4066 | ~v_180;
assign x_4609 = v_4066 | ~v_168;
assign x_4610 = v_4066 | ~v_167;
assign x_4611 = v_4066 | ~v_166;
assign x_4612 = v_4066 | ~v_165;
assign x_4613 = v_4066 | ~v_145;
assign x_4614 = v_4066 | ~v_144;
assign x_4615 = v_4066 | ~v_143;
assign x_4616 = v_4066 | ~v_142;
assign x_4617 = v_4066 | ~v_60;
assign x_4618 = v_4066 | ~v_59;
assign x_4619 = v_4065 | ~v_943;
assign x_4620 = v_4065 | ~v_944;
assign x_4621 = v_4065 | ~v_3241;
assign x_4622 = v_4065 | ~v_3242;
assign x_4623 = v_4065 | ~v_855;
assign x_4624 = v_4065 | ~v_3243;
assign x_4625 = v_4065 | ~v_3244;
assign x_4626 = v_4065 | ~v_856;
assign x_4627 = v_4065 | ~v_2554;
assign x_4628 = v_4065 | ~v_2555;
assign x_4629 = v_4065 | ~v_2556;
assign x_4630 = v_4065 | ~v_2557;
assign x_4631 = v_4065 | ~v_3099;
assign x_4632 = v_4065 | ~v_3100;
assign x_4633 = v_4065 | ~v_945;
assign x_4634 = v_4065 | ~v_3101;
assign x_4635 = v_4065 | ~v_3102;
assign x_4636 = v_4065 | ~v_946;
assign x_4637 = v_4065 | ~v_2412;
assign x_4638 = v_4065 | ~v_2413;
assign x_4639 = v_4065 | ~v_2414;
assign x_4640 = v_4065 | ~v_2415;
assign x_4641 = v_4065 | ~v_4045;
assign x_4642 = v_4065 | ~v_4046;
assign x_4643 = v_4065 | ~v_2416;
assign x_4644 = v_4065 | ~v_4047;
assign x_4645 = v_4065 | ~v_4048;
assign x_4646 = v_4065 | ~v_2419;
assign x_4647 = v_4065 | ~v_947;
assign x_4648 = v_4065 | ~v_948;
assign x_4649 = v_4065 | ~v_182;
assign x_4650 = v_4065 | ~v_179;
assign x_4651 = v_4065 | ~v_164;
assign x_4652 = v_4065 | ~v_163;
assign x_4653 = v_4065 | ~v_162;
assign x_4654 = v_4065 | ~v_161;
assign x_4655 = v_4065 | ~v_137;
assign x_4656 = v_4065 | ~v_136;
assign x_4657 = v_4065 | ~v_135;
assign x_4658 = v_4065 | ~v_134;
assign x_4659 = v_4065 | ~v_3107;
assign x_4660 = v_4065 | ~v_3108;
assign x_4661 = v_4065 | ~v_17;
assign x_4662 = v_4065 | ~v_16;
assign x_4663 = ~v_4063 | ~v_4062 | ~v_4061 | v_4064;
assign x_4664 = v_4063 | ~v_881;
assign x_4665 = v_4063 | ~v_882;
assign x_4666 = v_4063 | ~v_883;
assign x_4667 = v_4063 | ~v_884;
assign x_4668 = v_4063 | ~v_3251;
assign x_4669 = v_4063 | ~v_3252;
assign x_4670 = v_4063 | ~v_885;
assign x_4671 = v_4063 | ~v_3253;
assign x_4672 = v_4063 | ~v_3254;
assign x_4673 = v_4063 | ~v_886;
assign x_4674 = v_4063 | ~v_2564;
assign x_4675 = v_4063 | ~v_2565;
assign x_4676 = v_4063 | ~v_2566;
assign x_4677 = v_4063 | ~v_2567;
assign x_4678 = v_4063 | ~v_3183;
assign x_4679 = v_4063 | ~v_3184;
assign x_4680 = v_4063 | ~v_837;
assign x_4681 = v_4063 | ~v_3185;
assign x_4682 = v_4063 | ~v_3186;
assign x_4683 = v_4063 | ~v_838;
assign x_4684 = v_4063 | ~v_2496;
assign x_4685 = v_4063 | ~v_2497;
assign x_4686 = v_4063 | ~v_2498;
assign x_4687 = v_4063 | ~v_2499;
assign x_4688 = v_4063 | ~v_3133;
assign x_4689 = v_4063 | ~v_3136;
assign x_4690 = v_4063 | ~v_4055;
assign x_4691 = v_4063 | ~v_4056;
assign x_4692 = v_4063 | ~v_2446;
assign x_4693 = v_4063 | ~v_4057;
assign x_4694 = v_4063 | ~v_4058;
assign x_4695 = v_4063 | ~v_2449;
assign x_4696 = v_4063 | ~v_184;
assign x_4697 = v_4063 | ~v_181;
assign x_4698 = v_4063 | ~v_171;
assign x_4699 = v_4063 | ~v_170;
assign x_4700 = v_4063 | ~v_169;
assign x_4701 = v_4063 | ~v_160;
assign x_4702 = v_4063 | ~v_150;
assign x_4703 = v_4063 | ~v_149;
assign x_4704 = v_4063 | ~v_148;
assign x_4705 = v_4063 | ~v_103;
assign x_4706 = v_4063 | ~v_102;
assign x_4707 = v_4063 | ~v_95;
assign x_4708 = v_4062 | ~v_866;
assign x_4709 = v_4062 | ~v_867;
assign x_4710 = v_4062 | ~v_868;
assign x_4711 = v_4062 | ~v_869;
assign x_4712 = v_4062 | ~v_3246;
assign x_4713 = v_4062 | ~v_3247;
assign x_4714 = v_4062 | ~v_870;
assign x_4715 = v_4062 | ~v_3248;
assign x_4716 = v_4062 | ~v_3249;
assign x_4717 = v_4062 | ~v_871;
assign x_4718 = v_4062 | ~v_2559;
assign x_4719 = v_4062 | ~v_2560;
assign x_4720 = v_4062 | ~v_2561;
assign x_4721 = v_4062 | ~v_2562;
assign x_4722 = v_4062 | ~v_3178;
assign x_4723 = v_4062 | ~v_3179;
assign x_4724 = v_4062 | ~v_804;
assign x_4725 = v_4062 | ~v_3180;
assign x_4726 = v_4062 | ~v_3181;
assign x_4727 = v_4062 | ~v_805;
assign x_4728 = v_4062 | ~v_2491;
assign x_4729 = v_4062 | ~v_2492;
assign x_4730 = v_4062 | ~v_2493;
assign x_4731 = v_4062 | ~v_2494;
assign x_4732 = v_4062 | ~v_3118;
assign x_4733 = v_4062 | ~v_3121;
assign x_4734 = v_4062 | ~v_4050;
assign x_4735 = v_4062 | ~v_4051;
assign x_4736 = v_4062 | ~v_2431;
assign x_4737 = v_4062 | ~v_4052;
assign x_4738 = v_4062 | ~v_4053;
assign x_4739 = v_4062 | ~v_2434;
assign x_4740 = v_4062 | ~v_183;
assign x_4741 = v_4062 | ~v_180;
assign x_4742 = v_4062 | ~v_167;
assign x_4743 = v_4062 | ~v_166;
assign x_4744 = v_4062 | ~v_165;
assign x_4745 = v_4062 | ~v_159;
assign x_4746 = v_4062 | ~v_145;
assign x_4747 = v_4062 | ~v_144;
assign x_4748 = v_4062 | ~v_143;
assign x_4749 = v_4062 | ~v_61;
assign x_4750 = v_4062 | ~v_60;
assign x_4751 = v_4062 | ~v_53;
assign x_4752 = v_4061 | ~v_851;
assign x_4753 = v_4061 | ~v_852;
assign x_4754 = v_4061 | ~v_853;
assign x_4755 = v_4061 | ~v_854;
assign x_4756 = v_4061 | ~v_3241;
assign x_4757 = v_4061 | ~v_3242;
assign x_4758 = v_4061 | ~v_855;
assign x_4759 = v_4061 | ~v_3243;
assign x_4760 = v_4061 | ~v_3244;
assign x_4761 = v_4061 | ~v_856;
assign x_4762 = v_4061 | ~v_2554;
assign x_4763 = v_4061 | ~v_2555;
assign x_4764 = v_4061 | ~v_2556;
assign x_4765 = v_4061 | ~v_2557;
assign x_4766 = v_4061 | ~v_3173;
assign x_4767 = v_4061 | ~v_3174;
assign x_4768 = v_4061 | ~v_771;
assign x_4769 = v_4061 | ~v_3175;
assign x_4770 = v_4061 | ~v_3176;
assign x_4771 = v_4061 | ~v_772;
assign x_4772 = v_4061 | ~v_2486;
assign x_4773 = v_4061 | ~v_2487;
assign x_4774 = v_4061 | ~v_2488;
assign x_4775 = v_4061 | ~v_2489;
assign x_4776 = v_4061 | ~v_4045;
assign x_4777 = v_4061 | ~v_4046;
assign x_4778 = v_4061 | ~v_2416;
assign x_4779 = v_4061 | ~v_4047;
assign x_4780 = v_4061 | ~v_4048;
assign x_4781 = v_4061 | ~v_2419;
assign x_4782 = v_4061 | ~v_182;
assign x_4783 = v_4061 | ~v_179;
assign x_4784 = v_4061 | ~v_163;
assign x_4785 = v_4061 | ~v_162;
assign x_4786 = v_4061 | ~v_161;
assign x_4787 = v_4061 | ~v_155;
assign x_4788 = v_4061 | ~v_137;
assign x_4789 = v_4061 | ~v_136;
assign x_4790 = v_4061 | ~v_135;
assign x_4791 = v_4061 | ~v_3107;
assign x_4792 = v_4061 | ~v_3108;
assign x_4793 = v_4061 | ~v_18;
assign x_4794 = v_4061 | ~v_17;
assign x_4795 = v_4061 | ~v_10;
assign x_4796 = ~v_4059 | ~v_4054 | ~v_4049 | v_4060;
assign x_4797 = v_4059 | ~v_833;
assign x_4798 = v_4059 | ~v_834;
assign x_4799 = v_4059 | ~v_835;
assign x_4800 = v_4059 | ~v_836;
assign x_4801 = v_4059 | ~v_3183;
assign x_4802 = v_4059 | ~v_3184;
assign x_4803 = v_4059 | ~v_837;
assign x_4804 = v_4059 | ~v_3185;
assign x_4805 = v_4059 | ~v_3186;
assign x_4806 = v_4059 | ~v_838;
assign x_4807 = v_4059 | ~v_2496;
assign x_4808 = v_4059 | ~v_2497;
assign x_4809 = v_4059 | ~v_2498;
assign x_4810 = v_4059 | ~v_2499;
assign x_4811 = v_4059 | ~v_3133;
assign x_4812 = v_4059 | ~v_3134;
assign x_4813 = v_4059 | ~v_3135;
assign x_4814 = v_4059 | ~v_839;
assign x_4815 = v_4059 | ~v_3136;
assign x_4816 = v_4059 | ~v_3137;
assign x_4817 = v_4059 | ~v_3138;
assign x_4818 = v_4059 | ~v_840;
assign x_4819 = v_4059 | ~v_4055;
assign x_4820 = v_4059 | ~v_4056;
assign x_4821 = v_4059 | ~v_2446;
assign x_4822 = v_4059 | ~v_2447;
assign x_4823 = v_4059 | ~v_2448;
assign x_4824 = v_4059 | ~v_4057;
assign x_4825 = v_4059 | ~v_4058;
assign x_4826 = v_4059 | ~v_2449;
assign x_4827 = v_4059 | ~v_2450;
assign x_4828 = v_4059 | ~v_2451;
assign x_4829 = v_4059 | ~v_184;
assign x_4830 = v_4059 | ~v_170;
assign x_4831 = v_4059 | ~v_160;
assign x_4832 = v_4059 | ~v_150;
assign x_4833 = v_4059 | ~v_149;
assign x_4834 = v_4059 | ~v_148;
assign x_4835 = v_4059 | ~v_147;
assign x_4836 = v_4059 | ~v_103;
assign x_4837 = v_4059 | ~v_102;
assign x_4838 = v_4059 | ~v_100;
assign x_4839 = v_4059 | ~v_98;
assign x_4840 = v_4059 | ~v_93;
assign x_4841 = ~v_123 | ~v_140 | v_4058;
assign x_4842 = ~v_120 | ~v_139 | v_4057;
assign x_4843 = ~v_108 | v_140 | v_4056;
assign x_4844 = ~v_105 | v_139 | v_4055;
assign x_4845 = v_4054 | ~v_800;
assign x_4846 = v_4054 | ~v_801;
assign x_4847 = v_4054 | ~v_802;
assign x_4848 = v_4054 | ~v_803;
assign x_4849 = v_4054 | ~v_3178;
assign x_4850 = v_4054 | ~v_3179;
assign x_4851 = v_4054 | ~v_804;
assign x_4852 = v_4054 | ~v_3180;
assign x_4853 = v_4054 | ~v_3181;
assign x_4854 = v_4054 | ~v_805;
assign x_4855 = v_4054 | ~v_2491;
assign x_4856 = v_4054 | ~v_2492;
assign x_4857 = v_4054 | ~v_2493;
assign x_4858 = v_4054 | ~v_2494;
assign x_4859 = v_4054 | ~v_3118;
assign x_4860 = v_4054 | ~v_3119;
assign x_4861 = v_4054 | ~v_3120;
assign x_4862 = v_4054 | ~v_806;
assign x_4863 = v_4054 | ~v_3121;
assign x_4864 = v_4054 | ~v_3122;
assign x_4865 = v_4054 | ~v_4050;
assign x_4866 = v_4054 | ~v_4051;
assign x_4867 = v_4054 | ~v_2431;
assign x_4868 = v_4054 | ~v_2432;
assign x_4869 = v_4054 | ~v_2433;
assign x_4870 = v_4054 | ~v_4052;
assign x_4871 = v_4054 | ~v_4053;
assign x_4872 = v_4054 | ~v_2434;
assign x_4873 = v_4054 | ~v_2435;
assign x_4874 = v_4054 | ~v_2436;
assign x_4875 = v_4054 | ~v_3123;
assign x_4876 = v_4054 | ~v_807;
assign x_4877 = v_4054 | ~v_183;
assign x_4878 = v_4054 | ~v_166;
assign x_4879 = v_4054 | ~v_159;
assign x_4880 = v_4054 | ~v_145;
assign x_4881 = v_4054 | ~v_144;
assign x_4882 = v_4054 | ~v_143;
assign x_4883 = v_4054 | ~v_142;
assign x_4884 = v_4054 | ~v_61;
assign x_4885 = v_4054 | ~v_60;
assign x_4886 = v_4054 | ~v_58;
assign x_4887 = v_4054 | ~v_56;
assign x_4888 = v_4054 | ~v_51;
assign x_4889 = ~v_81 | ~v_140 | v_4053;
assign x_4890 = ~v_78 | ~v_139 | v_4052;
assign x_4891 = ~v_66 | v_140 | v_4051;
assign x_4892 = ~v_63 | v_139 | v_4050;
assign x_4893 = v_4049 | ~v_767;
assign x_4894 = v_4049 | ~v_768;
assign x_4895 = v_4049 | ~v_769;
assign x_4896 = v_4049 | ~v_770;
assign x_4897 = v_4049 | ~v_3173;
assign x_4898 = v_4049 | ~v_3174;
assign x_4899 = v_4049 | ~v_771;
assign x_4900 = v_4049 | ~v_3175;
assign x_4901 = v_4049 | ~v_3176;
assign x_4902 = v_4049 | ~v_772;
assign x_4903 = v_4049 | ~v_2486;
assign x_4904 = v_4049 | ~v_2487;
assign x_4905 = v_4049 | ~v_2488;
assign x_4906 = v_4049 | ~v_2489;
assign x_4907 = v_4049 | ~v_3103;
assign x_4908 = v_4049 | ~v_3104;
assign x_4909 = v_4049 | ~v_773;
assign x_4910 = v_4049 | ~v_3105;
assign x_4911 = v_4049 | ~v_3106;
assign x_4912 = v_4049 | ~v_774;
assign x_4913 = v_4049 | ~v_4045;
assign x_4914 = v_4049 | ~v_4046;
assign x_4915 = v_4049 | ~v_2416;
assign x_4916 = v_4049 | ~v_2417;
assign x_4917 = v_4049 | ~v_2418;
assign x_4918 = v_4049 | ~v_4047;
assign x_4919 = v_4049 | ~v_4048;
assign x_4920 = v_4049 | ~v_2419;
assign x_4921 = v_4049 | ~v_2420;
assign x_4922 = v_4049 | ~v_2421;
assign x_4923 = v_4049 | ~v_182;
assign x_4924 = v_4049 | ~v_162;
assign x_4925 = v_4049 | ~v_155;
assign x_4926 = v_4049 | ~v_137;
assign x_4927 = v_4049 | ~v_136;
assign x_4928 = v_4049 | ~v_135;
assign x_4929 = v_4049 | ~v_134;
assign x_4930 = v_4049 | ~v_3107;
assign x_4931 = v_4049 | ~v_3108;
assign x_4932 = v_4049 | ~v_18;
assign x_4933 = v_4049 | ~v_17;
assign x_4934 = v_4049 | ~v_15;
assign x_4935 = v_4049 | ~v_13;
assign x_4936 = v_4049 | ~v_8;
assign x_4937 = ~v_39 | ~v_140 | v_4048;
assign x_4938 = ~v_36 | ~v_139 | v_4047;
assign x_4939 = ~v_24 | v_140 | v_4046;
assign x_4940 = ~v_21 | v_139 | v_4045;
assign x_4941 = v_4044 | ~v_1562;
assign x_4942 = v_4044 | ~v_737;
assign x_4943 = v_4043 | ~v_733;
assign x_4944 = v_4043 | ~v_727;
assign x_4945 = ~v_725 | ~v_724 | ~v_723 | ~v_722 | ~v_4041 | ~v_4037 | ~v_4033 | ~v_4029 | ~v_4025 | ~v_4021 | ~v_4017 | ~v_4013 | ~v_4009 | ~v_4005 | ~v_4001 | ~v_3997 | ~v_3993 | ~v_3989 | ~v_3985 | ~v_3981 | ~v_3965 | v_4042;
assign x_4946 = v_4041 | ~v_4038;
assign x_4947 = v_4041 | ~v_4039;
assign x_4948 = v_4041 | ~v_4040;
assign x_4949 = v_98 | v_103 | v_101 | v_96 | v_100 | v_95 | v_99 | v_93 | v_102 | ~v_719 | ~v_718 | v_170 | v_149 | v_184 | ~v_2331 | ~v_2267 | ~v_2330 | ~v_2266 | ~v_2265 | ~v_3979 | ~v_3978 | ~v_2329 | ~v_2264 | ~v_2328 | ~v_2263 | ~v_2262 | ~v_3977 | ~v_3976 | ~v_483 | ~v_717 | ~v_3021 | ~v_299 | ~v_2957 | ~v_3020 | ~v_2956 | ~v_2955 | ~v_482 | ~v_716 | ~v_3019 | ~v_298 | ~v_2954 | ~v_3018 | ~v_2953 | ~v_2952 | v_4040;
assign x_4950 = v_54 | v_53 | v_56 | v_61 | v_51 | v_60 | v_59 | v_58 | v_57 | ~v_714 | ~v_713 | ~v_3016 | v_144 | v_166 | v_183 | ~v_3015 | ~v_266 | ~v_2942 | ~v_2326 | ~v_2252 | ~v_2325 | ~v_2251 | ~v_2250 | ~v_3974 | ~v_3973 | ~v_2324 | ~v_2249 | ~v_2323 | ~v_2248 | ~v_2247 | ~v_3972 | ~v_3971 | ~v_468 | ~v_712 | ~v_2941 | ~v_2940 | ~v_467 | ~v_711 | ~v_3014 | ~v_265 | ~v_2939 | ~v_3013 | ~v_2938 | ~v_2937 | v_4039;
assign x_4951 = v_13 | v_18 | v_17 | v_16 | v_8 | v_15 | v_14 | v_11 | v_10 | ~v_453 | ~v_709 | ~v_2927 | ~v_452 | ~v_708 | ~v_2926 | v_136 | ~v_707 | ~v_706 | v_162 | v_182 | ~v_2321 | ~v_2237 | ~v_2320 | ~v_2236 | ~v_2235 | ~v_3969 | ~v_3968 | ~v_2319 | ~v_2234 | ~v_2318 | ~v_2233 | ~v_2232 | ~v_3967 | ~v_3966 | ~v_3011 | ~v_233 | ~v_2925 | ~v_3010 | ~v_2924 | ~v_3009 | ~v_232 | ~v_2923 | ~v_3008 | ~v_2922 | v_4038;
assign x_4952 = v_4037 | ~v_4034;
assign x_4953 = v_4037 | ~v_4035;
assign x_4954 = v_4037 | ~v_4036;
assign x_4955 = v_101 | v_96 | v_100 | v_94 | v_99 | v_102 | v_172 | v_171 | v_169 | v_149 | v_147 | v_184 | ~v_2331 | ~v_2330 | ~v_2265 | ~v_3979 | ~v_3978 | ~v_2329 | ~v_2328 | ~v_2262 | ~v_3977 | ~v_3976 | ~v_483 | ~v_3021 | ~v_3020 | ~v_2955 | ~v_482 | ~v_3019 | ~v_3018 | ~v_2952 | ~v_2351 | ~v_2350 | ~v_2349 | ~v_2348 | ~v_593 | ~v_592 | ~v_545 | ~v_3041 | ~v_3040 | ~v_591 | ~v_590 | ~v_544 | ~v_3039 | ~v_3038 | v_4036;
assign x_4956 = v_54 | v_52 | v_60 | v_59 | v_58 | v_57 | ~v_3016 | v_144 | v_142 | v_168 | v_167 | v_165 | v_183 | ~v_3015 | ~v_2326 | ~v_2325 | ~v_2250 | ~v_3974 | ~v_3973 | ~v_2324 | ~v_2323 | ~v_2247 | ~v_3972 | ~v_3971 | ~v_468 | ~v_2940 | ~v_467 | ~v_3014 | ~v_3013 | ~v_2937 | ~v_2346 | ~v_2345 | ~v_2344 | ~v_2343 | ~v_588 | ~v_587 | ~v_530 | ~v_3036 | ~v_3035 | ~v_586 | ~v_585 | ~v_529 | ~v_3034 | ~v_3033 | v_4035;
assign x_4957 = v_9 | v_17 | v_16 | v_15 | v_14 | v_11 | ~v_453 | ~v_2927 | ~v_452 | ~v_2926 | v_136 | v_134 | v_164 | v_163 | v_161 | v_182 | ~v_2321 | ~v_2320 | ~v_2235 | ~v_3969 | ~v_3968 | ~v_2319 | ~v_2318 | ~v_2232 | ~v_3967 | ~v_3966 | ~v_3011 | ~v_3010 | ~v_3009 | ~v_3008 | ~v_2341 | ~v_2340 | ~v_2339 | ~v_2338 | ~v_583 | ~v_582 | ~v_515 | ~v_3031 | ~v_3030 | ~v_581 | ~v_580 | ~v_514 | ~v_3029 | ~v_3028 | v_4034;
assign x_4958 = v_4033 | ~v_4030;
assign x_4959 = v_4033 | ~v_4031;
assign x_4960 = v_4033 | ~v_4032;
assign x_4961 = v_103 | v_101 | v_97 | v_100 | v_95 | v_94 | v_102 | v_171 | v_169 | v_150 | v_148 | v_184 | ~v_2265 | ~v_3979 | ~v_3978 | ~v_2262 | ~v_3977 | ~v_3976 | ~v_2955 | ~v_2952 | ~v_2351 | ~v_2350 | ~v_2349 | ~v_2348 | ~v_545 | ~v_3041 | ~v_3040 | ~v_544 | ~v_3039 | ~v_3038 | ~v_2299 | ~v_2298 | ~v_2297 | ~v_2296 | ~v_561 | ~v_560 | ~v_559 | ~v_558 | ~v_387 | ~v_2989 | ~v_2988 | ~v_386 | ~v_2987 | ~v_2986 | v_4032;
assign x_4962 = v_53 | v_55 | v_61 | v_52 | v_60 | v_59 | v_58 | v_145 | v_143 | v_167 | v_165 | v_183 | ~v_2250 | ~v_3974 | ~v_3973 | ~v_2247 | ~v_3972 | ~v_3971 | ~v_2940 | ~v_2937 | ~v_2346 | ~v_2345 | ~v_2344 | ~v_2343 | ~v_530 | ~v_3036 | ~v_3035 | ~v_529 | ~v_3034 | ~v_3033 | ~v_2294 | ~v_2293 | ~v_2292 | ~v_2291 | ~v_556 | ~v_555 | ~v_554 | ~v_553 | ~v_372 | ~v_2984 | ~v_2983 | ~v_371 | ~v_2982 | ~v_2981 | v_4031;
assign x_4963 = v_9 | v_18 | v_17 | v_16 | v_15 | v_12 | v_10 | ~v_2927 | ~v_2926 | v_135 | v_137 | v_163 | v_161 | v_182 | ~v_2235 | ~v_3969 | ~v_3968 | ~v_2232 | ~v_3967 | ~v_3966 | ~v_2341 | ~v_2340 | ~v_2339 | ~v_2338 | ~v_515 | ~v_3031 | ~v_3030 | ~v_514 | ~v_3029 | ~v_3028 | ~v_2289 | ~v_2288 | ~v_2287 | ~v_2286 | ~v_551 | ~v_550 | ~v_549 | ~v_548 | ~v_357 | ~v_2979 | ~v_2978 | ~v_356 | ~v_2977 | ~v_2976 | v_4030;
assign x_4964 = v_4029 | ~v_4026;
assign x_4965 = v_4029 | ~v_4027;
assign x_4966 = v_4029 | ~v_4028;
assign x_4967 = v_103 | v_101 | v_100 | v_94 | v_151 | v_171 | v_169 | v_150 | v_149 | v_148 | v_147 | v_184 | ~v_577 | ~v_576 | ~v_2265 | ~v_3979 | ~v_3978 | ~v_2262 | ~v_3977 | ~v_3976 | ~v_2955 | ~v_2952 | ~v_2351 | ~v_2350 | ~v_2349 | ~v_2348 | ~v_545 | ~v_3041 | ~v_3040 | ~v_544 | ~v_3039 | ~v_3038 | ~v_2261 | ~v_2260 | ~v_2259 | ~v_2258 | ~v_575 | ~v_574 | ~v_435 | ~v_2951 | ~v_2950 | ~v_434 | ~v_2949 | ~v_2948 | v_4028;
assign x_4968 = v_61 | v_52 | v_59 | v_58 | v_144 | v_145 | v_143 | v_142 | v_167 | v_165 | v_146 | v_183 | ~v_572 | ~v_571 | ~v_2250 | ~v_3974 | ~v_3973 | ~v_2247 | ~v_3972 | ~v_3971 | ~v_2940 | ~v_2937 | ~v_2346 | ~v_2345 | ~v_2344 | ~v_2343 | ~v_530 | ~v_3036 | ~v_3035 | ~v_529 | ~v_3034 | ~v_3033 | ~v_2246 | ~v_2245 | ~v_2244 | ~v_2243 | ~v_570 | ~v_569 | ~v_420 | ~v_2936 | ~v_2935 | ~v_419 | ~v_2934 | ~v_2933 | v_4027;
assign x_4969 = v_9 | v_18 | v_16 | v_15 | ~v_2927 | ~v_2926 | v_136 | v_135 | v_134 | v_137 | v_138 | v_163 | v_161 | v_182 | ~v_567 | ~v_566 | ~v_2235 | ~v_3969 | ~v_3968 | ~v_2232 | ~v_3967 | ~v_3966 | ~v_2341 | ~v_2340 | ~v_2339 | ~v_2338 | ~v_515 | ~v_3031 | ~v_3030 | ~v_514 | ~v_3029 | ~v_3028 | ~v_2231 | ~v_2230 | ~v_2229 | ~v_2228 | ~v_565 | ~v_564 | ~v_405 | ~v_2921 | ~v_2920 | ~v_404 | ~v_2919 | ~v_2918 | v_4026;
assign x_4970 = v_4025 | ~v_4022;
assign x_4971 = v_4025 | ~v_4023;
assign x_4972 = v_4025 | ~v_4024;
assign x_4973 = v_103 | v_100 | v_94 | v_102 | v_171 | v_169 | v_160 | v_150 | v_149 | v_148 | v_147 | v_184 | ~v_2265 | ~v_3979 | ~v_3978 | ~v_2262 | ~v_3977 | ~v_3976 | ~v_2955 | ~v_2952 | ~v_2351 | ~v_2350 | ~v_2349 | ~v_2348 | ~v_545 | ~v_3041 | ~v_3040 | ~v_544 | ~v_3039 | ~v_3038 | ~v_2315 | ~v_2314 | ~v_2313 | ~v_2312 | ~v_543 | ~v_542 | ~v_541 | ~v_540 | ~v_297 | ~v_3005 | ~v_3004 | ~v_296 | ~v_3003 | ~v_3002 | v_4024;
assign x_4974 = v_61 | v_52 | v_60 | v_58 | v_144 | v_159 | v_145 | v_143 | v_142 | v_167 | v_165 | v_183 | ~v_2250 | ~v_3974 | ~v_3973 | ~v_2247 | ~v_3972 | ~v_3971 | ~v_2940 | ~v_2937 | ~v_2346 | ~v_2345 | ~v_2344 | ~v_2343 | ~v_530 | ~v_3036 | ~v_3035 | ~v_529 | ~v_3034 | ~v_3033 | ~v_2310 | ~v_2309 | ~v_2308 | ~v_2307 | ~v_528 | ~v_527 | ~v_526 | ~v_525 | ~v_264 | ~v_3000 | ~v_2999 | ~v_263 | ~v_2998 | ~v_2997 | v_4023;
assign x_4975 = v_9 | v_18 | v_17 | v_15 | ~v_2927 | ~v_2926 | v_136 | v_135 | v_134 | v_137 | v_163 | v_161 | v_155 | v_182 | ~v_2235 | ~v_3969 | ~v_3968 | ~v_2232 | ~v_3967 | ~v_3966 | ~v_2341 | ~v_2340 | ~v_2339 | ~v_2338 | ~v_515 | ~v_3031 | ~v_3030 | ~v_514 | ~v_3029 | ~v_3028 | ~v_2305 | ~v_2304 | ~v_2303 | ~v_2302 | ~v_513 | ~v_512 | ~v_511 | ~v_510 | ~v_231 | ~v_2995 | ~v_2994 | ~v_230 | ~v_2993 | ~v_2992 | v_4022;
assign x_4976 = v_4021 | ~v_4018;
assign x_4977 = v_4021 | ~v_4019;
assign x_4978 = v_4021 | ~v_4020;
assign x_4979 = v_98 | v_103 | v_101 | v_97 | v_100 | v_93 | v_151 | v_170 | v_150 | v_148 | v_147 | v_184 | ~v_2267 | ~v_2266 | ~v_2265 | ~v_3979 | ~v_3978 | ~v_2264 | ~v_2263 | ~v_2262 | ~v_3977 | ~v_3976 | ~v_299 | ~v_2957 | ~v_2956 | ~v_2955 | ~v_298 | ~v_2954 | ~v_2953 | ~v_2952 | ~v_2299 | ~v_2298 | ~v_2297 | ~v_2296 | ~v_387 | ~v_2989 | ~v_2988 | ~v_386 | ~v_2987 | ~v_2986 | ~v_499 | ~v_498 | ~v_497 | ~v_496 | v_4020;
assign x_4980 = v_56 | v_55 | v_61 | v_51 | v_59 | v_58 | v_145 | v_143 | v_142 | v_166 | v_146 | v_183 | ~v_266 | ~v_2942 | ~v_2252 | ~v_2251 | ~v_2250 | ~v_3974 | ~v_3973 | ~v_2249 | ~v_2248 | ~v_2247 | ~v_3972 | ~v_3971 | ~v_2941 | ~v_2940 | ~v_265 | ~v_2939 | ~v_2938 | ~v_2937 | ~v_2294 | ~v_2293 | ~v_2292 | ~v_2291 | ~v_372 | ~v_2984 | ~v_2983 | ~v_371 | ~v_2982 | ~v_2981 | ~v_494 | ~v_493 | ~v_492 | ~v_491 | v_4019;
assign x_4981 = v_13 | v_18 | v_16 | v_8 | v_15 | v_12 | ~v_2927 | ~v_2926 | v_135 | v_134 | v_137 | v_138 | v_162 | v_182 | ~v_2237 | ~v_2236 | ~v_2235 | ~v_3969 | ~v_3968 | ~v_2234 | ~v_2233 | ~v_2232 | ~v_3967 | ~v_3966 | ~v_233 | ~v_2925 | ~v_2924 | ~v_232 | ~v_2923 | ~v_2922 | ~v_2289 | ~v_2288 | ~v_2287 | ~v_2286 | ~v_357 | ~v_2979 | ~v_2978 | ~v_356 | ~v_2977 | ~v_2976 | ~v_489 | ~v_488 | ~v_487 | ~v_486 | v_4018;
assign x_4982 = v_4017 | ~v_4014;
assign x_4983 = v_4017 | ~v_4015;
assign x_4984 = v_4017 | ~v_4016;
assign x_4985 = v_103 | v_101 | v_96 | v_100 | v_99 | v_102 | v_171 | v_170 | v_169 | v_149 | v_147 | v_184 | ~v_703 | ~v_702 | ~v_2331 | ~v_2330 | ~v_2265 | ~v_3979 | ~v_3978 | ~v_2329 | ~v_2328 | ~v_2262 | ~v_3977 | ~v_3976 | ~v_483 | ~v_3021 | ~v_3020 | ~v_2955 | ~v_482 | ~v_3019 | ~v_3018 | ~v_2952 | ~v_2283 | ~v_2282 | ~v_2281 | ~v_2280 | ~v_701 | ~v_653 | ~v_2973 | ~v_2972 | ~v_700 | ~v_652 | ~v_2971 | ~v_2970 | v_4016;
assign x_4986 = v_54 | v_61 | v_60 | v_59 | v_58 | v_57 | ~v_3016 | v_144 | v_142 | v_167 | v_166 | v_165 | v_183 | ~v_698 | ~v_697 | ~v_3015 | ~v_2326 | ~v_2325 | ~v_2250 | ~v_3974 | ~v_3973 | ~v_2324 | ~v_2323 | ~v_2247 | ~v_3972 | ~v_3971 | ~v_468 | ~v_2940 | ~v_467 | ~v_3014 | ~v_3013 | ~v_2937 | ~v_2278 | ~v_2277 | ~v_2276 | ~v_2275 | ~v_696 | ~v_638 | ~v_2968 | ~v_2967 | ~v_695 | ~v_637 | ~v_2966 | ~v_2965 | v_4015;
assign x_4987 = v_18 | v_17 | v_16 | v_15 | v_14 | v_11 | ~v_453 | ~v_2927 | ~v_452 | ~v_2926 | v_136 | v_134 | v_163 | v_162 | v_161 | v_182 | ~v_693 | ~v_692 | ~v_2321 | ~v_2320 | ~v_2235 | ~v_3969 | ~v_3968 | ~v_2319 | ~v_2318 | ~v_2232 | ~v_3967 | ~v_3966 | ~v_3011 | ~v_3010 | ~v_3009 | ~v_3008 | ~v_2273 | ~v_2272 | ~v_2271 | ~v_2270 | ~v_691 | ~v_623 | ~v_2963 | ~v_2962 | ~v_690 | ~v_622 | ~v_2961 | ~v_2960 | v_4014;
assign x_4988 = v_4013 | ~v_4010;
assign x_4989 = v_4013 | ~v_4011;
assign x_4990 = v_4013 | ~v_4012;
assign x_4991 = v_101 | v_97 | v_100 | v_102 | v_172 | v_171 | v_170 | v_169 | v_150 | v_148 | v_147 | v_184 | ~v_671 | ~v_670 | ~v_2265 | ~v_3979 | ~v_3978 | ~v_2262 | ~v_3977 | ~v_3976 | ~v_2955 | ~v_2952 | ~v_2299 | ~v_2298 | ~v_2297 | ~v_2296 | ~v_387 | ~v_2989 | ~v_2988 | ~v_386 | ~v_2987 | ~v_2986 | ~v_2283 | ~v_2282 | ~v_2281 | ~v_2280 | ~v_653 | ~v_2973 | ~v_2972 | ~v_652 | ~v_2971 | ~v_2970 | ~v_669 | ~v_668 | v_4012;
assign x_4992 = v_55 | v_60 | v_59 | v_58 | v_145 | v_143 | v_142 | v_168 | v_167 | v_166 | v_165 | v_183 | ~v_666 | ~v_665 | ~v_2250 | ~v_3974 | ~v_3973 | ~v_2247 | ~v_3972 | ~v_3971 | ~v_2940 | ~v_2937 | ~v_2294 | ~v_2293 | ~v_2292 | ~v_2291 | ~v_372 | ~v_2984 | ~v_2983 | ~v_371 | ~v_2982 | ~v_2981 | ~v_2278 | ~v_2277 | ~v_2276 | ~v_2275 | ~v_638 | ~v_2968 | ~v_2967 | ~v_637 | ~v_2966 | ~v_2965 | ~v_664 | ~v_663 | v_4011;
assign x_4993 = v_17 | v_16 | v_15 | v_12 | ~v_2927 | ~v_2926 | v_135 | v_134 | v_137 | v_164 | v_163 | v_162 | v_161 | v_182 | ~v_661 | ~v_660 | ~v_2235 | ~v_3969 | ~v_3968 | ~v_2232 | ~v_3967 | ~v_3966 | ~v_2289 | ~v_2288 | ~v_2287 | ~v_2286 | ~v_357 | ~v_2979 | ~v_2978 | ~v_356 | ~v_2977 | ~v_2976 | ~v_2273 | ~v_2272 | ~v_2271 | ~v_2270 | ~v_623 | ~v_2963 | ~v_2962 | ~v_622 | ~v_2961 | ~v_2960 | ~v_659 | ~v_658 | v_4010;
assign x_4994 = v_4009 | ~v_4006;
assign x_4995 = v_4009 | ~v_4007;
assign x_4996 = v_4009 | ~v_4008;
assign x_4997 = v_103 | v_101 | v_100 | v_95 | v_102 | v_171 | v_170 | v_169 | v_150 | v_149 | v_148 | v_184 | ~v_2265 | ~v_3979 | ~v_3978 | ~v_2262 | ~v_3977 | ~v_3976 | ~v_2955 | ~v_2952 | ~v_2261 | ~v_2260 | ~v_2259 | ~v_2258 | ~v_435 | ~v_2951 | ~v_2950 | ~v_434 | ~v_2949 | ~v_2948 | ~v_2283 | ~v_2282 | ~v_2281 | ~v_2280 | ~v_653 | ~v_2973 | ~v_2972 | ~v_652 | ~v_2971 | ~v_2970 | ~v_687 | ~v_686 | ~v_685 | ~v_684 | v_4008;
assign x_4998 = v_53 | v_61 | v_60 | v_59 | v_58 | v_144 | v_145 | v_143 | v_167 | v_166 | v_165 | v_183 | ~v_2250 | ~v_3974 | ~v_3973 | ~v_2247 | ~v_3972 | ~v_3971 | ~v_2940 | ~v_2937 | ~v_2246 | ~v_2245 | ~v_2244 | ~v_2243 | ~v_420 | ~v_2936 | ~v_2935 | ~v_419 | ~v_2934 | ~v_2933 | ~v_2278 | ~v_2277 | ~v_2276 | ~v_2275 | ~v_638 | ~v_2968 | ~v_2967 | ~v_637 | ~v_2966 | ~v_2965 | ~v_682 | ~v_681 | ~v_680 | ~v_679 | v_4007;
assign x_4999 = v_18 | v_17 | v_16 | v_15 | v_10 | ~v_2927 | ~v_2926 | v_136 | v_135 | v_137 | v_163 | v_162 | v_161 | v_182 | ~v_2235 | ~v_3969 | ~v_3968 | ~v_2232 | ~v_3967 | ~v_3966 | ~v_2231 | ~v_2230 | ~v_2229 | ~v_2228 | ~v_405 | ~v_2921 | ~v_2920 | ~v_404 | ~v_2919 | ~v_2918 | ~v_2273 | ~v_2272 | ~v_2271 | ~v_2270 | ~v_623 | ~v_2963 | ~v_2962 | ~v_622 | ~v_2961 | ~v_2960 | ~v_677 | ~v_676 | ~v_675 | ~v_674 | v_4006;
assign x_5000 = v_4005 | ~v_4002;
assign x_5001 = v_4005 | ~v_4003;
assign x_5002 = v_4005 | ~v_4004;
assign x_5003 = v_103 | v_100 | v_151 | v_171 | v_170 | v_169 | v_160 | v_150 | v_149 | v_148 | v_147 | v_184 | ~v_655 | ~v_654 | ~v_2265 | ~v_3979 | ~v_3978 | ~v_2262 | ~v_3977 | ~v_3976 | ~v_2955 | ~v_2952 | ~v_2315 | ~v_2314 | ~v_2313 | ~v_2312 | ~v_297 | ~v_3005 | ~v_3004 | ~v_296 | ~v_3003 | ~v_3002 | ~v_2283 | ~v_2282 | ~v_2281 | ~v_2280 | ~v_653 | ~v_2973 | ~v_2972 | ~v_652 | ~v_2971 | ~v_2970 | ~v_651 | ~v_650 | v_4004;
assign x_5004 = v_61 | v_58 | v_144 | v_159 | v_145 | v_143 | v_142 | v_167 | v_166 | v_165 | v_146 | v_183 | ~v_640 | ~v_639 | ~v_2250 | ~v_3974 | ~v_3973 | ~v_2247 | ~v_3972 | ~v_3971 | ~v_2940 | ~v_2937 | ~v_2310 | ~v_2309 | ~v_2308 | ~v_2307 | ~v_264 | ~v_3000 | ~v_2999 | ~v_263 | ~v_2998 | ~v_2997 | ~v_2278 | ~v_2277 | ~v_2276 | ~v_2275 | ~v_638 | ~v_2968 | ~v_2967 | ~v_637 | ~v_2966 | ~v_2965 | ~v_636 | ~v_635 | v_4003;
assign x_5005 = v_18 | v_15 | ~v_2927 | ~v_2926 | v_136 | v_135 | v_134 | v_137 | v_138 | v_163 | v_162 | v_161 | v_155 | v_182 | ~v_625 | ~v_624 | ~v_2235 | ~v_3969 | ~v_3968 | ~v_2232 | ~v_3967 | ~v_3966 | ~v_2305 | ~v_2304 | ~v_2303 | ~v_2302 | ~v_231 | ~v_2995 | ~v_2994 | ~v_230 | ~v_2993 | ~v_2992 | ~v_2273 | ~v_2272 | ~v_2271 | ~v_2270 | ~v_623 | ~v_2963 | ~v_2962 | ~v_622 | ~v_2961 | ~v_2960 | ~v_621 | ~v_620 | v_4002;
assign x_5006 = v_4001 | ~v_3998;
assign x_5007 = v_4001 | ~v_3999;
assign x_5008 = v_4001 | ~v_4000;
assign x_5009 = v_98 | v_103 | v_101 | v_100 | v_93 | v_102 | v_170 | v_150 | v_149 | v_148 | v_147 | v_184 | ~v_609 | ~v_608 | ~v_2267 | ~v_2266 | ~v_2265 | ~v_3979 | ~v_3978 | ~v_2264 | ~v_2263 | ~v_2262 | ~v_3977 | ~v_3976 | ~v_299 | ~v_2957 | ~v_2956 | ~v_2955 | ~v_298 | ~v_2954 | ~v_2953 | ~v_2952 | ~v_2261 | ~v_2260 | ~v_2259 | ~v_2258 | ~v_435 | ~v_2951 | ~v_2950 | ~v_434 | ~v_2949 | ~v_2948 | ~v_607 | ~v_606 | v_4000;
assign x_5010 = v_56 | v_61 | v_51 | v_60 | v_59 | v_58 | v_144 | v_145 | v_143 | v_142 | v_166 | v_183 | ~v_604 | ~v_603 | ~v_266 | ~v_2942 | ~v_2252 | ~v_2251 | ~v_2250 | ~v_3974 | ~v_3973 | ~v_2249 | ~v_2248 | ~v_2247 | ~v_3972 | ~v_3971 | ~v_2941 | ~v_2940 | ~v_265 | ~v_2939 | ~v_2938 | ~v_2937 | ~v_2246 | ~v_2245 | ~v_2244 | ~v_2243 | ~v_420 | ~v_2936 | ~v_2935 | ~v_419 | ~v_2934 | ~v_2933 | ~v_602 | ~v_601 | v_3999;
assign x_5011 = v_13 | v_18 | v_17 | v_16 | v_8 | v_15 | ~v_2927 | ~v_2926 | v_136 | v_135 | v_134 | v_137 | v_162 | v_182 | ~v_599 | ~v_598 | ~v_2237 | ~v_2236 | ~v_2235 | ~v_3969 | ~v_3968 | ~v_2234 | ~v_2233 | ~v_2232 | ~v_3967 | ~v_3966 | ~v_233 | ~v_2925 | ~v_2924 | ~v_232 | ~v_2923 | ~v_2922 | ~v_2231 | ~v_2230 | ~v_2229 | ~v_2228 | ~v_405 | ~v_2921 | ~v_2920 | ~v_404 | ~v_2919 | ~v_2918 | ~v_597 | ~v_596 | v_3998;
assign x_5012 = v_3997 | ~v_3994;
assign x_5013 = v_3997 | ~v_3995;
assign x_5014 = v_3997 | ~v_3996;
assign x_5015 = v_103 | v_101 | v_96 | v_99 | v_102 | v_171 | v_170 | v_169 | v_149 | v_147 | v_184 | v_181 | ~v_2331 | ~v_2330 | ~v_2265 | ~v_3979 | ~v_3978 | ~v_2329 | ~v_2328 | ~v_2262 | ~v_3977 | ~v_3976 | ~v_483 | ~v_3021 | ~v_3020 | ~v_2955 | ~v_482 | ~v_3019 | ~v_3018 | ~v_2952 | ~v_2383 | ~v_2382 | ~v_2381 | ~v_2380 | ~v_481 | ~v_480 | ~v_345 | ~v_3073 | ~v_3072 | ~v_479 | ~v_478 | ~v_344 | ~v_3071 | ~v_3070 | v_3996;
assign x_5016 = v_54 | v_61 | v_60 | v_59 | v_57 | ~v_3016 | v_144 | v_180 | v_142 | v_167 | v_166 | v_165 | v_183 | ~v_3015 | ~v_2326 | ~v_2325 | ~v_2250 | ~v_3974 | ~v_3973 | ~v_2324 | ~v_2323 | ~v_2247 | ~v_3972 | ~v_3971 | ~v_468 | ~v_2940 | ~v_467 | ~v_3014 | ~v_3013 | ~v_2937 | ~v_2378 | ~v_2377 | ~v_2376 | ~v_2375 | ~v_466 | ~v_465 | ~v_330 | ~v_3068 | ~v_3067 | ~v_464 | ~v_463 | ~v_329 | ~v_3066 | ~v_3065 | v_3995;
assign x_5017 = v_18 | v_17 | v_16 | v_14 | v_11 | ~v_453 | ~v_2927 | ~v_452 | ~v_2926 | v_136 | v_134 | v_179 | v_163 | v_162 | v_161 | v_182 | ~v_2321 | ~v_2320 | ~v_2235 | ~v_3969 | ~v_3968 | ~v_2319 | ~v_2318 | ~v_2232 | ~v_3967 | ~v_3966 | ~v_3011 | ~v_3010 | ~v_3009 | ~v_3008 | ~v_2373 | ~v_2372 | ~v_2371 | ~v_2370 | ~v_451 | ~v_450 | ~v_315 | ~v_3063 | ~v_3062 | ~v_449 | ~v_448 | ~v_314 | ~v_3061 | ~v_3060 | v_3994;
assign x_5018 = v_3993 | ~v_3990;
assign x_5019 = v_3993 | ~v_3991;
assign x_5020 = v_3993 | ~v_3992;
assign x_5021 = v_103 | v_101 | v_97 | v_102 | v_171 | v_170 | v_169 | v_150 | v_148 | v_147 | v_184 | v_181 | ~v_391 | ~v_390 | ~v_2265 | ~v_3979 | ~v_3978 | ~v_2262 | ~v_3977 | ~v_3976 | ~v_2955 | ~v_2952 | ~v_2299 | ~v_2298 | ~v_2297 | ~v_2296 | ~v_387 | ~v_2989 | ~v_2988 | ~v_386 | ~v_2987 | ~v_2986 | ~v_2383 | ~v_2382 | ~v_2381 | ~v_2380 | ~v_345 | ~v_3073 | ~v_3072 | ~v_344 | ~v_3071 | ~v_3070 | ~v_385 | ~v_384 | v_3992;
assign x_5022 = v_55 | v_61 | v_60 | v_59 | v_180 | v_145 | v_143 | v_142 | v_167 | v_166 | v_165 | v_183 | ~v_376 | ~v_375 | ~v_2250 | ~v_3974 | ~v_3973 | ~v_2247 | ~v_3972 | ~v_3971 | ~v_2940 | ~v_2937 | ~v_2294 | ~v_2293 | ~v_2292 | ~v_2291 | ~v_372 | ~v_2984 | ~v_2983 | ~v_371 | ~v_2982 | ~v_2981 | ~v_2378 | ~v_2377 | ~v_2376 | ~v_2375 | ~v_330 | ~v_3068 | ~v_3067 | ~v_329 | ~v_3066 | ~v_3065 | ~v_370 | ~v_369 | v_3991;
assign x_5023 = v_18 | v_17 | v_16 | v_12 | ~v_2927 | ~v_2926 | v_135 | v_134 | v_137 | v_179 | v_163 | v_162 | v_161 | v_182 | ~v_361 | ~v_360 | ~v_2235 | ~v_3969 | ~v_3968 | ~v_2232 | ~v_3967 | ~v_3966 | ~v_2289 | ~v_2288 | ~v_2287 | ~v_2286 | ~v_357 | ~v_2979 | ~v_2978 | ~v_356 | ~v_2977 | ~v_2976 | ~v_2373 | ~v_2372 | ~v_2371 | ~v_2370 | ~v_315 | ~v_3063 | ~v_3062 | ~v_314 | ~v_3061 | ~v_3060 | ~v_355 | ~v_354 | v_3990;
assign x_5024 = v_3989 | ~v_3986;
assign x_5025 = v_3989 | ~v_3987;
assign x_5026 = v_3989 | ~v_3988;
assign x_5027 = v_101 | v_102 | v_172 | v_171 | v_170 | v_169 | v_150 | v_149 | v_148 | v_147 | v_184 | v_181 | ~v_437 | ~v_436 | ~v_2265 | ~v_3979 | ~v_3978 | ~v_2262 | ~v_3977 | ~v_3976 | ~v_2955 | ~v_2952 | ~v_2261 | ~v_2260 | ~v_2259 | ~v_2258 | ~v_435 | ~v_2951 | ~v_2950 | ~v_434 | ~v_2949 | ~v_2948 | ~v_2383 | ~v_2382 | ~v_2381 | ~v_2380 | ~v_345 | ~v_3073 | ~v_3072 | ~v_344 | ~v_3071 | ~v_3070 | ~v_433 | ~v_432 | v_3988;
assign x_5028 = v_60 | v_59 | v_144 | v_180 | v_145 | v_143 | v_142 | v_168 | v_167 | v_166 | v_165 | v_183 | ~v_422 | ~v_421 | ~v_2250 | ~v_3974 | ~v_3973 | ~v_2247 | ~v_3972 | ~v_3971 | ~v_2940 | ~v_2937 | ~v_2246 | ~v_2245 | ~v_2244 | ~v_2243 | ~v_420 | ~v_2936 | ~v_2935 | ~v_419 | ~v_2934 | ~v_2933 | ~v_2378 | ~v_2377 | ~v_2376 | ~v_2375 | ~v_330 | ~v_3068 | ~v_3067 | ~v_329 | ~v_3066 | ~v_3065 | ~v_418 | ~v_417 | v_3987;
assign x_5029 = v_17 | v_16 | ~v_2927 | ~v_2926 | v_136 | v_135 | v_134 | v_137 | v_179 | v_164 | v_163 | v_162 | v_161 | v_182 | ~v_407 | ~v_406 | ~v_2235 | ~v_3969 | ~v_3968 | ~v_2232 | ~v_3967 | ~v_3966 | ~v_2231 | ~v_2230 | ~v_2229 | ~v_2228 | ~v_405 | ~v_2921 | ~v_2920 | ~v_404 | ~v_2919 | ~v_2918 | ~v_2373 | ~v_2372 | ~v_2371 | ~v_2370 | ~v_315 | ~v_3063 | ~v_3062 | ~v_314 | ~v_3061 | ~v_3060 | ~v_403 | ~v_402 | v_3986;
assign x_5030 = v_3985 | ~v_3982;
assign x_5031 = v_3985 | ~v_3983;
assign x_5032 = v_3985 | ~v_3984;
assign x_5033 = v_103 | v_95 | v_102 | v_171 | v_170 | v_169 | v_160 | v_150 | v_149 | v_148 | v_184 | v_181 | ~v_2265 | ~v_3979 | ~v_3978 | ~v_2262 | ~v_3977 | ~v_3976 | ~v_2955 | ~v_2952 | ~v_2315 | ~v_2314 | ~v_2313 | ~v_2312 | ~v_297 | ~v_3005 | ~v_3004 | ~v_296 | ~v_3003 | ~v_3002 | ~v_2383 | ~v_2382 | ~v_2381 | ~v_2380 | ~v_345 | ~v_3073 | ~v_3072 | ~v_344 | ~v_3071 | ~v_3070 | ~v_343 | ~v_342 | ~v_341 | ~v_340 | v_3984;
assign x_5034 = v_53 | v_61 | v_60 | v_144 | v_180 | v_159 | v_145 | v_143 | v_167 | v_166 | v_165 | v_183 | ~v_2250 | ~v_3974 | ~v_3973 | ~v_2247 | ~v_3972 | ~v_3971 | ~v_2940 | ~v_2937 | ~v_2310 | ~v_2309 | ~v_2308 | ~v_2307 | ~v_264 | ~v_3000 | ~v_2999 | ~v_263 | ~v_2998 | ~v_2997 | ~v_2378 | ~v_2377 | ~v_2376 | ~v_2375 | ~v_330 | ~v_3068 | ~v_3067 | ~v_329 | ~v_3066 | ~v_3065 | ~v_328 | ~v_327 | ~v_326 | ~v_325 | v_3983;
assign x_5035 = v_18 | v_17 | v_10 | ~v_2927 | ~v_2926 | v_136 | v_135 | v_137 | v_179 | v_163 | v_162 | v_161 | v_155 | v_182 | ~v_2235 | ~v_3969 | ~v_3968 | ~v_2232 | ~v_3967 | ~v_3966 | ~v_2305 | ~v_2304 | ~v_2303 | ~v_2302 | ~v_231 | ~v_2995 | ~v_2994 | ~v_230 | ~v_2993 | ~v_2992 | ~v_2373 | ~v_2372 | ~v_2371 | ~v_2370 | ~v_315 | ~v_3063 | ~v_3062 | ~v_314 | ~v_3061 | ~v_3060 | ~v_313 | ~v_312 | ~v_311 | ~v_310 | v_3982;
assign x_5036 = v_3981 | ~v_3970;
assign x_5037 = v_3981 | ~v_3975;
assign x_5038 = v_3981 | ~v_3980;
assign x_5039 = v_98 | v_103 | v_100 | v_93 | v_102 | v_170 | v_160 | v_150 | v_149 | v_148 | v_147 | v_184 | ~v_2267 | ~v_2266 | ~v_2265 | ~v_3979 | ~v_3978 | ~v_2264 | ~v_2263 | ~v_2262 | ~v_3977 | ~v_3976 | ~v_299 | ~v_2957 | ~v_2956 | ~v_2955 | ~v_298 | ~v_2954 | ~v_2953 | ~v_2952 | ~v_2315 | ~v_2314 | ~v_2313 | ~v_2312 | ~v_297 | ~v_3005 | ~v_3004 | ~v_296 | ~v_3003 | ~v_3002 | ~v_295 | ~v_294 | ~v_293 | ~v_292 | v_3980;
assign x_5040 = v_3979 | v_140;
assign x_5041 = v_3979 | v_123;
assign x_5042 = v_3978 | v_139;
assign x_5043 = v_3978 | v_120;
assign x_5044 = v_3977 | ~v_140;
assign x_5045 = v_3977 | v_108;
assign x_5046 = v_3976 | ~v_139;
assign x_5047 = v_3976 | v_105;
assign x_5048 = v_56 | v_61 | v_51 | v_60 | v_58 | v_144 | v_159 | v_145 | v_143 | v_142 | v_166 | v_183 | ~v_266 | ~v_2942 | ~v_2252 | ~v_2251 | ~v_2250 | ~v_3974 | ~v_3973 | ~v_2249 | ~v_2248 | ~v_2247 | ~v_3972 | ~v_3971 | ~v_2941 | ~v_2940 | ~v_265 | ~v_2939 | ~v_2938 | ~v_2937 | ~v_2310 | ~v_2309 | ~v_2308 | ~v_2307 | ~v_264 | ~v_3000 | ~v_2999 | ~v_263 | ~v_2998 | ~v_2997 | ~v_262 | ~v_261 | ~v_260 | ~v_259 | v_3975;
assign x_5049 = v_3974 | v_140;
assign x_5050 = v_3974 | v_81;
assign x_5051 = v_3973 | v_139;
assign x_5052 = v_3973 | v_78;
assign x_5053 = v_3972 | ~v_140;
assign x_5054 = v_3972 | v_66;
assign x_5055 = v_3971 | ~v_139;
assign x_5056 = v_3971 | v_63;
assign x_5057 = v_13 | v_18 | v_17 | v_8 | v_15 | ~v_2927 | ~v_2926 | v_136 | v_135 | v_134 | v_137 | v_162 | v_155 | v_182 | ~v_2237 | ~v_2236 | ~v_2235 | ~v_3969 | ~v_3968 | ~v_2234 | ~v_2233 | ~v_2232 | ~v_3967 | ~v_3966 | ~v_233 | ~v_2925 | ~v_2924 | ~v_232 | ~v_2923 | ~v_2922 | ~v_2305 | ~v_2304 | ~v_2303 | ~v_2302 | ~v_231 | ~v_2995 | ~v_2994 | ~v_230 | ~v_2993 | ~v_2992 | ~v_229 | ~v_228 | ~v_227 | ~v_226 | v_3970;
assign x_5058 = v_3969 | v_140;
assign x_5059 = v_3969 | v_39;
assign x_5060 = v_3968 | v_139;
assign x_5061 = v_3968 | v_36;
assign x_5062 = v_3967 | ~v_140;
assign x_5063 = v_3967 | v_24;
assign x_5064 = v_3966 | ~v_139;
assign x_5065 = v_3966 | v_21;
assign x_5066 = v_3965 | ~v_3963;
assign x_5067 = v_3965 | ~v_3964;
assign x_5068 = v_3965 | ~v_2219;
assign x_5069 = v_3965 | ~v_2220;
assign x_5070 = v_3965 | ~v_140;
assign x_5071 = v_3965 | ~v_139;
assign x_5072 = ~v_193 | ~v_1272 | v_3964;
assign x_5073 = ~v_185 | ~v_191 | v_3963;
assign x_5074 = v_3962 | ~v_3881;
assign x_5075 = v_3962 | ~v_3961;
assign x_5076 = v_152 | v_153 | ~v_3960 | ~v_1565 | ~v_1564 | ~v_3883 | ~v_3882 | v_3961;
assign x_5077 = v_3960 | ~v_3899;
assign x_5078 = v_3960 | ~v_3903;
assign x_5079 = v_3960 | ~v_3907;
assign x_5080 = v_3960 | ~v_3911;
assign x_5081 = v_3960 | ~v_3915;
assign x_5082 = v_3960 | ~v_3919;
assign x_5083 = v_3960 | ~v_3923;
assign x_5084 = v_3960 | ~v_3927;
assign x_5085 = v_3960 | ~v_3931;
assign x_5086 = v_3960 | ~v_3935;
assign x_5087 = v_3960 | ~v_3939;
assign x_5088 = v_3960 | ~v_3943;
assign x_5089 = v_3960 | ~v_3947;
assign x_5090 = v_3960 | ~v_3951;
assign x_5091 = v_3960 | ~v_3955;
assign x_5092 = v_3960 | ~v_3959;
assign x_5093 = v_3960 | ~v_1263;
assign x_5094 = v_3960 | ~v_1264;
assign x_5095 = v_3960 | ~v_1265;
assign x_5096 = v_3960 | ~v_1266;
assign x_5097 = ~v_3958 | ~v_3957 | ~v_3956 | v_3959;
assign x_5098 = v_3958 | ~v_827;
assign x_5099 = v_3958 | ~v_3894;
assign x_5100 = v_3958 | ~v_828;
assign x_5101 = v_3958 | ~v_1015;
assign x_5102 = v_3958 | ~v_3895;
assign x_5103 = v_3958 | ~v_829;
assign x_5104 = v_3958 | ~v_1016;
assign x_5105 = v_3958 | ~v_830;
assign x_5106 = v_3958 | ~v_3896;
assign x_5107 = v_3958 | ~v_831;
assign x_5108 = v_3958 | ~v_1017;
assign x_5109 = v_3958 | ~v_3897;
assign x_5110 = v_3958 | ~v_832;
assign x_5111 = v_3958 | ~v_1018;
assign x_5112 = v_3958 | ~v_3496;
assign x_5113 = v_3958 | ~v_3497;
assign x_5114 = v_3958 | ~v_3564;
assign x_5115 = v_3958 | ~v_3498;
assign x_5116 = v_3958 | ~v_3565;
assign x_5117 = v_3958 | ~v_3499;
assign x_5118 = v_3958 | ~v_3500;
assign x_5119 = v_3958 | ~v_3566;
assign x_5120 = v_3958 | ~v_3501;
assign x_5121 = v_3958 | ~v_3567;
assign x_5122 = v_3958 | ~v_839;
assign x_5123 = v_3958 | ~v_1257;
assign x_5124 = v_3958 | ~v_1023;
assign x_5125 = v_3958 | ~v_840;
assign x_5126 = v_3958 | ~v_1258;
assign x_5127 = v_3958 | ~v_1024;
assign x_5128 = v_3958 | ~v_184;
assign x_5129 = v_3958 | ~v_169;
assign x_5130 = v_3958 | ~v_148;
assign x_5131 = v_3958 | ~v_1259;
assign x_5132 = v_3958 | ~v_1260;
assign x_5133 = v_3958 | ~v_103;
assign x_5134 = v_3958 | ~v_102;
assign x_5135 = v_3958 | ~v_101;
assign x_5136 = v_3958 | ~v_100;
assign x_5137 = v_3958 | ~v_99;
assign x_5138 = v_3958 | ~v_98;
assign x_5139 = v_3958 | ~v_97;
assign x_5140 = v_3958 | ~v_95;
assign x_5141 = v_3958 | ~v_94;
assign x_5142 = v_3957 | ~v_794;
assign x_5143 = v_3957 | ~v_3889;
assign x_5144 = v_3957 | ~v_795;
assign x_5145 = v_3957 | ~v_1000;
assign x_5146 = v_3957 | ~v_3890;
assign x_5147 = v_3957 | ~v_796;
assign x_5148 = v_3957 | ~v_1001;
assign x_5149 = v_3957 | ~v_797;
assign x_5150 = v_3957 | ~v_3891;
assign x_5151 = v_3957 | ~v_798;
assign x_5152 = v_3957 | ~v_1002;
assign x_5153 = v_3957 | ~v_3892;
assign x_5154 = v_3957 | ~v_799;
assign x_5155 = v_3957 | ~v_1003;
assign x_5156 = v_3957 | ~v_3481;
assign x_5157 = v_3957 | ~v_3482;
assign x_5158 = v_3957 | ~v_3559;
assign x_5159 = v_3957 | ~v_3483;
assign x_5160 = v_3957 | ~v_3560;
assign x_5161 = v_3957 | ~v_3484;
assign x_5162 = v_3957 | ~v_3485;
assign x_5163 = v_3957 | ~v_806;
assign x_5164 = v_3957 | ~v_1252;
assign x_5165 = v_3957 | ~v_1008;
assign x_5166 = v_3957 | ~v_1253;
assign x_5167 = v_3957 | ~v_1009;
assign x_5168 = v_3957 | ~v_3561;
assign x_5169 = v_3957 | ~v_807;
assign x_5170 = v_3957 | ~v_3486;
assign x_5171 = v_3957 | ~v_3562;
assign x_5172 = v_3957 | ~v_183;
assign x_5173 = v_3957 | ~v_165;
assign x_5174 = v_3957 | ~v_143;
assign x_5175 = v_3957 | ~v_1254;
assign x_5176 = v_3957 | ~v_1255;
assign x_5177 = v_3957 | ~v_61;
assign x_5178 = v_3957 | ~v_60;
assign x_5179 = v_3957 | ~v_59;
assign x_5180 = v_3957 | ~v_58;
assign x_5181 = v_3957 | ~v_57;
assign x_5182 = v_3957 | ~v_56;
assign x_5183 = v_3957 | ~v_55;
assign x_5184 = v_3957 | ~v_53;
assign x_5185 = v_3957 | ~v_52;
assign x_5186 = v_3956 | ~v_761;
assign x_5187 = v_3956 | ~v_3884;
assign x_5188 = v_3956 | ~v_762;
assign x_5189 = v_3956 | ~v_985;
assign x_5190 = v_3956 | ~v_3885;
assign x_5191 = v_3956 | ~v_763;
assign x_5192 = v_3956 | ~v_986;
assign x_5193 = v_3956 | ~v_764;
assign x_5194 = v_3956 | ~v_3886;
assign x_5195 = v_3956 | ~v_765;
assign x_5196 = v_3956 | ~v_987;
assign x_5197 = v_3956 | ~v_3887;
assign x_5198 = v_3956 | ~v_766;
assign x_5199 = v_3956 | ~v_988;
assign x_5200 = v_3956 | ~v_3466;
assign x_5201 = v_3956 | ~v_3467;
assign x_5202 = v_3956 | ~v_3554;
assign x_5203 = v_3956 | ~v_3468;
assign x_5204 = v_3956 | ~v_3555;
assign x_5205 = v_3956 | ~v_3469;
assign x_5206 = v_3956 | ~v_3556;
assign x_5207 = v_3956 | ~v_3470;
assign x_5208 = v_3956 | ~v_3557;
assign x_5209 = v_3956 | ~v_773;
assign x_5210 = v_3956 | ~v_774;
assign x_5211 = v_3956 | ~v_182;
assign x_5212 = v_3956 | ~v_161;
assign x_5213 = v_3956 | ~v_3473;
assign x_5214 = v_3956 | ~v_1247;
assign x_5215 = v_3956 | ~v_1248;
assign x_5216 = v_3956 | ~v_135;
assign x_5217 = v_3956 | ~v_1249;
assign x_5218 = v_3956 | ~v_993;
assign x_5219 = v_3956 | ~v_1250;
assign x_5220 = v_3956 | ~v_994;
assign x_5221 = v_3956 | ~v_18;
assign x_5222 = v_3956 | ~v_17;
assign x_5223 = v_3956 | ~v_16;
assign x_5224 = v_3956 | ~v_15;
assign x_5225 = v_3956 | ~v_14;
assign x_5226 = v_3956 | ~v_13;
assign x_5227 = v_3956 | ~v_12;
assign x_5228 = v_3956 | ~v_10;
assign x_5229 = v_3956 | ~v_9;
assign x_5230 = ~v_3954 | ~v_3953 | ~v_3952 | v_3955;
assign x_5231 = v_3954 | ~v_1187;
assign x_5232 = v_3954 | ~v_1188;
assign x_5233 = v_3954 | ~v_1189;
assign x_5234 = v_3954 | ~v_1190;
assign x_5235 = v_3954 | ~v_827;
assign x_5236 = v_3954 | ~v_3894;
assign x_5237 = v_3954 | ~v_1015;
assign x_5238 = v_3954 | ~v_3895;
assign x_5239 = v_3954 | ~v_1016;
assign x_5240 = v_3954 | ~v_830;
assign x_5241 = v_3954 | ~v_3896;
assign x_5242 = v_3954 | ~v_1017;
assign x_5243 = v_3954 | ~v_3897;
assign x_5244 = v_3954 | ~v_1018;
assign x_5245 = v_3954 | ~v_3516;
assign x_5246 = v_3954 | ~v_3517;
assign x_5247 = v_3954 | ~v_3518;
assign x_5248 = v_3954 | ~v_3519;
assign x_5249 = v_3954 | ~v_3496;
assign x_5250 = v_3954 | ~v_3564;
assign x_5251 = v_3954 | ~v_3565;
assign x_5252 = v_3954 | ~v_3499;
assign x_5253 = v_3954 | ~v_3566;
assign x_5254 = v_3954 | ~v_3567;
assign x_5255 = v_3954 | ~v_1193;
assign x_5256 = v_3954 | ~v_1241;
assign x_5257 = v_3954 | ~v_1194;
assign x_5258 = v_3954 | ~v_1242;
assign x_5259 = v_3954 | ~v_1023;
assign x_5260 = v_3954 | ~v_1024;
assign x_5261 = v_3954 | ~v_1243;
assign x_5262 = v_3954 | ~v_1244;
assign x_5263 = v_3954 | ~v_184;
assign x_5264 = v_3954 | ~v_171;
assign x_5265 = v_3954 | ~v_170;
assign x_5266 = v_3954 | ~v_148;
assign x_5267 = v_3954 | ~v_147;
assign x_5268 = v_3954 | ~v_103;
assign x_5269 = v_3954 | ~v_102;
assign x_5270 = v_3954 | ~v_101;
assign x_5271 = v_3954 | ~v_100;
assign x_5272 = v_3954 | ~v_99;
assign x_5273 = v_3954 | ~v_97;
assign x_5274 = v_3954 | ~v_93;
assign x_5275 = v_3953 | ~v_1172;
assign x_5276 = v_3953 | ~v_1173;
assign x_5277 = v_3953 | ~v_1174;
assign x_5278 = v_3953 | ~v_1175;
assign x_5279 = v_3953 | ~v_794;
assign x_5280 = v_3953 | ~v_3889;
assign x_5281 = v_3953 | ~v_1000;
assign x_5282 = v_3953 | ~v_3890;
assign x_5283 = v_3953 | ~v_1001;
assign x_5284 = v_3953 | ~v_797;
assign x_5285 = v_3953 | ~v_3891;
assign x_5286 = v_3953 | ~v_1002;
assign x_5287 = v_3953 | ~v_3892;
assign x_5288 = v_3953 | ~v_1003;
assign x_5289 = v_3953 | ~v_3511;
assign x_5290 = v_3953 | ~v_3512;
assign x_5291 = v_3953 | ~v_3513;
assign x_5292 = v_3953 | ~v_3514;
assign x_5293 = v_3953 | ~v_3481;
assign x_5294 = v_3953 | ~v_3559;
assign x_5295 = v_3953 | ~v_3560;
assign x_5296 = v_3953 | ~v_3484;
assign x_5297 = v_3953 | ~v_1178;
assign x_5298 = v_3953 | ~v_1236;
assign x_5299 = v_3953 | ~v_1179;
assign x_5300 = v_3953 | ~v_1237;
assign x_5301 = v_3953 | ~v_1008;
assign x_5302 = v_3953 | ~v_1009;
assign x_5303 = v_3953 | ~v_3561;
assign x_5304 = v_3953 | ~v_3562;
assign x_5305 = v_3953 | ~v_1238;
assign x_5306 = v_3953 | ~v_1239;
assign x_5307 = v_3953 | ~v_183;
assign x_5308 = v_3953 | ~v_167;
assign x_5309 = v_3953 | ~v_166;
assign x_5310 = v_3953 | ~v_143;
assign x_5311 = v_3953 | ~v_142;
assign x_5312 = v_3953 | ~v_61;
assign x_5313 = v_3953 | ~v_60;
assign x_5314 = v_3953 | ~v_59;
assign x_5315 = v_3953 | ~v_58;
assign x_5316 = v_3953 | ~v_57;
assign x_5317 = v_3953 | ~v_55;
assign x_5318 = v_3953 | ~v_51;
assign x_5319 = v_3952 | ~v_1157;
assign x_5320 = v_3952 | ~v_1158;
assign x_5321 = v_3952 | ~v_1159;
assign x_5322 = v_3952 | ~v_1160;
assign x_5323 = v_3952 | ~v_761;
assign x_5324 = v_3952 | ~v_3884;
assign x_5325 = v_3952 | ~v_985;
assign x_5326 = v_3952 | ~v_3885;
assign x_5327 = v_3952 | ~v_986;
assign x_5328 = v_3952 | ~v_764;
assign x_5329 = v_3952 | ~v_3886;
assign x_5330 = v_3952 | ~v_987;
assign x_5331 = v_3952 | ~v_3887;
assign x_5332 = v_3952 | ~v_988;
assign x_5333 = v_3952 | ~v_3506;
assign x_5334 = v_3952 | ~v_3507;
assign x_5335 = v_3952 | ~v_3508;
assign x_5336 = v_3952 | ~v_3509;
assign x_5337 = v_3952 | ~v_3466;
assign x_5338 = v_3952 | ~v_3554;
assign x_5339 = v_3952 | ~v_3555;
assign x_5340 = v_3952 | ~v_3469;
assign x_5341 = v_3952 | ~v_3556;
assign x_5342 = v_3952 | ~v_3557;
assign x_5343 = v_3952 | ~v_1163;
assign x_5344 = v_3952 | ~v_1231;
assign x_5345 = v_3952 | ~v_1164;
assign x_5346 = v_3952 | ~v_1232;
assign x_5347 = v_3952 | ~v_1233;
assign x_5348 = v_3952 | ~v_1234;
assign x_5349 = v_3952 | ~v_182;
assign x_5350 = v_3952 | ~v_163;
assign x_5351 = v_3952 | ~v_162;
assign x_5352 = v_3952 | ~v_135;
assign x_5353 = v_3952 | ~v_134;
assign x_5354 = v_3952 | ~v_993;
assign x_5355 = v_3952 | ~v_994;
assign x_5356 = v_3952 | ~v_18;
assign x_5357 = v_3952 | ~v_17;
assign x_5358 = v_3952 | ~v_16;
assign x_5359 = v_3952 | ~v_15;
assign x_5360 = v_3952 | ~v_14;
assign x_5361 = v_3952 | ~v_12;
assign x_5362 = v_3952 | ~v_8;
assign x_5363 = ~v_3950 | ~v_3949 | ~v_3948 | v_3951;
assign x_5364 = v_3950 | ~v_969;
assign x_5365 = v_3950 | ~v_970;
assign x_5366 = v_3950 | ~v_971;
assign x_5367 = v_3950 | ~v_972;
assign x_5368 = v_3950 | ~v_1187;
assign x_5369 = v_3950 | ~v_1188;
assign x_5370 = v_3950 | ~v_1189;
assign x_5371 = v_3950 | ~v_1190;
assign x_5372 = v_3950 | ~v_827;
assign x_5373 = v_3950 | ~v_3894;
assign x_5374 = v_3950 | ~v_3895;
assign x_5375 = v_3950 | ~v_830;
assign x_5376 = v_3950 | ~v_3896;
assign x_5377 = v_3950 | ~v_3897;
assign x_5378 = v_3950 | ~v_3516;
assign x_5379 = v_3950 | ~v_3517;
assign x_5380 = v_3950 | ~v_3518;
assign x_5381 = v_3950 | ~v_3519;
assign x_5382 = v_3950 | ~v_3494;
assign x_5383 = v_3950 | ~v_3495;
assign x_5384 = v_3950 | ~v_3496;
assign x_5385 = v_3950 | ~v_3499;
assign x_5386 = v_3950 | ~v_1225;
assign x_5387 = v_3950 | ~v_1226;
assign x_5388 = v_3950 | ~v_1227;
assign x_5389 = v_3950 | ~v_1228;
assign x_5390 = v_3950 | ~v_1193;
assign x_5391 = v_3950 | ~v_1194;
assign x_5392 = v_3950 | ~v_975;
assign x_5393 = v_3950 | ~v_976;
assign x_5394 = v_3950 | ~v_3502;
assign x_5395 = v_3950 | ~v_3503;
assign x_5396 = v_3950 | ~v_184;
assign x_5397 = v_3950 | ~v_171;
assign x_5398 = v_3950 | ~v_170;
assign x_5399 = v_3950 | ~v_150;
assign x_5400 = v_3950 | ~v_149;
assign x_5401 = v_3950 | ~v_103;
assign x_5402 = v_3950 | ~v_102;
assign x_5403 = v_3950 | ~v_101;
assign x_5404 = v_3950 | ~v_100;
assign x_5405 = v_3950 | ~v_96;
assign x_5406 = v_3950 | ~v_95;
assign x_5407 = v_3950 | ~v_93;
assign x_5408 = v_3949 | ~v_954;
assign x_5409 = v_3949 | ~v_955;
assign x_5410 = v_3949 | ~v_956;
assign x_5411 = v_3949 | ~v_957;
assign x_5412 = v_3949 | ~v_1172;
assign x_5413 = v_3949 | ~v_1173;
assign x_5414 = v_3949 | ~v_1174;
assign x_5415 = v_3949 | ~v_1175;
assign x_5416 = v_3949 | ~v_794;
assign x_5417 = v_3949 | ~v_3889;
assign x_5418 = v_3949 | ~v_3890;
assign x_5419 = v_3949 | ~v_797;
assign x_5420 = v_3949 | ~v_3891;
assign x_5421 = v_3949 | ~v_3892;
assign x_5422 = v_3949 | ~v_3511;
assign x_5423 = v_3949 | ~v_3512;
assign x_5424 = v_3949 | ~v_3513;
assign x_5425 = v_3949 | ~v_3514;
assign x_5426 = v_3949 | ~v_3479;
assign x_5427 = v_3949 | ~v_3480;
assign x_5428 = v_3949 | ~v_3481;
assign x_5429 = v_3949 | ~v_3484;
assign x_5430 = v_3949 | ~v_1220;
assign x_5431 = v_3949 | ~v_1221;
assign x_5432 = v_3949 | ~v_1222;
assign x_5433 = v_3949 | ~v_1223;
assign x_5434 = v_3949 | ~v_1178;
assign x_5435 = v_3949 | ~v_1179;
assign x_5436 = v_3949 | ~v_960;
assign x_5437 = v_3949 | ~v_961;
assign x_5438 = v_3949 | ~v_3487;
assign x_5439 = v_3949 | ~v_3488;
assign x_5440 = v_3949 | ~v_183;
assign x_5441 = v_3949 | ~v_167;
assign x_5442 = v_3949 | ~v_166;
assign x_5443 = v_3949 | ~v_145;
assign x_5444 = v_3949 | ~v_144;
assign x_5445 = v_3949 | ~v_61;
assign x_5446 = v_3949 | ~v_60;
assign x_5447 = v_3949 | ~v_59;
assign x_5448 = v_3949 | ~v_58;
assign x_5449 = v_3949 | ~v_54;
assign x_5450 = v_3949 | ~v_53;
assign x_5451 = v_3949 | ~v_51;
assign x_5452 = v_3948 | ~v_939;
assign x_5453 = v_3948 | ~v_940;
assign x_5454 = v_3948 | ~v_941;
assign x_5455 = v_3948 | ~v_942;
assign x_5456 = v_3948 | ~v_1157;
assign x_5457 = v_3948 | ~v_1158;
assign x_5458 = v_3948 | ~v_1159;
assign x_5459 = v_3948 | ~v_1160;
assign x_5460 = v_3948 | ~v_761;
assign x_5461 = v_3948 | ~v_3884;
assign x_5462 = v_3948 | ~v_3885;
assign x_5463 = v_3948 | ~v_764;
assign x_5464 = v_3948 | ~v_3886;
assign x_5465 = v_3948 | ~v_3887;
assign x_5466 = v_3948 | ~v_3506;
assign x_5467 = v_3948 | ~v_3507;
assign x_5468 = v_3948 | ~v_3508;
assign x_5469 = v_3948 | ~v_3509;
assign x_5470 = v_3948 | ~v_3464;
assign x_5471 = v_3948 | ~v_3465;
assign x_5472 = v_3948 | ~v_3466;
assign x_5473 = v_3948 | ~v_3469;
assign x_5474 = v_3948 | ~v_1215;
assign x_5475 = v_3948 | ~v_1216;
assign x_5476 = v_3948 | ~v_1217;
assign x_5477 = v_3948 | ~v_1218;
assign x_5478 = v_3948 | ~v_1163;
assign x_5479 = v_3948 | ~v_1164;
assign x_5480 = v_3948 | ~v_945;
assign x_5481 = v_3948 | ~v_946;
assign x_5482 = v_3948 | ~v_3471;
assign x_5483 = v_3948 | ~v_3472;
assign x_5484 = v_3948 | ~v_182;
assign x_5485 = v_3948 | ~v_163;
assign x_5486 = v_3948 | ~v_162;
assign x_5487 = v_3948 | ~v_137;
assign x_5488 = v_3948 | ~v_136;
assign x_5489 = v_3948 | ~v_18;
assign x_5490 = v_3948 | ~v_17;
assign x_5491 = v_3948 | ~v_16;
assign x_5492 = v_3948 | ~v_15;
assign x_5493 = v_3948 | ~v_11;
assign x_5494 = v_3948 | ~v_10;
assign x_5495 = v_3948 | ~v_8;
assign x_5496 = ~v_3946 | ~v_3945 | ~v_3944 | v_3947;
assign x_5497 = v_3946 | ~v_921;
assign x_5498 = v_3946 | ~v_922;
assign x_5499 = v_3946 | ~v_923;
assign x_5500 = v_3946 | ~v_924;
assign x_5501 = v_3946 | ~v_1187;
assign x_5502 = v_3946 | ~v_1188;
assign x_5503 = v_3946 | ~v_1189;
assign x_5504 = v_3946 | ~v_1190;
assign x_5505 = v_3946 | ~v_827;
assign x_5506 = v_3946 | ~v_3894;
assign x_5507 = v_3946 | ~v_3895;
assign x_5508 = v_3946 | ~v_830;
assign x_5509 = v_3946 | ~v_3896;
assign x_5510 = v_3946 | ~v_3897;
assign x_5511 = v_3946 | ~v_3516;
assign x_5512 = v_3946 | ~v_3517;
assign x_5513 = v_3946 | ~v_3518;
assign x_5514 = v_3946 | ~v_3519;
assign x_5515 = v_3946 | ~v_3532;
assign x_5516 = v_3946 | ~v_3533;
assign x_5517 = v_3946 | ~v_3534;
assign x_5518 = v_3946 | ~v_3535;
assign x_5519 = v_3946 | ~v_3496;
assign x_5520 = v_3946 | ~v_3499;
assign x_5521 = v_3946 | ~v_1209;
assign x_5522 = v_3946 | ~v_1210;
assign x_5523 = v_3946 | ~v_1193;
assign x_5524 = v_3946 | ~v_1194;
assign x_5525 = v_3946 | ~v_927;
assign x_5526 = v_3946 | ~v_928;
assign x_5527 = v_3946 | ~v_1211;
assign x_5528 = v_3946 | ~v_1212;
assign x_5529 = v_3946 | ~v_184;
assign x_5530 = v_3946 | ~v_172;
assign x_5531 = v_3946 | ~v_171;
assign x_5532 = v_3946 | ~v_170;
assign x_5533 = v_3946 | ~v_150;
assign x_5534 = v_3946 | ~v_149;
assign x_5535 = v_3946 | ~v_148;
assign x_5536 = v_3946 | ~v_147;
assign x_5537 = v_3946 | ~v_102;
assign x_5538 = v_3946 | ~v_101;
assign x_5539 = v_3946 | ~v_100;
assign x_5540 = v_3946 | ~v_93;
assign x_5541 = v_3945 | ~v_906;
assign x_5542 = v_3945 | ~v_907;
assign x_5543 = v_3945 | ~v_908;
assign x_5544 = v_3945 | ~v_909;
assign x_5545 = v_3945 | ~v_1172;
assign x_5546 = v_3945 | ~v_1173;
assign x_5547 = v_3945 | ~v_1174;
assign x_5548 = v_3945 | ~v_1175;
assign x_5549 = v_3945 | ~v_794;
assign x_5550 = v_3945 | ~v_3889;
assign x_5551 = v_3945 | ~v_3890;
assign x_5552 = v_3945 | ~v_797;
assign x_5553 = v_3945 | ~v_3891;
assign x_5554 = v_3945 | ~v_3892;
assign x_5555 = v_3945 | ~v_3511;
assign x_5556 = v_3945 | ~v_3512;
assign x_5557 = v_3945 | ~v_3513;
assign x_5558 = v_3945 | ~v_3514;
assign x_5559 = v_3945 | ~v_3527;
assign x_5560 = v_3945 | ~v_3528;
assign x_5561 = v_3945 | ~v_3529;
assign x_5562 = v_3945 | ~v_3530;
assign x_5563 = v_3945 | ~v_3481;
assign x_5564 = v_3945 | ~v_3484;
assign x_5565 = v_3945 | ~v_1204;
assign x_5566 = v_3945 | ~v_1205;
assign x_5567 = v_3945 | ~v_1178;
assign x_5568 = v_3945 | ~v_1179;
assign x_5569 = v_3945 | ~v_912;
assign x_5570 = v_3945 | ~v_913;
assign x_5571 = v_3945 | ~v_1206;
assign x_5572 = v_3945 | ~v_1207;
assign x_5573 = v_3945 | ~v_183;
assign x_5574 = v_3945 | ~v_168;
assign x_5575 = v_3945 | ~v_167;
assign x_5576 = v_3945 | ~v_166;
assign x_5577 = v_3945 | ~v_145;
assign x_5578 = v_3945 | ~v_144;
assign x_5579 = v_3945 | ~v_143;
assign x_5580 = v_3945 | ~v_142;
assign x_5581 = v_3945 | ~v_60;
assign x_5582 = v_3945 | ~v_59;
assign x_5583 = v_3945 | ~v_58;
assign x_5584 = v_3945 | ~v_51;
assign x_5585 = v_3944 | ~v_891;
assign x_5586 = v_3944 | ~v_892;
assign x_5587 = v_3944 | ~v_893;
assign x_5588 = v_3944 | ~v_894;
assign x_5589 = v_3944 | ~v_1157;
assign x_5590 = v_3944 | ~v_1158;
assign x_5591 = v_3944 | ~v_1159;
assign x_5592 = v_3944 | ~v_1160;
assign x_5593 = v_3944 | ~v_761;
assign x_5594 = v_3944 | ~v_3884;
assign x_5595 = v_3944 | ~v_3885;
assign x_5596 = v_3944 | ~v_764;
assign x_5597 = v_3944 | ~v_3886;
assign x_5598 = v_3944 | ~v_3887;
assign x_5599 = v_3944 | ~v_3506;
assign x_5600 = v_3944 | ~v_3507;
assign x_5601 = v_3944 | ~v_3508;
assign x_5602 = v_3944 | ~v_3509;
assign x_5603 = v_3944 | ~v_3522;
assign x_5604 = v_3944 | ~v_3523;
assign x_5605 = v_3944 | ~v_3524;
assign x_5606 = v_3944 | ~v_3525;
assign x_5607 = v_3944 | ~v_3466;
assign x_5608 = v_3944 | ~v_3469;
assign x_5609 = v_3944 | ~v_1199;
assign x_5610 = v_3944 | ~v_1200;
assign x_5611 = v_3944 | ~v_1163;
assign x_5612 = v_3944 | ~v_1164;
assign x_5613 = v_3944 | ~v_897;
assign x_5614 = v_3944 | ~v_898;
assign x_5615 = v_3944 | ~v_1201;
assign x_5616 = v_3944 | ~v_1202;
assign x_5617 = v_3944 | ~v_182;
assign x_5618 = v_3944 | ~v_164;
assign x_5619 = v_3944 | ~v_163;
assign x_5620 = v_3944 | ~v_162;
assign x_5621 = v_3944 | ~v_137;
assign x_5622 = v_3944 | ~v_136;
assign x_5623 = v_3944 | ~v_135;
assign x_5624 = v_3944 | ~v_134;
assign x_5625 = v_3944 | ~v_17;
assign x_5626 = v_3944 | ~v_16;
assign x_5627 = v_3944 | ~v_15;
assign x_5628 = v_3944 | ~v_8;
assign x_5629 = ~v_3942 | ~v_3941 | ~v_3940 | v_3943;
assign x_5630 = v_3942 | ~v_823;
assign x_5631 = v_3942 | ~v_824;
assign x_5632 = v_3942 | ~v_825;
assign x_5633 = v_3942 | ~v_826;
assign x_5634 = v_3942 | ~v_1187;
assign x_5635 = v_3942 | ~v_1188;
assign x_5636 = v_3942 | ~v_1189;
assign x_5637 = v_3942 | ~v_1190;
assign x_5638 = v_3942 | ~v_827;
assign x_5639 = v_3942 | ~v_3894;
assign x_5640 = v_3942 | ~v_3895;
assign x_5641 = v_3942 | ~v_830;
assign x_5642 = v_3942 | ~v_3896;
assign x_5643 = v_3942 | ~v_3897;
assign x_5644 = v_3942 | ~v_3516;
assign x_5645 = v_3942 | ~v_3517;
assign x_5646 = v_3942 | ~v_3518;
assign x_5647 = v_3942 | ~v_3519;
assign x_5648 = v_3942 | ~v_3548;
assign x_5649 = v_3942 | ~v_3549;
assign x_5650 = v_3942 | ~v_3550;
assign x_5651 = v_3942 | ~v_3551;
assign x_5652 = v_3942 | ~v_3496;
assign x_5653 = v_3942 | ~v_3499;
assign x_5654 = v_3942 | ~v_1191;
assign x_5655 = v_3942 | ~v_1192;
assign x_5656 = v_3942 | ~v_1193;
assign x_5657 = v_3942 | ~v_1194;
assign x_5658 = v_3942 | ~v_837;
assign x_5659 = v_3942 | ~v_838;
assign x_5660 = v_3942 | ~v_1195;
assign x_5661 = v_3942 | ~v_1196;
assign x_5662 = v_3942 | ~v_184;
assign x_5663 = v_3942 | ~v_171;
assign x_5664 = v_3942 | ~v_170;
assign x_5665 = v_3942 | ~v_160;
assign x_5666 = v_3942 | ~v_151;
assign x_5667 = v_3942 | ~v_150;
assign x_5668 = v_3942 | ~v_149;
assign x_5669 = v_3942 | ~v_148;
assign x_5670 = v_3942 | ~v_147;
assign x_5671 = v_3942 | ~v_103;
assign x_5672 = v_3942 | ~v_100;
assign x_5673 = v_3942 | ~v_93;
assign x_5674 = v_3941 | ~v_790;
assign x_5675 = v_3941 | ~v_791;
assign x_5676 = v_3941 | ~v_792;
assign x_5677 = v_3941 | ~v_793;
assign x_5678 = v_3941 | ~v_1172;
assign x_5679 = v_3941 | ~v_1173;
assign x_5680 = v_3941 | ~v_1174;
assign x_5681 = v_3941 | ~v_1175;
assign x_5682 = v_3941 | ~v_794;
assign x_5683 = v_3941 | ~v_3889;
assign x_5684 = v_3941 | ~v_3890;
assign x_5685 = v_3941 | ~v_797;
assign x_5686 = v_3941 | ~v_3891;
assign x_5687 = v_3941 | ~v_3892;
assign x_5688 = v_3941 | ~v_3511;
assign x_5689 = v_3941 | ~v_3512;
assign x_5690 = v_3941 | ~v_3513;
assign x_5691 = v_3941 | ~v_3514;
assign x_5692 = v_3941 | ~v_3543;
assign x_5693 = v_3941 | ~v_3544;
assign x_5694 = v_3941 | ~v_3545;
assign x_5695 = v_3941 | ~v_3546;
assign x_5696 = v_3941 | ~v_3481;
assign x_5697 = v_3941 | ~v_3484;
assign x_5698 = v_3941 | ~v_1176;
assign x_5699 = v_3941 | ~v_1177;
assign x_5700 = v_3941 | ~v_1178;
assign x_5701 = v_3941 | ~v_1179;
assign x_5702 = v_3941 | ~v_804;
assign x_5703 = v_3941 | ~v_805;
assign x_5704 = v_3941 | ~v_1180;
assign x_5705 = v_3941 | ~v_1181;
assign x_5706 = v_3941 | ~v_183;
assign x_5707 = v_3941 | ~v_167;
assign x_5708 = v_3941 | ~v_166;
assign x_5709 = v_3941 | ~v_159;
assign x_5710 = v_3941 | ~v_146;
assign x_5711 = v_3941 | ~v_145;
assign x_5712 = v_3941 | ~v_144;
assign x_5713 = v_3941 | ~v_143;
assign x_5714 = v_3941 | ~v_142;
assign x_5715 = v_3941 | ~v_61;
assign x_5716 = v_3941 | ~v_58;
assign x_5717 = v_3941 | ~v_51;
assign x_5718 = v_3940 | ~v_757;
assign x_5719 = v_3940 | ~v_758;
assign x_5720 = v_3940 | ~v_759;
assign x_5721 = v_3940 | ~v_760;
assign x_5722 = v_3940 | ~v_1157;
assign x_5723 = v_3940 | ~v_1158;
assign x_5724 = v_3940 | ~v_1159;
assign x_5725 = v_3940 | ~v_1160;
assign x_5726 = v_3940 | ~v_761;
assign x_5727 = v_3940 | ~v_3884;
assign x_5728 = v_3940 | ~v_3885;
assign x_5729 = v_3940 | ~v_764;
assign x_5730 = v_3940 | ~v_3886;
assign x_5731 = v_3940 | ~v_3887;
assign x_5732 = v_3940 | ~v_3506;
assign x_5733 = v_3940 | ~v_3507;
assign x_5734 = v_3940 | ~v_3508;
assign x_5735 = v_3940 | ~v_3509;
assign x_5736 = v_3940 | ~v_3538;
assign x_5737 = v_3940 | ~v_3539;
assign x_5738 = v_3940 | ~v_3540;
assign x_5739 = v_3940 | ~v_3541;
assign x_5740 = v_3940 | ~v_3466;
assign x_5741 = v_3940 | ~v_3469;
assign x_5742 = v_3940 | ~v_1161;
assign x_5743 = v_3940 | ~v_1162;
assign x_5744 = v_3940 | ~v_1163;
assign x_5745 = v_3940 | ~v_1164;
assign x_5746 = v_3940 | ~v_771;
assign x_5747 = v_3940 | ~v_772;
assign x_5748 = v_3940 | ~v_1165;
assign x_5749 = v_3940 | ~v_1166;
assign x_5750 = v_3940 | ~v_182;
assign x_5751 = v_3940 | ~v_163;
assign x_5752 = v_3940 | ~v_162;
assign x_5753 = v_3940 | ~v_155;
assign x_5754 = v_3940 | ~v_138;
assign x_5755 = v_3940 | ~v_137;
assign x_5756 = v_3940 | ~v_136;
assign x_5757 = v_3940 | ~v_135;
assign x_5758 = v_3940 | ~v_134;
assign x_5759 = v_3940 | ~v_18;
assign x_5760 = v_3940 | ~v_15;
assign x_5761 = v_3940 | ~v_8;
assign x_5762 = ~v_3938 | ~v_3937 | ~v_3936 | v_3939;
assign x_5763 = v_3938 | ~v_969;
assign x_5764 = v_3938 | ~v_970;
assign x_5765 = v_3938 | ~v_971;
assign x_5766 = v_3938 | ~v_972;
assign x_5767 = v_3938 | ~v_827;
assign x_5768 = v_3938 | ~v_3894;
assign x_5769 = v_3938 | ~v_828;
assign x_5770 = v_3938 | ~v_3895;
assign x_5771 = v_3938 | ~v_829;
assign x_5772 = v_3938 | ~v_830;
assign x_5773 = v_3938 | ~v_3896;
assign x_5774 = v_3938 | ~v_831;
assign x_5775 = v_3938 | ~v_3897;
assign x_5776 = v_3938 | ~v_832;
assign x_5777 = v_3938 | ~v_3494;
assign x_5778 = v_3938 | ~v_3495;
assign x_5779 = v_3938 | ~v_3496;
assign x_5780 = v_3938 | ~v_3497;
assign x_5781 = v_3938 | ~v_3498;
assign x_5782 = v_3938 | ~v_3499;
assign x_5783 = v_3938 | ~v_3500;
assign x_5784 = v_3938 | ~v_3501;
assign x_5785 = v_3938 | ~v_1147;
assign x_5786 = v_3938 | ~v_1148;
assign x_5787 = v_3938 | ~v_975;
assign x_5788 = v_3938 | ~v_976;
assign x_5789 = v_3938 | ~v_839;
assign x_5790 = v_3938 | ~v_840;
assign x_5791 = v_3938 | ~v_1149;
assign x_5792 = v_3938 | ~v_1150;
assign x_5793 = v_3938 | ~v_3502;
assign x_5794 = v_3938 | ~v_3503;
assign x_5795 = v_3938 | ~v_184;
assign x_5796 = v_3938 | ~v_169;
assign x_5797 = v_3938 | ~v_150;
assign x_5798 = v_3938 | ~v_149;
assign x_5799 = v_3938 | ~v_147;
assign x_5800 = v_3938 | ~v_103;
assign x_5801 = v_3938 | ~v_102;
assign x_5802 = v_3938 | ~v_101;
assign x_5803 = v_3938 | ~v_100;
assign x_5804 = v_3938 | ~v_98;
assign x_5805 = v_3938 | ~v_96;
assign x_5806 = v_3938 | ~v_94;
assign x_5807 = v_3937 | ~v_954;
assign x_5808 = v_3937 | ~v_955;
assign x_5809 = v_3937 | ~v_956;
assign x_5810 = v_3937 | ~v_957;
assign x_5811 = v_3937 | ~v_794;
assign x_5812 = v_3937 | ~v_3889;
assign x_5813 = v_3937 | ~v_795;
assign x_5814 = v_3937 | ~v_3890;
assign x_5815 = v_3937 | ~v_796;
assign x_5816 = v_3937 | ~v_797;
assign x_5817 = v_3937 | ~v_3891;
assign x_5818 = v_3937 | ~v_798;
assign x_5819 = v_3937 | ~v_3892;
assign x_5820 = v_3937 | ~v_799;
assign x_5821 = v_3937 | ~v_3479;
assign x_5822 = v_3937 | ~v_3480;
assign x_5823 = v_3937 | ~v_3481;
assign x_5824 = v_3937 | ~v_3482;
assign x_5825 = v_3937 | ~v_3483;
assign x_5826 = v_3937 | ~v_3484;
assign x_5827 = v_3937 | ~v_3485;
assign x_5828 = v_3937 | ~v_1142;
assign x_5829 = v_3937 | ~v_1143;
assign x_5830 = v_3937 | ~v_960;
assign x_5831 = v_3937 | ~v_961;
assign x_5832 = v_3937 | ~v_806;
assign x_5833 = v_3937 | ~v_807;
assign x_5834 = v_3937 | ~v_3486;
assign x_5835 = v_3937 | ~v_1144;
assign x_5836 = v_3937 | ~v_1145;
assign x_5837 = v_3937 | ~v_3487;
assign x_5838 = v_3937 | ~v_3488;
assign x_5839 = v_3937 | ~v_183;
assign x_5840 = v_3937 | ~v_165;
assign x_5841 = v_3937 | ~v_145;
assign x_5842 = v_3937 | ~v_144;
assign x_5843 = v_3937 | ~v_142;
assign x_5844 = v_3937 | ~v_61;
assign x_5845 = v_3937 | ~v_60;
assign x_5846 = v_3937 | ~v_59;
assign x_5847 = v_3937 | ~v_58;
assign x_5848 = v_3937 | ~v_56;
assign x_5849 = v_3937 | ~v_54;
assign x_5850 = v_3937 | ~v_52;
assign x_5851 = v_3936 | ~v_939;
assign x_5852 = v_3936 | ~v_940;
assign x_5853 = v_3936 | ~v_941;
assign x_5854 = v_3936 | ~v_942;
assign x_5855 = v_3936 | ~v_761;
assign x_5856 = v_3936 | ~v_3884;
assign x_5857 = v_3936 | ~v_762;
assign x_5858 = v_3936 | ~v_3885;
assign x_5859 = v_3936 | ~v_763;
assign x_5860 = v_3936 | ~v_764;
assign x_5861 = v_3936 | ~v_3886;
assign x_5862 = v_3936 | ~v_765;
assign x_5863 = v_3936 | ~v_3887;
assign x_5864 = v_3936 | ~v_766;
assign x_5865 = v_3936 | ~v_3464;
assign x_5866 = v_3936 | ~v_3465;
assign x_5867 = v_3936 | ~v_3466;
assign x_5868 = v_3936 | ~v_3467;
assign x_5869 = v_3936 | ~v_3468;
assign x_5870 = v_3936 | ~v_3469;
assign x_5871 = v_3936 | ~v_3470;
assign x_5872 = v_3936 | ~v_1137;
assign x_5873 = v_3936 | ~v_1138;
assign x_5874 = v_3936 | ~v_945;
assign x_5875 = v_3936 | ~v_946;
assign x_5876 = v_3936 | ~v_773;
assign x_5877 = v_3936 | ~v_774;
assign x_5878 = v_3936 | ~v_1139;
assign x_5879 = v_3936 | ~v_1140;
assign x_5880 = v_3936 | ~v_3471;
assign x_5881 = v_3936 | ~v_3472;
assign x_5882 = v_3936 | ~v_182;
assign x_5883 = v_3936 | ~v_161;
assign x_5884 = v_3936 | ~v_137;
assign x_5885 = v_3936 | ~v_3473;
assign x_5886 = v_3936 | ~v_136;
assign x_5887 = v_3936 | ~v_134;
assign x_5888 = v_3936 | ~v_18;
assign x_5889 = v_3936 | ~v_17;
assign x_5890 = v_3936 | ~v_16;
assign x_5891 = v_3936 | ~v_15;
assign x_5892 = v_3936 | ~v_13;
assign x_5893 = v_3936 | ~v_11;
assign x_5894 = v_3936 | ~v_9;
assign x_5895 = ~v_3934 | ~v_3933 | ~v_3932 | v_3935;
assign x_5896 = v_3934 | ~v_1077;
assign x_5897 = v_3934 | ~v_1078;
assign x_5898 = v_3934 | ~v_1079;
assign x_5899 = v_3934 | ~v_1080;
assign x_5900 = v_3934 | ~v_827;
assign x_5901 = v_3934 | ~v_3894;
assign x_5902 = v_3934 | ~v_1015;
assign x_5903 = v_3934 | ~v_3895;
assign x_5904 = v_3934 | ~v_1016;
assign x_5905 = v_3934 | ~v_830;
assign x_5906 = v_3934 | ~v_3896;
assign x_5907 = v_3934 | ~v_1017;
assign x_5908 = v_3934 | ~v_3897;
assign x_5909 = v_3934 | ~v_1018;
assign x_5910 = v_3934 | ~v_3584;
assign x_5911 = v_3934 | ~v_3585;
assign x_5912 = v_3934 | ~v_3586;
assign x_5913 = v_3934 | ~v_3587;
assign x_5914 = v_3934 | ~v_3496;
assign x_5915 = v_3934 | ~v_3564;
assign x_5916 = v_3934 | ~v_3565;
assign x_5917 = v_3934 | ~v_3499;
assign x_5918 = v_3934 | ~v_3566;
assign x_5919 = v_3934 | ~v_3567;
assign x_5920 = v_3934 | ~v_1085;
assign x_5921 = v_3934 | ~v_1131;
assign x_5922 = v_3934 | ~v_1132;
assign x_5923 = v_3934 | ~v_1086;
assign x_5924 = v_3934 | ~v_1133;
assign x_5925 = v_3934 | ~v_1134;
assign x_5926 = v_3934 | ~v_1023;
assign x_5927 = v_3934 | ~v_1024;
assign x_5928 = v_3934 | ~v_184;
assign x_5929 = v_3934 | ~v_172;
assign x_5930 = v_3934 | ~v_171;
assign x_5931 = v_3934 | ~v_170;
assign x_5932 = v_3934 | ~v_169;
assign x_5933 = v_3934 | ~v_148;
assign x_5934 = v_3934 | ~v_147;
assign x_5935 = v_3934 | ~v_102;
assign x_5936 = v_3934 | ~v_101;
assign x_5937 = v_3934 | ~v_100;
assign x_5938 = v_3934 | ~v_99;
assign x_5939 = v_3934 | ~v_97;
assign x_5940 = v_3933 | ~v_1062;
assign x_5941 = v_3933 | ~v_1063;
assign x_5942 = v_3933 | ~v_1064;
assign x_5943 = v_3933 | ~v_1065;
assign x_5944 = v_3933 | ~v_794;
assign x_5945 = v_3933 | ~v_3889;
assign x_5946 = v_3933 | ~v_1000;
assign x_5947 = v_3933 | ~v_3890;
assign x_5948 = v_3933 | ~v_1001;
assign x_5949 = v_3933 | ~v_797;
assign x_5950 = v_3933 | ~v_3891;
assign x_5951 = v_3933 | ~v_1002;
assign x_5952 = v_3933 | ~v_3892;
assign x_5953 = v_3933 | ~v_1003;
assign x_5954 = v_3933 | ~v_3579;
assign x_5955 = v_3933 | ~v_3580;
assign x_5956 = v_3933 | ~v_3581;
assign x_5957 = v_3933 | ~v_3582;
assign x_5958 = v_3933 | ~v_3481;
assign x_5959 = v_3933 | ~v_3559;
assign x_5960 = v_3933 | ~v_3560;
assign x_5961 = v_3933 | ~v_3484;
assign x_5962 = v_3933 | ~v_1070;
assign x_5963 = v_3933 | ~v_1126;
assign x_5964 = v_3933 | ~v_1127;
assign x_5965 = v_3933 | ~v_1071;
assign x_5966 = v_3933 | ~v_1128;
assign x_5967 = v_3933 | ~v_1129;
assign x_5968 = v_3933 | ~v_1008;
assign x_5969 = v_3933 | ~v_1009;
assign x_5970 = v_3933 | ~v_3561;
assign x_5971 = v_3933 | ~v_3562;
assign x_5972 = v_3933 | ~v_183;
assign x_5973 = v_3933 | ~v_168;
assign x_5974 = v_3933 | ~v_167;
assign x_5975 = v_3933 | ~v_166;
assign x_5976 = v_3933 | ~v_165;
assign x_5977 = v_3933 | ~v_143;
assign x_5978 = v_3933 | ~v_142;
assign x_5979 = v_3933 | ~v_60;
assign x_5980 = v_3933 | ~v_59;
assign x_5981 = v_3933 | ~v_58;
assign x_5982 = v_3933 | ~v_57;
assign x_5983 = v_3933 | ~v_55;
assign x_5984 = v_3932 | ~v_1047;
assign x_5985 = v_3932 | ~v_1048;
assign x_5986 = v_3932 | ~v_1049;
assign x_5987 = v_3932 | ~v_1050;
assign x_5988 = v_3932 | ~v_761;
assign x_5989 = v_3932 | ~v_3884;
assign x_5990 = v_3932 | ~v_985;
assign x_5991 = v_3932 | ~v_3885;
assign x_5992 = v_3932 | ~v_986;
assign x_5993 = v_3932 | ~v_764;
assign x_5994 = v_3932 | ~v_3886;
assign x_5995 = v_3932 | ~v_987;
assign x_5996 = v_3932 | ~v_3887;
assign x_5997 = v_3932 | ~v_988;
assign x_5998 = v_3932 | ~v_3574;
assign x_5999 = v_3932 | ~v_3575;
assign x_6000 = v_3932 | ~v_3576;
assign x_6001 = v_3932 | ~v_3577;
assign x_6002 = v_3932 | ~v_3466;
assign x_6003 = v_3932 | ~v_3554;
assign x_6004 = v_3932 | ~v_3555;
assign x_6005 = v_3932 | ~v_3469;
assign x_6006 = v_3932 | ~v_3556;
assign x_6007 = v_3932 | ~v_3557;
assign x_6008 = v_3932 | ~v_1055;
assign x_6009 = v_3932 | ~v_1121;
assign x_6010 = v_3932 | ~v_1122;
assign x_6011 = v_3932 | ~v_1056;
assign x_6012 = v_3932 | ~v_1123;
assign x_6013 = v_3932 | ~v_1124;
assign x_6014 = v_3932 | ~v_182;
assign x_6015 = v_3932 | ~v_164;
assign x_6016 = v_3932 | ~v_163;
assign x_6017 = v_3932 | ~v_162;
assign x_6018 = v_3932 | ~v_161;
assign x_6019 = v_3932 | ~v_135;
assign x_6020 = v_3932 | ~v_134;
assign x_6021 = v_3932 | ~v_993;
assign x_6022 = v_3932 | ~v_994;
assign x_6023 = v_3932 | ~v_17;
assign x_6024 = v_3932 | ~v_16;
assign x_6025 = v_3932 | ~v_15;
assign x_6026 = v_3932 | ~v_14;
assign x_6027 = v_3932 | ~v_12;
assign x_6028 = ~v_3930 | ~v_3929 | ~v_3928 | v_3931;
assign x_6029 = v_3930 | ~v_1077;
assign x_6030 = v_3930 | ~v_1078;
assign x_6031 = v_3930 | ~v_1079;
assign x_6032 = v_3930 | ~v_1080;
assign x_6033 = v_3930 | ~v_969;
assign x_6034 = v_3930 | ~v_970;
assign x_6035 = v_3930 | ~v_971;
assign x_6036 = v_3930 | ~v_972;
assign x_6037 = v_3930 | ~v_827;
assign x_6038 = v_3930 | ~v_3894;
assign x_6039 = v_3930 | ~v_3895;
assign x_6040 = v_3930 | ~v_830;
assign x_6041 = v_3930 | ~v_3896;
assign x_6042 = v_3930 | ~v_3897;
assign x_6043 = v_3930 | ~v_3494;
assign x_6044 = v_3930 | ~v_3495;
assign x_6045 = v_3930 | ~v_3584;
assign x_6046 = v_3930 | ~v_3585;
assign x_6047 = v_3930 | ~v_3586;
assign x_6048 = v_3930 | ~v_3587;
assign x_6049 = v_3930 | ~v_3496;
assign x_6050 = v_3930 | ~v_3499;
assign x_6051 = v_3930 | ~v_975;
assign x_6052 = v_3930 | ~v_976;
assign x_6053 = v_3930 | ~v_1115;
assign x_6054 = v_3930 | ~v_1116;
assign x_6055 = v_3930 | ~v_1085;
assign x_6056 = v_3930 | ~v_1086;
assign x_6057 = v_3930 | ~v_1117;
assign x_6058 = v_3930 | ~v_1118;
assign x_6059 = v_3930 | ~v_3502;
assign x_6060 = v_3930 | ~v_3503;
assign x_6061 = v_3930 | ~v_184;
assign x_6062 = v_3930 | ~v_171;
assign x_6063 = v_3930 | ~v_170;
assign x_6064 = v_3930 | ~v_169;
assign x_6065 = v_3930 | ~v_151;
assign x_6066 = v_3930 | ~v_150;
assign x_6067 = v_3930 | ~v_149;
assign x_6068 = v_3930 | ~v_147;
assign x_6069 = v_3930 | ~v_103;
assign x_6070 = v_3930 | ~v_101;
assign x_6071 = v_3930 | ~v_100;
assign x_6072 = v_3930 | ~v_96;
assign x_6073 = v_3929 | ~v_1062;
assign x_6074 = v_3929 | ~v_1063;
assign x_6075 = v_3929 | ~v_1064;
assign x_6076 = v_3929 | ~v_1065;
assign x_6077 = v_3929 | ~v_954;
assign x_6078 = v_3929 | ~v_955;
assign x_6079 = v_3929 | ~v_956;
assign x_6080 = v_3929 | ~v_957;
assign x_6081 = v_3929 | ~v_794;
assign x_6082 = v_3929 | ~v_3889;
assign x_6083 = v_3929 | ~v_3890;
assign x_6084 = v_3929 | ~v_797;
assign x_6085 = v_3929 | ~v_3891;
assign x_6086 = v_3929 | ~v_3892;
assign x_6087 = v_3929 | ~v_3479;
assign x_6088 = v_3929 | ~v_3480;
assign x_6089 = v_3929 | ~v_3579;
assign x_6090 = v_3929 | ~v_3580;
assign x_6091 = v_3929 | ~v_3581;
assign x_6092 = v_3929 | ~v_3582;
assign x_6093 = v_3929 | ~v_3481;
assign x_6094 = v_3929 | ~v_3484;
assign x_6095 = v_3929 | ~v_960;
assign x_6096 = v_3929 | ~v_961;
assign x_6097 = v_3929 | ~v_1110;
assign x_6098 = v_3929 | ~v_1111;
assign x_6099 = v_3929 | ~v_1070;
assign x_6100 = v_3929 | ~v_1071;
assign x_6101 = v_3929 | ~v_1112;
assign x_6102 = v_3929 | ~v_1113;
assign x_6103 = v_3929 | ~v_3487;
assign x_6104 = v_3929 | ~v_3488;
assign x_6105 = v_3929 | ~v_183;
assign x_6106 = v_3929 | ~v_167;
assign x_6107 = v_3929 | ~v_166;
assign x_6108 = v_3929 | ~v_165;
assign x_6109 = v_3929 | ~v_146;
assign x_6110 = v_3929 | ~v_145;
assign x_6111 = v_3929 | ~v_144;
assign x_6112 = v_3929 | ~v_142;
assign x_6113 = v_3929 | ~v_61;
assign x_6114 = v_3929 | ~v_59;
assign x_6115 = v_3929 | ~v_58;
assign x_6116 = v_3929 | ~v_54;
assign x_6117 = v_3928 | ~v_1047;
assign x_6118 = v_3928 | ~v_1048;
assign x_6119 = v_3928 | ~v_1049;
assign x_6120 = v_3928 | ~v_1050;
assign x_6121 = v_3928 | ~v_939;
assign x_6122 = v_3928 | ~v_940;
assign x_6123 = v_3928 | ~v_941;
assign x_6124 = v_3928 | ~v_942;
assign x_6125 = v_3928 | ~v_761;
assign x_6126 = v_3928 | ~v_3884;
assign x_6127 = v_3928 | ~v_3885;
assign x_6128 = v_3928 | ~v_764;
assign x_6129 = v_3928 | ~v_3886;
assign x_6130 = v_3928 | ~v_3887;
assign x_6131 = v_3928 | ~v_3464;
assign x_6132 = v_3928 | ~v_3465;
assign x_6133 = v_3928 | ~v_3574;
assign x_6134 = v_3928 | ~v_3575;
assign x_6135 = v_3928 | ~v_3576;
assign x_6136 = v_3928 | ~v_3577;
assign x_6137 = v_3928 | ~v_3466;
assign x_6138 = v_3928 | ~v_3469;
assign x_6139 = v_3928 | ~v_945;
assign x_6140 = v_3928 | ~v_946;
assign x_6141 = v_3928 | ~v_1105;
assign x_6142 = v_3928 | ~v_1106;
assign x_6143 = v_3928 | ~v_1055;
assign x_6144 = v_3928 | ~v_1056;
assign x_6145 = v_3928 | ~v_1107;
assign x_6146 = v_3928 | ~v_1108;
assign x_6147 = v_3928 | ~v_3471;
assign x_6148 = v_3928 | ~v_3472;
assign x_6149 = v_3928 | ~v_182;
assign x_6150 = v_3928 | ~v_163;
assign x_6151 = v_3928 | ~v_162;
assign x_6152 = v_3928 | ~v_161;
assign x_6153 = v_3928 | ~v_138;
assign x_6154 = v_3928 | ~v_137;
assign x_6155 = v_3928 | ~v_136;
assign x_6156 = v_3928 | ~v_134;
assign x_6157 = v_3928 | ~v_18;
assign x_6158 = v_3928 | ~v_16;
assign x_6159 = v_3928 | ~v_15;
assign x_6160 = v_3928 | ~v_11;
assign x_6161 = ~v_3926 | ~v_3925 | ~v_3924 | v_3927;
assign x_6162 = v_3926 | ~v_1077;
assign x_6163 = v_3926 | ~v_1078;
assign x_6164 = v_3926 | ~v_1079;
assign x_6165 = v_3926 | ~v_1080;
assign x_6166 = v_3926 | ~v_921;
assign x_6167 = v_3926 | ~v_922;
assign x_6168 = v_3926 | ~v_923;
assign x_6169 = v_3926 | ~v_924;
assign x_6170 = v_3926 | ~v_827;
assign x_6171 = v_3926 | ~v_3894;
assign x_6172 = v_3926 | ~v_3895;
assign x_6173 = v_3926 | ~v_830;
assign x_6174 = v_3926 | ~v_3896;
assign x_6175 = v_3926 | ~v_3897;
assign x_6176 = v_3926 | ~v_3532;
assign x_6177 = v_3926 | ~v_3533;
assign x_6178 = v_3926 | ~v_3534;
assign x_6179 = v_3926 | ~v_3535;
assign x_6180 = v_3926 | ~v_3584;
assign x_6181 = v_3926 | ~v_3585;
assign x_6182 = v_3926 | ~v_3586;
assign x_6183 = v_3926 | ~v_3587;
assign x_6184 = v_3926 | ~v_3496;
assign x_6185 = v_3926 | ~v_3499;
assign x_6186 = v_3926 | ~v_927;
assign x_6187 = v_3926 | ~v_928;
assign x_6188 = v_3926 | ~v_1099;
assign x_6189 = v_3926 | ~v_1100;
assign x_6190 = v_3926 | ~v_1101;
assign x_6191 = v_3926 | ~v_1102;
assign x_6192 = v_3926 | ~v_1085;
assign x_6193 = v_3926 | ~v_1086;
assign x_6194 = v_3926 | ~v_184;
assign x_6195 = v_3926 | ~v_171;
assign x_6196 = v_3926 | ~v_170;
assign x_6197 = v_3926 | ~v_169;
assign x_6198 = v_3926 | ~v_150;
assign x_6199 = v_3926 | ~v_149;
assign x_6200 = v_3926 | ~v_148;
assign x_6201 = v_3926 | ~v_103;
assign x_6202 = v_3926 | ~v_102;
assign x_6203 = v_3926 | ~v_101;
assign x_6204 = v_3926 | ~v_100;
assign x_6205 = v_3926 | ~v_95;
assign x_6206 = v_3925 | ~v_1062;
assign x_6207 = v_3925 | ~v_1063;
assign x_6208 = v_3925 | ~v_1064;
assign x_6209 = v_3925 | ~v_1065;
assign x_6210 = v_3925 | ~v_906;
assign x_6211 = v_3925 | ~v_907;
assign x_6212 = v_3925 | ~v_908;
assign x_6213 = v_3925 | ~v_909;
assign x_6214 = v_3925 | ~v_794;
assign x_6215 = v_3925 | ~v_3889;
assign x_6216 = v_3925 | ~v_3890;
assign x_6217 = v_3925 | ~v_797;
assign x_6218 = v_3925 | ~v_3891;
assign x_6219 = v_3925 | ~v_3892;
assign x_6220 = v_3925 | ~v_3527;
assign x_6221 = v_3925 | ~v_3528;
assign x_6222 = v_3925 | ~v_3529;
assign x_6223 = v_3925 | ~v_3530;
assign x_6224 = v_3925 | ~v_3579;
assign x_6225 = v_3925 | ~v_3580;
assign x_6226 = v_3925 | ~v_3581;
assign x_6227 = v_3925 | ~v_3582;
assign x_6228 = v_3925 | ~v_3481;
assign x_6229 = v_3925 | ~v_3484;
assign x_6230 = v_3925 | ~v_912;
assign x_6231 = v_3925 | ~v_913;
assign x_6232 = v_3925 | ~v_1094;
assign x_6233 = v_3925 | ~v_1095;
assign x_6234 = v_3925 | ~v_1096;
assign x_6235 = v_3925 | ~v_1097;
assign x_6236 = v_3925 | ~v_1070;
assign x_6237 = v_3925 | ~v_1071;
assign x_6238 = v_3925 | ~v_183;
assign x_6239 = v_3925 | ~v_167;
assign x_6240 = v_3925 | ~v_166;
assign x_6241 = v_3925 | ~v_165;
assign x_6242 = v_3925 | ~v_145;
assign x_6243 = v_3925 | ~v_144;
assign x_6244 = v_3925 | ~v_143;
assign x_6245 = v_3925 | ~v_61;
assign x_6246 = v_3925 | ~v_60;
assign x_6247 = v_3925 | ~v_59;
assign x_6248 = v_3925 | ~v_58;
assign x_6249 = v_3925 | ~v_53;
assign x_6250 = v_3924 | ~v_1047;
assign x_6251 = v_3924 | ~v_1048;
assign x_6252 = v_3924 | ~v_1049;
assign x_6253 = v_3924 | ~v_1050;
assign x_6254 = v_3924 | ~v_891;
assign x_6255 = v_3924 | ~v_892;
assign x_6256 = v_3924 | ~v_893;
assign x_6257 = v_3924 | ~v_894;
assign x_6258 = v_3924 | ~v_761;
assign x_6259 = v_3924 | ~v_3884;
assign x_6260 = v_3924 | ~v_3885;
assign x_6261 = v_3924 | ~v_764;
assign x_6262 = v_3924 | ~v_3886;
assign x_6263 = v_3924 | ~v_3887;
assign x_6264 = v_3924 | ~v_3522;
assign x_6265 = v_3924 | ~v_3523;
assign x_6266 = v_3924 | ~v_3524;
assign x_6267 = v_3924 | ~v_3525;
assign x_6268 = v_3924 | ~v_3574;
assign x_6269 = v_3924 | ~v_3575;
assign x_6270 = v_3924 | ~v_3576;
assign x_6271 = v_3924 | ~v_3577;
assign x_6272 = v_3924 | ~v_3466;
assign x_6273 = v_3924 | ~v_3469;
assign x_6274 = v_3924 | ~v_897;
assign x_6275 = v_3924 | ~v_898;
assign x_6276 = v_3924 | ~v_1089;
assign x_6277 = v_3924 | ~v_1090;
assign x_6278 = v_3924 | ~v_1091;
assign x_6279 = v_3924 | ~v_1092;
assign x_6280 = v_3924 | ~v_1055;
assign x_6281 = v_3924 | ~v_1056;
assign x_6282 = v_3924 | ~v_182;
assign x_6283 = v_3924 | ~v_163;
assign x_6284 = v_3924 | ~v_162;
assign x_6285 = v_3924 | ~v_161;
assign x_6286 = v_3924 | ~v_137;
assign x_6287 = v_3924 | ~v_136;
assign x_6288 = v_3924 | ~v_135;
assign x_6289 = v_3924 | ~v_18;
assign x_6290 = v_3924 | ~v_17;
assign x_6291 = v_3924 | ~v_16;
assign x_6292 = v_3924 | ~v_15;
assign x_6293 = v_3924 | ~v_10;
assign x_6294 = ~v_3922 | ~v_3921 | ~v_3920 | v_3923;
assign x_6295 = v_3922 | ~v_1077;
assign x_6296 = v_3922 | ~v_1078;
assign x_6297 = v_3922 | ~v_1079;
assign x_6298 = v_3922 | ~v_1080;
assign x_6299 = v_3922 | ~v_823;
assign x_6300 = v_3922 | ~v_824;
assign x_6301 = v_3922 | ~v_825;
assign x_6302 = v_3922 | ~v_826;
assign x_6303 = v_3922 | ~v_827;
assign x_6304 = v_3922 | ~v_3894;
assign x_6305 = v_3922 | ~v_3895;
assign x_6306 = v_3922 | ~v_830;
assign x_6307 = v_3922 | ~v_3896;
assign x_6308 = v_3922 | ~v_3897;
assign x_6309 = v_3922 | ~v_3548;
assign x_6310 = v_3922 | ~v_3549;
assign x_6311 = v_3922 | ~v_3550;
assign x_6312 = v_3922 | ~v_3551;
assign x_6313 = v_3922 | ~v_3584;
assign x_6314 = v_3922 | ~v_3585;
assign x_6315 = v_3922 | ~v_3586;
assign x_6316 = v_3922 | ~v_3587;
assign x_6317 = v_3922 | ~v_3496;
assign x_6318 = v_3922 | ~v_3499;
assign x_6319 = v_3922 | ~v_837;
assign x_6320 = v_3922 | ~v_838;
assign x_6321 = v_3922 | ~v_1081;
assign x_6322 = v_3922 | ~v_1082;
assign x_6323 = v_3922 | ~v_1083;
assign x_6324 = v_3922 | ~v_1084;
assign x_6325 = v_3922 | ~v_1085;
assign x_6326 = v_3922 | ~v_1086;
assign x_6327 = v_3922 | ~v_184;
assign x_6328 = v_3922 | ~v_171;
assign x_6329 = v_3922 | ~v_170;
assign x_6330 = v_3922 | ~v_169;
assign x_6331 = v_3922 | ~v_160;
assign x_6332 = v_3922 | ~v_150;
assign x_6333 = v_3922 | ~v_149;
assign x_6334 = v_3922 | ~v_148;
assign x_6335 = v_3922 | ~v_147;
assign x_6336 = v_3922 | ~v_103;
assign x_6337 = v_3922 | ~v_102;
assign x_6338 = v_3922 | ~v_100;
assign x_6339 = v_3921 | ~v_1062;
assign x_6340 = v_3921 | ~v_1063;
assign x_6341 = v_3921 | ~v_1064;
assign x_6342 = v_3921 | ~v_1065;
assign x_6343 = v_3921 | ~v_790;
assign x_6344 = v_3921 | ~v_791;
assign x_6345 = v_3921 | ~v_792;
assign x_6346 = v_3921 | ~v_793;
assign x_6347 = v_3921 | ~v_794;
assign x_6348 = v_3921 | ~v_3889;
assign x_6349 = v_3921 | ~v_3890;
assign x_6350 = v_3921 | ~v_797;
assign x_6351 = v_3921 | ~v_3891;
assign x_6352 = v_3921 | ~v_3892;
assign x_6353 = v_3921 | ~v_3543;
assign x_6354 = v_3921 | ~v_3544;
assign x_6355 = v_3921 | ~v_3545;
assign x_6356 = v_3921 | ~v_3546;
assign x_6357 = v_3921 | ~v_3579;
assign x_6358 = v_3921 | ~v_3580;
assign x_6359 = v_3921 | ~v_3581;
assign x_6360 = v_3921 | ~v_3582;
assign x_6361 = v_3921 | ~v_3481;
assign x_6362 = v_3921 | ~v_3484;
assign x_6363 = v_3921 | ~v_804;
assign x_6364 = v_3921 | ~v_805;
assign x_6365 = v_3921 | ~v_1066;
assign x_6366 = v_3921 | ~v_1067;
assign x_6367 = v_3921 | ~v_1068;
assign x_6368 = v_3921 | ~v_1069;
assign x_6369 = v_3921 | ~v_1070;
assign x_6370 = v_3921 | ~v_1071;
assign x_6371 = v_3921 | ~v_183;
assign x_6372 = v_3921 | ~v_167;
assign x_6373 = v_3921 | ~v_166;
assign x_6374 = v_3921 | ~v_165;
assign x_6375 = v_3921 | ~v_159;
assign x_6376 = v_3921 | ~v_145;
assign x_6377 = v_3921 | ~v_144;
assign x_6378 = v_3921 | ~v_143;
assign x_6379 = v_3921 | ~v_142;
assign x_6380 = v_3921 | ~v_61;
assign x_6381 = v_3921 | ~v_60;
assign x_6382 = v_3921 | ~v_58;
assign x_6383 = v_3920 | ~v_1047;
assign x_6384 = v_3920 | ~v_1048;
assign x_6385 = v_3920 | ~v_1049;
assign x_6386 = v_3920 | ~v_1050;
assign x_6387 = v_3920 | ~v_757;
assign x_6388 = v_3920 | ~v_758;
assign x_6389 = v_3920 | ~v_759;
assign x_6390 = v_3920 | ~v_760;
assign x_6391 = v_3920 | ~v_761;
assign x_6392 = v_3920 | ~v_3884;
assign x_6393 = v_3920 | ~v_3885;
assign x_6394 = v_3920 | ~v_764;
assign x_6395 = v_3920 | ~v_3886;
assign x_6396 = v_3920 | ~v_3887;
assign x_6397 = v_3920 | ~v_3538;
assign x_6398 = v_3920 | ~v_3539;
assign x_6399 = v_3920 | ~v_3540;
assign x_6400 = v_3920 | ~v_3541;
assign x_6401 = v_3920 | ~v_3574;
assign x_6402 = v_3920 | ~v_3575;
assign x_6403 = v_3920 | ~v_3576;
assign x_6404 = v_3920 | ~v_3577;
assign x_6405 = v_3920 | ~v_3466;
assign x_6406 = v_3920 | ~v_3469;
assign x_6407 = v_3920 | ~v_771;
assign x_6408 = v_3920 | ~v_772;
assign x_6409 = v_3920 | ~v_1051;
assign x_6410 = v_3920 | ~v_1052;
assign x_6411 = v_3920 | ~v_1053;
assign x_6412 = v_3920 | ~v_1054;
assign x_6413 = v_3920 | ~v_1055;
assign x_6414 = v_3920 | ~v_1056;
assign x_6415 = v_3920 | ~v_182;
assign x_6416 = v_3920 | ~v_163;
assign x_6417 = v_3920 | ~v_162;
assign x_6418 = v_3920 | ~v_161;
assign x_6419 = v_3920 | ~v_155;
assign x_6420 = v_3920 | ~v_137;
assign x_6421 = v_3920 | ~v_136;
assign x_6422 = v_3920 | ~v_135;
assign x_6423 = v_3920 | ~v_134;
assign x_6424 = v_3920 | ~v_18;
assign x_6425 = v_3920 | ~v_17;
assign x_6426 = v_3920 | ~v_15;
assign x_6427 = ~v_3918 | ~v_3917 | ~v_3916 | v_3919;
assign x_6428 = v_3918 | ~v_921;
assign x_6429 = v_3918 | ~v_922;
assign x_6430 = v_3918 | ~v_923;
assign x_6431 = v_3918 | ~v_924;
assign x_6432 = v_3918 | ~v_827;
assign x_6433 = v_3918 | ~v_3894;
assign x_6434 = v_3918 | ~v_828;
assign x_6435 = v_3918 | ~v_3895;
assign x_6436 = v_3918 | ~v_829;
assign x_6437 = v_3918 | ~v_830;
assign x_6438 = v_3918 | ~v_3896;
assign x_6439 = v_3918 | ~v_831;
assign x_6440 = v_3918 | ~v_3897;
assign x_6441 = v_3918 | ~v_832;
assign x_6442 = v_3918 | ~v_3532;
assign x_6443 = v_3918 | ~v_3533;
assign x_6444 = v_3918 | ~v_3534;
assign x_6445 = v_3918 | ~v_3535;
assign x_6446 = v_3918 | ~v_3496;
assign x_6447 = v_3918 | ~v_3497;
assign x_6448 = v_3918 | ~v_3498;
assign x_6449 = v_3918 | ~v_3499;
assign x_6450 = v_3918 | ~v_3500;
assign x_6451 = v_3918 | ~v_3501;
assign x_6452 = v_3918 | ~v_1037;
assign x_6453 = v_3918 | ~v_1038;
assign x_6454 = v_3918 | ~v_1039;
assign x_6455 = v_3918 | ~v_1040;
assign x_6456 = v_3918 | ~v_927;
assign x_6457 = v_3918 | ~v_928;
assign x_6458 = v_3918 | ~v_839;
assign x_6459 = v_3918 | ~v_840;
assign x_6460 = v_3918 | ~v_184;
assign x_6461 = v_3918 | ~v_169;
assign x_6462 = v_3918 | ~v_151;
assign x_6463 = v_3918 | ~v_150;
assign x_6464 = v_3918 | ~v_149;
assign x_6465 = v_3918 | ~v_148;
assign x_6466 = v_3918 | ~v_147;
assign x_6467 = v_3918 | ~v_103;
assign x_6468 = v_3918 | ~v_101;
assign x_6469 = v_3918 | ~v_100;
assign x_6470 = v_3918 | ~v_98;
assign x_6471 = v_3918 | ~v_94;
assign x_6472 = v_3917 | ~v_906;
assign x_6473 = v_3917 | ~v_907;
assign x_6474 = v_3917 | ~v_908;
assign x_6475 = v_3917 | ~v_909;
assign x_6476 = v_3917 | ~v_794;
assign x_6477 = v_3917 | ~v_3889;
assign x_6478 = v_3917 | ~v_795;
assign x_6479 = v_3917 | ~v_3890;
assign x_6480 = v_3917 | ~v_796;
assign x_6481 = v_3917 | ~v_797;
assign x_6482 = v_3917 | ~v_3891;
assign x_6483 = v_3917 | ~v_798;
assign x_6484 = v_3917 | ~v_3892;
assign x_6485 = v_3917 | ~v_799;
assign x_6486 = v_3917 | ~v_3527;
assign x_6487 = v_3917 | ~v_3528;
assign x_6488 = v_3917 | ~v_3529;
assign x_6489 = v_3917 | ~v_3530;
assign x_6490 = v_3917 | ~v_3481;
assign x_6491 = v_3917 | ~v_3482;
assign x_6492 = v_3917 | ~v_3483;
assign x_6493 = v_3917 | ~v_3484;
assign x_6494 = v_3917 | ~v_3485;
assign x_6495 = v_3917 | ~v_1032;
assign x_6496 = v_3917 | ~v_1033;
assign x_6497 = v_3917 | ~v_1034;
assign x_6498 = v_3917 | ~v_1035;
assign x_6499 = v_3917 | ~v_912;
assign x_6500 = v_3917 | ~v_913;
assign x_6501 = v_3917 | ~v_806;
assign x_6502 = v_3917 | ~v_807;
assign x_6503 = v_3917 | ~v_3486;
assign x_6504 = v_3917 | ~v_183;
assign x_6505 = v_3917 | ~v_165;
assign x_6506 = v_3917 | ~v_146;
assign x_6507 = v_3917 | ~v_145;
assign x_6508 = v_3917 | ~v_144;
assign x_6509 = v_3917 | ~v_143;
assign x_6510 = v_3917 | ~v_142;
assign x_6511 = v_3917 | ~v_61;
assign x_6512 = v_3917 | ~v_59;
assign x_6513 = v_3917 | ~v_58;
assign x_6514 = v_3917 | ~v_56;
assign x_6515 = v_3917 | ~v_52;
assign x_6516 = v_3916 | ~v_891;
assign x_6517 = v_3916 | ~v_892;
assign x_6518 = v_3916 | ~v_893;
assign x_6519 = v_3916 | ~v_894;
assign x_6520 = v_3916 | ~v_761;
assign x_6521 = v_3916 | ~v_3884;
assign x_6522 = v_3916 | ~v_762;
assign x_6523 = v_3916 | ~v_3885;
assign x_6524 = v_3916 | ~v_763;
assign x_6525 = v_3916 | ~v_764;
assign x_6526 = v_3916 | ~v_3886;
assign x_6527 = v_3916 | ~v_765;
assign x_6528 = v_3916 | ~v_3887;
assign x_6529 = v_3916 | ~v_766;
assign x_6530 = v_3916 | ~v_3522;
assign x_6531 = v_3916 | ~v_3523;
assign x_6532 = v_3916 | ~v_3524;
assign x_6533 = v_3916 | ~v_3525;
assign x_6534 = v_3916 | ~v_3466;
assign x_6535 = v_3916 | ~v_3467;
assign x_6536 = v_3916 | ~v_3468;
assign x_6537 = v_3916 | ~v_3469;
assign x_6538 = v_3916 | ~v_3470;
assign x_6539 = v_3916 | ~v_1027;
assign x_6540 = v_3916 | ~v_1028;
assign x_6541 = v_3916 | ~v_1029;
assign x_6542 = v_3916 | ~v_1030;
assign x_6543 = v_3916 | ~v_897;
assign x_6544 = v_3916 | ~v_898;
assign x_6545 = v_3916 | ~v_773;
assign x_6546 = v_3916 | ~v_774;
assign x_6547 = v_3916 | ~v_182;
assign x_6548 = v_3916 | ~v_161;
assign x_6549 = v_3916 | ~v_138;
assign x_6550 = v_3916 | ~v_137;
assign x_6551 = v_3916 | ~v_3473;
assign x_6552 = v_3916 | ~v_136;
assign x_6553 = v_3916 | ~v_135;
assign x_6554 = v_3916 | ~v_134;
assign x_6555 = v_3916 | ~v_18;
assign x_6556 = v_3916 | ~v_16;
assign x_6557 = v_3916 | ~v_15;
assign x_6558 = v_3916 | ~v_13;
assign x_6559 = v_3916 | ~v_9;
assign x_6560 = ~v_3914 | ~v_3913 | ~v_3912 | v_3915;
assign x_6561 = v_3914 | ~v_877;
assign x_6562 = v_3914 | ~v_878;
assign x_6563 = v_3914 | ~v_879;
assign x_6564 = v_3914 | ~v_880;
assign x_6565 = v_3914 | ~v_827;
assign x_6566 = v_3914 | ~v_3894;
assign x_6567 = v_3914 | ~v_1015;
assign x_6568 = v_3914 | ~v_3895;
assign x_6569 = v_3914 | ~v_1016;
assign x_6570 = v_3914 | ~v_830;
assign x_6571 = v_3914 | ~v_3896;
assign x_6572 = v_3914 | ~v_1017;
assign x_6573 = v_3914 | ~v_3897;
assign x_6574 = v_3914 | ~v_1018;
assign x_6575 = v_3914 | ~v_3616;
assign x_6576 = v_3914 | ~v_3617;
assign x_6577 = v_3914 | ~v_3618;
assign x_6578 = v_3914 | ~v_3619;
assign x_6579 = v_3914 | ~v_3496;
assign x_6580 = v_3914 | ~v_3564;
assign x_6581 = v_3914 | ~v_3565;
assign x_6582 = v_3914 | ~v_3499;
assign x_6583 = v_3914 | ~v_3566;
assign x_6584 = v_3914 | ~v_3567;
assign x_6585 = v_3914 | ~v_885;
assign x_6586 = v_3914 | ~v_1019;
assign x_6587 = v_3914 | ~v_1020;
assign x_6588 = v_3914 | ~v_886;
assign x_6589 = v_3914 | ~v_1021;
assign x_6590 = v_3914 | ~v_1022;
assign x_6591 = v_3914 | ~v_1023;
assign x_6592 = v_3914 | ~v_1024;
assign x_6593 = v_3914 | ~v_184;
assign x_6594 = v_3914 | ~v_181;
assign x_6595 = v_3914 | ~v_171;
assign x_6596 = v_3914 | ~v_170;
assign x_6597 = v_3914 | ~v_169;
assign x_6598 = v_3914 | ~v_148;
assign x_6599 = v_3914 | ~v_147;
assign x_6600 = v_3914 | ~v_103;
assign x_6601 = v_3914 | ~v_102;
assign x_6602 = v_3914 | ~v_101;
assign x_6603 = v_3914 | ~v_99;
assign x_6604 = v_3914 | ~v_97;
assign x_6605 = v_3913 | ~v_862;
assign x_6606 = v_3913 | ~v_863;
assign x_6607 = v_3913 | ~v_864;
assign x_6608 = v_3913 | ~v_865;
assign x_6609 = v_3913 | ~v_794;
assign x_6610 = v_3913 | ~v_3889;
assign x_6611 = v_3913 | ~v_1000;
assign x_6612 = v_3913 | ~v_3890;
assign x_6613 = v_3913 | ~v_1001;
assign x_6614 = v_3913 | ~v_797;
assign x_6615 = v_3913 | ~v_3891;
assign x_6616 = v_3913 | ~v_1002;
assign x_6617 = v_3913 | ~v_3892;
assign x_6618 = v_3913 | ~v_1003;
assign x_6619 = v_3913 | ~v_3611;
assign x_6620 = v_3913 | ~v_3612;
assign x_6621 = v_3913 | ~v_3613;
assign x_6622 = v_3913 | ~v_3614;
assign x_6623 = v_3913 | ~v_3481;
assign x_6624 = v_3913 | ~v_3559;
assign x_6625 = v_3913 | ~v_3560;
assign x_6626 = v_3913 | ~v_3484;
assign x_6627 = v_3913 | ~v_870;
assign x_6628 = v_3913 | ~v_1004;
assign x_6629 = v_3913 | ~v_1005;
assign x_6630 = v_3913 | ~v_871;
assign x_6631 = v_3913 | ~v_1006;
assign x_6632 = v_3913 | ~v_1007;
assign x_6633 = v_3913 | ~v_1008;
assign x_6634 = v_3913 | ~v_1009;
assign x_6635 = v_3913 | ~v_3561;
assign x_6636 = v_3913 | ~v_3562;
assign x_6637 = v_3913 | ~v_183;
assign x_6638 = v_3913 | ~v_180;
assign x_6639 = v_3913 | ~v_167;
assign x_6640 = v_3913 | ~v_166;
assign x_6641 = v_3913 | ~v_165;
assign x_6642 = v_3913 | ~v_143;
assign x_6643 = v_3913 | ~v_142;
assign x_6644 = v_3913 | ~v_61;
assign x_6645 = v_3913 | ~v_60;
assign x_6646 = v_3913 | ~v_59;
assign x_6647 = v_3913 | ~v_57;
assign x_6648 = v_3913 | ~v_55;
assign x_6649 = v_3912 | ~v_847;
assign x_6650 = v_3912 | ~v_848;
assign x_6651 = v_3912 | ~v_849;
assign x_6652 = v_3912 | ~v_850;
assign x_6653 = v_3912 | ~v_761;
assign x_6654 = v_3912 | ~v_3884;
assign x_6655 = v_3912 | ~v_985;
assign x_6656 = v_3912 | ~v_3885;
assign x_6657 = v_3912 | ~v_986;
assign x_6658 = v_3912 | ~v_764;
assign x_6659 = v_3912 | ~v_3886;
assign x_6660 = v_3912 | ~v_987;
assign x_6661 = v_3912 | ~v_3887;
assign x_6662 = v_3912 | ~v_988;
assign x_6663 = v_3912 | ~v_3606;
assign x_6664 = v_3912 | ~v_3607;
assign x_6665 = v_3912 | ~v_3608;
assign x_6666 = v_3912 | ~v_3609;
assign x_6667 = v_3912 | ~v_3466;
assign x_6668 = v_3912 | ~v_3554;
assign x_6669 = v_3912 | ~v_3555;
assign x_6670 = v_3912 | ~v_3469;
assign x_6671 = v_3912 | ~v_3556;
assign x_6672 = v_3912 | ~v_3557;
assign x_6673 = v_3912 | ~v_855;
assign x_6674 = v_3912 | ~v_989;
assign x_6675 = v_3912 | ~v_990;
assign x_6676 = v_3912 | ~v_856;
assign x_6677 = v_3912 | ~v_991;
assign x_6678 = v_3912 | ~v_992;
assign x_6679 = v_3912 | ~v_182;
assign x_6680 = v_3912 | ~v_179;
assign x_6681 = v_3912 | ~v_163;
assign x_6682 = v_3912 | ~v_162;
assign x_6683 = v_3912 | ~v_161;
assign x_6684 = v_3912 | ~v_135;
assign x_6685 = v_3912 | ~v_134;
assign x_6686 = v_3912 | ~v_993;
assign x_6687 = v_3912 | ~v_994;
assign x_6688 = v_3912 | ~v_18;
assign x_6689 = v_3912 | ~v_17;
assign x_6690 = v_3912 | ~v_16;
assign x_6691 = v_3912 | ~v_14;
assign x_6692 = v_3912 | ~v_12;
assign x_6693 = ~v_3910 | ~v_3909 | ~v_3908 | v_3911;
assign x_6694 = v_3910 | ~v_877;
assign x_6695 = v_3910 | ~v_878;
assign x_6696 = v_3910 | ~v_879;
assign x_6697 = v_3910 | ~v_880;
assign x_6698 = v_3910 | ~v_969;
assign x_6699 = v_3910 | ~v_970;
assign x_6700 = v_3910 | ~v_971;
assign x_6701 = v_3910 | ~v_972;
assign x_6702 = v_3910 | ~v_827;
assign x_6703 = v_3910 | ~v_3894;
assign x_6704 = v_3910 | ~v_3895;
assign x_6705 = v_3910 | ~v_830;
assign x_6706 = v_3910 | ~v_3896;
assign x_6707 = v_3910 | ~v_3897;
assign x_6708 = v_3910 | ~v_3616;
assign x_6709 = v_3910 | ~v_3617;
assign x_6710 = v_3910 | ~v_3618;
assign x_6711 = v_3910 | ~v_3619;
assign x_6712 = v_3910 | ~v_3494;
assign x_6713 = v_3910 | ~v_3495;
assign x_6714 = v_3910 | ~v_3496;
assign x_6715 = v_3910 | ~v_3499;
assign x_6716 = v_3910 | ~v_973;
assign x_6717 = v_3910 | ~v_974;
assign x_6718 = v_3910 | ~v_885;
assign x_6719 = v_3910 | ~v_886;
assign x_6720 = v_3910 | ~v_975;
assign x_6721 = v_3910 | ~v_976;
assign x_6722 = v_3910 | ~v_977;
assign x_6723 = v_3910 | ~v_978;
assign x_6724 = v_3910 | ~v_3502;
assign x_6725 = v_3910 | ~v_3503;
assign x_6726 = v_3910 | ~v_184;
assign x_6727 = v_3910 | ~v_181;
assign x_6728 = v_3910 | ~v_172;
assign x_6729 = v_3910 | ~v_171;
assign x_6730 = v_3910 | ~v_170;
assign x_6731 = v_3910 | ~v_169;
assign x_6732 = v_3910 | ~v_150;
assign x_6733 = v_3910 | ~v_149;
assign x_6734 = v_3910 | ~v_147;
assign x_6735 = v_3910 | ~v_102;
assign x_6736 = v_3910 | ~v_101;
assign x_6737 = v_3910 | ~v_96;
assign x_6738 = v_3909 | ~v_862;
assign x_6739 = v_3909 | ~v_863;
assign x_6740 = v_3909 | ~v_864;
assign x_6741 = v_3909 | ~v_865;
assign x_6742 = v_3909 | ~v_954;
assign x_6743 = v_3909 | ~v_955;
assign x_6744 = v_3909 | ~v_956;
assign x_6745 = v_3909 | ~v_957;
assign x_6746 = v_3909 | ~v_794;
assign x_6747 = v_3909 | ~v_3889;
assign x_6748 = v_3909 | ~v_3890;
assign x_6749 = v_3909 | ~v_797;
assign x_6750 = v_3909 | ~v_3891;
assign x_6751 = v_3909 | ~v_3892;
assign x_6752 = v_3909 | ~v_3611;
assign x_6753 = v_3909 | ~v_3612;
assign x_6754 = v_3909 | ~v_3613;
assign x_6755 = v_3909 | ~v_3614;
assign x_6756 = v_3909 | ~v_3479;
assign x_6757 = v_3909 | ~v_3480;
assign x_6758 = v_3909 | ~v_3481;
assign x_6759 = v_3909 | ~v_3484;
assign x_6760 = v_3909 | ~v_958;
assign x_6761 = v_3909 | ~v_959;
assign x_6762 = v_3909 | ~v_870;
assign x_6763 = v_3909 | ~v_871;
assign x_6764 = v_3909 | ~v_960;
assign x_6765 = v_3909 | ~v_961;
assign x_6766 = v_3909 | ~v_962;
assign x_6767 = v_3909 | ~v_963;
assign x_6768 = v_3909 | ~v_3487;
assign x_6769 = v_3909 | ~v_3488;
assign x_6770 = v_3909 | ~v_183;
assign x_6771 = v_3909 | ~v_180;
assign x_6772 = v_3909 | ~v_168;
assign x_6773 = v_3909 | ~v_167;
assign x_6774 = v_3909 | ~v_166;
assign x_6775 = v_3909 | ~v_165;
assign x_6776 = v_3909 | ~v_145;
assign x_6777 = v_3909 | ~v_144;
assign x_6778 = v_3909 | ~v_142;
assign x_6779 = v_3909 | ~v_60;
assign x_6780 = v_3909 | ~v_59;
assign x_6781 = v_3909 | ~v_54;
assign x_6782 = v_3908 | ~v_847;
assign x_6783 = v_3908 | ~v_848;
assign x_6784 = v_3908 | ~v_849;
assign x_6785 = v_3908 | ~v_850;
assign x_6786 = v_3908 | ~v_939;
assign x_6787 = v_3908 | ~v_940;
assign x_6788 = v_3908 | ~v_941;
assign x_6789 = v_3908 | ~v_942;
assign x_6790 = v_3908 | ~v_761;
assign x_6791 = v_3908 | ~v_3884;
assign x_6792 = v_3908 | ~v_3885;
assign x_6793 = v_3908 | ~v_764;
assign x_6794 = v_3908 | ~v_3886;
assign x_6795 = v_3908 | ~v_3887;
assign x_6796 = v_3908 | ~v_3606;
assign x_6797 = v_3908 | ~v_3607;
assign x_6798 = v_3908 | ~v_3608;
assign x_6799 = v_3908 | ~v_3609;
assign x_6800 = v_3908 | ~v_3464;
assign x_6801 = v_3908 | ~v_3465;
assign x_6802 = v_3908 | ~v_3466;
assign x_6803 = v_3908 | ~v_3469;
assign x_6804 = v_3908 | ~v_943;
assign x_6805 = v_3908 | ~v_944;
assign x_6806 = v_3908 | ~v_855;
assign x_6807 = v_3908 | ~v_856;
assign x_6808 = v_3908 | ~v_945;
assign x_6809 = v_3908 | ~v_946;
assign x_6810 = v_3908 | ~v_947;
assign x_6811 = v_3908 | ~v_948;
assign x_6812 = v_3908 | ~v_3471;
assign x_6813 = v_3908 | ~v_3472;
assign x_6814 = v_3908 | ~v_182;
assign x_6815 = v_3908 | ~v_179;
assign x_6816 = v_3908 | ~v_164;
assign x_6817 = v_3908 | ~v_163;
assign x_6818 = v_3908 | ~v_162;
assign x_6819 = v_3908 | ~v_161;
assign x_6820 = v_3908 | ~v_137;
assign x_6821 = v_3908 | ~v_136;
assign x_6822 = v_3908 | ~v_134;
assign x_6823 = v_3908 | ~v_17;
assign x_6824 = v_3908 | ~v_16;
assign x_6825 = v_3908 | ~v_11;
assign x_6826 = ~v_3906 | ~v_3905 | ~v_3904 | v_3907;
assign x_6827 = v_3906 | ~v_877;
assign x_6828 = v_3906 | ~v_878;
assign x_6829 = v_3906 | ~v_879;
assign x_6830 = v_3906 | ~v_880;
assign x_6831 = v_3906 | ~v_921;
assign x_6832 = v_3906 | ~v_922;
assign x_6833 = v_3906 | ~v_923;
assign x_6834 = v_3906 | ~v_924;
assign x_6835 = v_3906 | ~v_827;
assign x_6836 = v_3906 | ~v_3894;
assign x_6837 = v_3906 | ~v_3895;
assign x_6838 = v_3906 | ~v_830;
assign x_6839 = v_3906 | ~v_3896;
assign x_6840 = v_3906 | ~v_3897;
assign x_6841 = v_3906 | ~v_3616;
assign x_6842 = v_3906 | ~v_3617;
assign x_6843 = v_3906 | ~v_3618;
assign x_6844 = v_3906 | ~v_3619;
assign x_6845 = v_3906 | ~v_3532;
assign x_6846 = v_3906 | ~v_3533;
assign x_6847 = v_3906 | ~v_3534;
assign x_6848 = v_3906 | ~v_3535;
assign x_6849 = v_3906 | ~v_3496;
assign x_6850 = v_3906 | ~v_3499;
assign x_6851 = v_3906 | ~v_925;
assign x_6852 = v_3906 | ~v_926;
assign x_6853 = v_3906 | ~v_885;
assign x_6854 = v_3906 | ~v_886;
assign x_6855 = v_3906 | ~v_927;
assign x_6856 = v_3906 | ~v_928;
assign x_6857 = v_3906 | ~v_929;
assign x_6858 = v_3906 | ~v_930;
assign x_6859 = v_3906 | ~v_184;
assign x_6860 = v_3906 | ~v_181;
assign x_6861 = v_3906 | ~v_171;
assign x_6862 = v_3906 | ~v_170;
assign x_6863 = v_3906 | ~v_169;
assign x_6864 = v_3906 | ~v_150;
assign x_6865 = v_3906 | ~v_149;
assign x_6866 = v_3906 | ~v_148;
assign x_6867 = v_3906 | ~v_147;
assign x_6868 = v_3906 | ~v_103;
assign x_6869 = v_3906 | ~v_102;
assign x_6870 = v_3906 | ~v_101;
assign x_6871 = v_3905 | ~v_862;
assign x_6872 = v_3905 | ~v_863;
assign x_6873 = v_3905 | ~v_864;
assign x_6874 = v_3905 | ~v_865;
assign x_6875 = v_3905 | ~v_906;
assign x_6876 = v_3905 | ~v_907;
assign x_6877 = v_3905 | ~v_908;
assign x_6878 = v_3905 | ~v_909;
assign x_6879 = v_3905 | ~v_794;
assign x_6880 = v_3905 | ~v_3889;
assign x_6881 = v_3905 | ~v_3890;
assign x_6882 = v_3905 | ~v_797;
assign x_6883 = v_3905 | ~v_3891;
assign x_6884 = v_3905 | ~v_3892;
assign x_6885 = v_3905 | ~v_3611;
assign x_6886 = v_3905 | ~v_3612;
assign x_6887 = v_3905 | ~v_3613;
assign x_6888 = v_3905 | ~v_3614;
assign x_6889 = v_3905 | ~v_3527;
assign x_6890 = v_3905 | ~v_3528;
assign x_6891 = v_3905 | ~v_3529;
assign x_6892 = v_3905 | ~v_3530;
assign x_6893 = v_3905 | ~v_3481;
assign x_6894 = v_3905 | ~v_3484;
assign x_6895 = v_3905 | ~v_910;
assign x_6896 = v_3905 | ~v_911;
assign x_6897 = v_3905 | ~v_870;
assign x_6898 = v_3905 | ~v_871;
assign x_6899 = v_3905 | ~v_912;
assign x_6900 = v_3905 | ~v_913;
assign x_6901 = v_3905 | ~v_914;
assign x_6902 = v_3905 | ~v_915;
assign x_6903 = v_3905 | ~v_183;
assign x_6904 = v_3905 | ~v_180;
assign x_6905 = v_3905 | ~v_167;
assign x_6906 = v_3905 | ~v_166;
assign x_6907 = v_3905 | ~v_165;
assign x_6908 = v_3905 | ~v_145;
assign x_6909 = v_3905 | ~v_144;
assign x_6910 = v_3905 | ~v_143;
assign x_6911 = v_3905 | ~v_142;
assign x_6912 = v_3905 | ~v_61;
assign x_6913 = v_3905 | ~v_60;
assign x_6914 = v_3905 | ~v_59;
assign x_6915 = v_3904 | ~v_847;
assign x_6916 = v_3904 | ~v_848;
assign x_6917 = v_3904 | ~v_849;
assign x_6918 = v_3904 | ~v_850;
assign x_6919 = v_3904 | ~v_891;
assign x_6920 = v_3904 | ~v_892;
assign x_6921 = v_3904 | ~v_893;
assign x_6922 = v_3904 | ~v_894;
assign x_6923 = v_3904 | ~v_761;
assign x_6924 = v_3904 | ~v_3884;
assign x_6925 = v_3904 | ~v_3885;
assign x_6926 = v_3904 | ~v_764;
assign x_6927 = v_3904 | ~v_3886;
assign x_6928 = v_3904 | ~v_3887;
assign x_6929 = v_3904 | ~v_3606;
assign x_6930 = v_3904 | ~v_3607;
assign x_6931 = v_3904 | ~v_3608;
assign x_6932 = v_3904 | ~v_3609;
assign x_6933 = v_3904 | ~v_3522;
assign x_6934 = v_3904 | ~v_3523;
assign x_6935 = v_3904 | ~v_3524;
assign x_6936 = v_3904 | ~v_3525;
assign x_6937 = v_3904 | ~v_3466;
assign x_6938 = v_3904 | ~v_3469;
assign x_6939 = v_3904 | ~v_895;
assign x_6940 = v_3904 | ~v_896;
assign x_6941 = v_3904 | ~v_855;
assign x_6942 = v_3904 | ~v_856;
assign x_6943 = v_3904 | ~v_897;
assign x_6944 = v_3904 | ~v_898;
assign x_6945 = v_3904 | ~v_899;
assign x_6946 = v_3904 | ~v_900;
assign x_6947 = v_3904 | ~v_182;
assign x_6948 = v_3904 | ~v_179;
assign x_6949 = v_3904 | ~v_163;
assign x_6950 = v_3904 | ~v_162;
assign x_6951 = v_3904 | ~v_161;
assign x_6952 = v_3904 | ~v_137;
assign x_6953 = v_3904 | ~v_136;
assign x_6954 = v_3904 | ~v_135;
assign x_6955 = v_3904 | ~v_134;
assign x_6956 = v_3904 | ~v_18;
assign x_6957 = v_3904 | ~v_17;
assign x_6958 = v_3904 | ~v_16;
assign x_6959 = ~v_3902 | ~v_3901 | ~v_3900 | v_3903;
assign x_6960 = v_3902 | ~v_877;
assign x_6961 = v_3902 | ~v_878;
assign x_6962 = v_3902 | ~v_879;
assign x_6963 = v_3902 | ~v_880;
assign x_6964 = v_3902 | ~v_823;
assign x_6965 = v_3902 | ~v_824;
assign x_6966 = v_3902 | ~v_825;
assign x_6967 = v_3902 | ~v_826;
assign x_6968 = v_3902 | ~v_827;
assign x_6969 = v_3902 | ~v_3894;
assign x_6970 = v_3902 | ~v_3895;
assign x_6971 = v_3902 | ~v_830;
assign x_6972 = v_3902 | ~v_3896;
assign x_6973 = v_3902 | ~v_3897;
assign x_6974 = v_3902 | ~v_3616;
assign x_6975 = v_3902 | ~v_3617;
assign x_6976 = v_3902 | ~v_3618;
assign x_6977 = v_3902 | ~v_3619;
assign x_6978 = v_3902 | ~v_3548;
assign x_6979 = v_3902 | ~v_3549;
assign x_6980 = v_3902 | ~v_3550;
assign x_6981 = v_3902 | ~v_3551;
assign x_6982 = v_3902 | ~v_3496;
assign x_6983 = v_3902 | ~v_3499;
assign x_6984 = v_3902 | ~v_881;
assign x_6985 = v_3902 | ~v_882;
assign x_6986 = v_3902 | ~v_883;
assign x_6987 = v_3902 | ~v_884;
assign x_6988 = v_3902 | ~v_885;
assign x_6989 = v_3902 | ~v_886;
assign x_6990 = v_3902 | ~v_837;
assign x_6991 = v_3902 | ~v_838;
assign x_6992 = v_3902 | ~v_184;
assign x_6993 = v_3902 | ~v_181;
assign x_6994 = v_3902 | ~v_171;
assign x_6995 = v_3902 | ~v_170;
assign x_6996 = v_3902 | ~v_169;
assign x_6997 = v_3902 | ~v_160;
assign x_6998 = v_3902 | ~v_150;
assign x_6999 = v_3902 | ~v_149;
assign x_7000 = v_3902 | ~v_148;
assign x_7001 = v_3902 | ~v_103;
assign x_7002 = v_3902 | ~v_102;
assign x_7003 = v_3902 | ~v_95;
assign x_7004 = v_3901 | ~v_862;
assign x_7005 = v_3901 | ~v_863;
assign x_7006 = v_3901 | ~v_864;
assign x_7007 = v_3901 | ~v_865;
assign x_7008 = v_3901 | ~v_790;
assign x_7009 = v_3901 | ~v_791;
assign x_7010 = v_3901 | ~v_792;
assign x_7011 = v_3901 | ~v_793;
assign x_7012 = v_3901 | ~v_794;
assign x_7013 = v_3901 | ~v_3889;
assign x_7014 = v_3901 | ~v_3890;
assign x_7015 = v_3901 | ~v_797;
assign x_7016 = v_3901 | ~v_3891;
assign x_7017 = v_3901 | ~v_3892;
assign x_7018 = v_3901 | ~v_3611;
assign x_7019 = v_3901 | ~v_3612;
assign x_7020 = v_3901 | ~v_3613;
assign x_7021 = v_3901 | ~v_3614;
assign x_7022 = v_3901 | ~v_3543;
assign x_7023 = v_3901 | ~v_3544;
assign x_7024 = v_3901 | ~v_3545;
assign x_7025 = v_3901 | ~v_3546;
assign x_7026 = v_3901 | ~v_3481;
assign x_7027 = v_3901 | ~v_3484;
assign x_7028 = v_3901 | ~v_866;
assign x_7029 = v_3901 | ~v_867;
assign x_7030 = v_3901 | ~v_868;
assign x_7031 = v_3901 | ~v_869;
assign x_7032 = v_3901 | ~v_870;
assign x_7033 = v_3901 | ~v_871;
assign x_7034 = v_3901 | ~v_804;
assign x_7035 = v_3901 | ~v_805;
assign x_7036 = v_3901 | ~v_183;
assign x_7037 = v_3901 | ~v_180;
assign x_7038 = v_3901 | ~v_167;
assign x_7039 = v_3901 | ~v_166;
assign x_7040 = v_3901 | ~v_165;
assign x_7041 = v_3901 | ~v_159;
assign x_7042 = v_3901 | ~v_145;
assign x_7043 = v_3901 | ~v_144;
assign x_7044 = v_3901 | ~v_143;
assign x_7045 = v_3901 | ~v_61;
assign x_7046 = v_3901 | ~v_60;
assign x_7047 = v_3901 | ~v_53;
assign x_7048 = v_3900 | ~v_847;
assign x_7049 = v_3900 | ~v_848;
assign x_7050 = v_3900 | ~v_849;
assign x_7051 = v_3900 | ~v_850;
assign x_7052 = v_3900 | ~v_757;
assign x_7053 = v_3900 | ~v_758;
assign x_7054 = v_3900 | ~v_759;
assign x_7055 = v_3900 | ~v_760;
assign x_7056 = v_3900 | ~v_761;
assign x_7057 = v_3900 | ~v_3884;
assign x_7058 = v_3900 | ~v_3885;
assign x_7059 = v_3900 | ~v_764;
assign x_7060 = v_3900 | ~v_3886;
assign x_7061 = v_3900 | ~v_3887;
assign x_7062 = v_3900 | ~v_3606;
assign x_7063 = v_3900 | ~v_3607;
assign x_7064 = v_3900 | ~v_3608;
assign x_7065 = v_3900 | ~v_3609;
assign x_7066 = v_3900 | ~v_3538;
assign x_7067 = v_3900 | ~v_3539;
assign x_7068 = v_3900 | ~v_3540;
assign x_7069 = v_3900 | ~v_3541;
assign x_7070 = v_3900 | ~v_3466;
assign x_7071 = v_3900 | ~v_3469;
assign x_7072 = v_3900 | ~v_851;
assign x_7073 = v_3900 | ~v_852;
assign x_7074 = v_3900 | ~v_853;
assign x_7075 = v_3900 | ~v_854;
assign x_7076 = v_3900 | ~v_855;
assign x_7077 = v_3900 | ~v_856;
assign x_7078 = v_3900 | ~v_771;
assign x_7079 = v_3900 | ~v_772;
assign x_7080 = v_3900 | ~v_182;
assign x_7081 = v_3900 | ~v_179;
assign x_7082 = v_3900 | ~v_163;
assign x_7083 = v_3900 | ~v_162;
assign x_7084 = v_3900 | ~v_161;
assign x_7085 = v_3900 | ~v_155;
assign x_7086 = v_3900 | ~v_137;
assign x_7087 = v_3900 | ~v_136;
assign x_7088 = v_3900 | ~v_135;
assign x_7089 = v_3900 | ~v_18;
assign x_7090 = v_3900 | ~v_17;
assign x_7091 = v_3900 | ~v_10;
assign x_7092 = ~v_3898 | ~v_3893 | ~v_3888 | v_3899;
assign x_7093 = v_3898 | ~v_823;
assign x_7094 = v_3898 | ~v_824;
assign x_7095 = v_3898 | ~v_825;
assign x_7096 = v_3898 | ~v_826;
assign x_7097 = v_3898 | ~v_827;
assign x_7098 = v_3898 | ~v_3894;
assign x_7099 = v_3898 | ~v_828;
assign x_7100 = v_3898 | ~v_3895;
assign x_7101 = v_3898 | ~v_829;
assign x_7102 = v_3898 | ~v_830;
assign x_7103 = v_3898 | ~v_3896;
assign x_7104 = v_3898 | ~v_831;
assign x_7105 = v_3898 | ~v_3897;
assign x_7106 = v_3898 | ~v_832;
assign x_7107 = v_3898 | ~v_3548;
assign x_7108 = v_3898 | ~v_3549;
assign x_7109 = v_3898 | ~v_3550;
assign x_7110 = v_3898 | ~v_3551;
assign x_7111 = v_3898 | ~v_3496;
assign x_7112 = v_3898 | ~v_3497;
assign x_7113 = v_3898 | ~v_3498;
assign x_7114 = v_3898 | ~v_3499;
assign x_7115 = v_3898 | ~v_3500;
assign x_7116 = v_3898 | ~v_3501;
assign x_7117 = v_3898 | ~v_833;
assign x_7118 = v_3898 | ~v_834;
assign x_7119 = v_3898 | ~v_835;
assign x_7120 = v_3898 | ~v_836;
assign x_7121 = v_3898 | ~v_837;
assign x_7122 = v_3898 | ~v_838;
assign x_7123 = v_3898 | ~v_839;
assign x_7124 = v_3898 | ~v_840;
assign x_7125 = v_3898 | ~v_184;
assign x_7126 = v_3898 | ~v_169;
assign x_7127 = v_3898 | ~v_160;
assign x_7128 = v_3898 | ~v_150;
assign x_7129 = v_3898 | ~v_149;
assign x_7130 = v_3898 | ~v_148;
assign x_7131 = v_3898 | ~v_147;
assign x_7132 = v_3898 | ~v_103;
assign x_7133 = v_3898 | ~v_102;
assign x_7134 = v_3898 | ~v_100;
assign x_7135 = v_3898 | ~v_98;
assign x_7136 = v_3898 | ~v_94;
assign x_7137 = ~v_123 | ~v_152 | v_3897;
assign x_7138 = ~v_120 | ~v_153 | v_3896;
assign x_7139 = ~v_108 | v_152 | v_3895;
assign x_7140 = ~v_105 | v_153 | v_3894;
assign x_7141 = v_3893 | ~v_790;
assign x_7142 = v_3893 | ~v_791;
assign x_7143 = v_3893 | ~v_792;
assign x_7144 = v_3893 | ~v_793;
assign x_7145 = v_3893 | ~v_794;
assign x_7146 = v_3893 | ~v_3889;
assign x_7147 = v_3893 | ~v_795;
assign x_7148 = v_3893 | ~v_3890;
assign x_7149 = v_3893 | ~v_796;
assign x_7150 = v_3893 | ~v_797;
assign x_7151 = v_3893 | ~v_3891;
assign x_7152 = v_3893 | ~v_798;
assign x_7153 = v_3893 | ~v_3892;
assign x_7154 = v_3893 | ~v_799;
assign x_7155 = v_3893 | ~v_3543;
assign x_7156 = v_3893 | ~v_3544;
assign x_7157 = v_3893 | ~v_3545;
assign x_7158 = v_3893 | ~v_3546;
assign x_7159 = v_3893 | ~v_3481;
assign x_7160 = v_3893 | ~v_3482;
assign x_7161 = v_3893 | ~v_3483;
assign x_7162 = v_3893 | ~v_3484;
assign x_7163 = v_3893 | ~v_3485;
assign x_7164 = v_3893 | ~v_800;
assign x_7165 = v_3893 | ~v_801;
assign x_7166 = v_3893 | ~v_802;
assign x_7167 = v_3893 | ~v_803;
assign x_7168 = v_3893 | ~v_804;
assign x_7169 = v_3893 | ~v_805;
assign x_7170 = v_3893 | ~v_806;
assign x_7171 = v_3893 | ~v_807;
assign x_7172 = v_3893 | ~v_3486;
assign x_7173 = v_3893 | ~v_183;
assign x_7174 = v_3893 | ~v_165;
assign x_7175 = v_3893 | ~v_159;
assign x_7176 = v_3893 | ~v_145;
assign x_7177 = v_3893 | ~v_144;
assign x_7178 = v_3893 | ~v_143;
assign x_7179 = v_3893 | ~v_142;
assign x_7180 = v_3893 | ~v_61;
assign x_7181 = v_3893 | ~v_60;
assign x_7182 = v_3893 | ~v_58;
assign x_7183 = v_3893 | ~v_56;
assign x_7184 = v_3893 | ~v_52;
assign x_7185 = ~v_81 | ~v_152 | v_3892;
assign x_7186 = ~v_78 | ~v_153 | v_3891;
assign x_7187 = ~v_66 | v_152 | v_3890;
assign x_7188 = ~v_63 | v_153 | v_3889;
assign x_7189 = v_3888 | ~v_757;
assign x_7190 = v_3888 | ~v_758;
assign x_7191 = v_3888 | ~v_759;
assign x_7192 = v_3888 | ~v_760;
assign x_7193 = v_3888 | ~v_761;
assign x_7194 = v_3888 | ~v_3884;
assign x_7195 = v_3888 | ~v_762;
assign x_7196 = v_3888 | ~v_3885;
assign x_7197 = v_3888 | ~v_763;
assign x_7198 = v_3888 | ~v_764;
assign x_7199 = v_3888 | ~v_3886;
assign x_7200 = v_3888 | ~v_765;
assign x_7201 = v_3888 | ~v_3887;
assign x_7202 = v_3888 | ~v_766;
assign x_7203 = v_3888 | ~v_3538;
assign x_7204 = v_3888 | ~v_3539;
assign x_7205 = v_3888 | ~v_3540;
assign x_7206 = v_3888 | ~v_3541;
assign x_7207 = v_3888 | ~v_3466;
assign x_7208 = v_3888 | ~v_3467;
assign x_7209 = v_3888 | ~v_3468;
assign x_7210 = v_3888 | ~v_3469;
assign x_7211 = v_3888 | ~v_3470;
assign x_7212 = v_3888 | ~v_767;
assign x_7213 = v_3888 | ~v_768;
assign x_7214 = v_3888 | ~v_769;
assign x_7215 = v_3888 | ~v_770;
assign x_7216 = v_3888 | ~v_771;
assign x_7217 = v_3888 | ~v_772;
assign x_7218 = v_3888 | ~v_773;
assign x_7219 = v_3888 | ~v_774;
assign x_7220 = v_3888 | ~v_182;
assign x_7221 = v_3888 | ~v_161;
assign x_7222 = v_3888 | ~v_155;
assign x_7223 = v_3888 | ~v_137;
assign x_7224 = v_3888 | ~v_3473;
assign x_7225 = v_3888 | ~v_136;
assign x_7226 = v_3888 | ~v_135;
assign x_7227 = v_3888 | ~v_134;
assign x_7228 = v_3888 | ~v_18;
assign x_7229 = v_3888 | ~v_17;
assign x_7230 = v_3888 | ~v_15;
assign x_7231 = v_3888 | ~v_13;
assign x_7232 = v_3888 | ~v_9;
assign x_7233 = ~v_39 | ~v_152 | v_3887;
assign x_7234 = ~v_36 | ~v_153 | v_3886;
assign x_7235 = ~v_24 | v_152 | v_3885;
assign x_7236 = ~v_21 | v_153 | v_3884;
assign x_7237 = v_3883 | ~v_2406;
assign x_7238 = v_3883 | ~v_731;
assign x_7239 = v_3882 | ~v_739;
assign x_7240 = v_3882 | ~v_730;
assign x_7241 = ~v_725 | ~v_724 | ~v_723 | ~v_722 | ~v_3880 | ~v_3876 | ~v_3872 | ~v_3868 | ~v_3864 | ~v_3860 | ~v_3856 | ~v_3852 | ~v_3848 | ~v_3844 | ~v_3840 | ~v_3836 | ~v_3832 | ~v_3828 | ~v_3824 | ~v_3820 | ~v_3804 | v_3881;
assign x_7242 = v_3880 | ~v_3877;
assign x_7243 = v_3880 | ~v_3878;
assign x_7244 = v_3880 | ~v_3879;
assign x_7245 = v_98 | v_103 | v_101 | v_97 | v_100 | v_95 | v_94 | v_99 | v_102 | ~v_719 | ~v_718 | v_169 | v_148 | v_184 | ~v_483 | ~v_717 | ~v_299 | ~v_482 | ~v_716 | ~v_298 | ~v_3386 | ~v_3320 | ~v_3385 | ~v_3319 | ~v_3318 | ~v_3384 | ~v_3317 | ~v_3383 | ~v_3316 | ~v_3315 | ~v_477 | ~v_291 | ~v_3818 | ~v_476 | ~v_290 | ~v_3817 | ~v_289 | ~v_475 | ~v_288 | ~v_3816 | ~v_474 | ~v_287 | ~v_3815 | ~v_286 | v_3879;
assign x_7246 = v_53 | v_56 | v_55 | v_61 | v_52 | v_60 | v_59 | v_58 | v_57 | ~v_714 | ~v_713 | v_143 | v_165 | v_183 | ~v_3381 | ~v_3305 | ~v_266 | ~v_3380 | ~v_468 | ~v_712 | ~v_467 | ~v_711 | ~v_265 | ~v_3304 | ~v_3303 | ~v_3379 | ~v_3302 | ~v_3378 | ~v_3301 | ~v_3300 | ~v_462 | ~v_258 | ~v_3813 | ~v_461 | ~v_257 | ~v_3812 | ~v_256 | ~v_460 | ~v_255 | ~v_3811 | ~v_459 | ~v_254 | ~v_3810 | ~v_253 | v_3878;
assign x_7247 = v_13 | v_9 | v_18 | v_17 | v_16 | v_15 | v_14 | v_12 | v_10 | ~v_453 | ~v_709 | ~v_452 | ~v_708 | v_135 | ~v_707 | ~v_706 | ~v_3292 | v_161 | v_182 | ~v_233 | ~v_232 | ~v_3376 | ~v_3289 | ~v_3375 | ~v_3288 | ~v_3374 | ~v_3287 | ~v_3373 | ~v_3286 | ~v_3285 | ~v_447 | ~v_225 | ~v_3808 | ~v_446 | ~v_224 | ~v_3807 | ~v_223 | ~v_445 | ~v_222 | ~v_3806 | ~v_444 | ~v_221 | ~v_3805 | ~v_220 | v_3877;
assign x_7248 = v_3876 | ~v_3873;
assign x_7249 = v_3876 | ~v_3874;
assign x_7250 = v_3876 | ~v_3875;
assign x_7251 = v_103 | v_101 | v_97 | v_100 | v_99 | v_93 | v_102 | v_171 | v_170 | v_148 | v_147 | v_184 | ~v_703 | ~v_702 | ~v_483 | ~v_482 | ~v_701 | ~v_653 | ~v_700 | ~v_652 | ~v_3386 | ~v_3385 | ~v_3318 | ~v_3384 | ~v_3383 | ~v_3315 | ~v_3338 | ~v_3337 | ~v_3336 | ~v_3335 | ~v_477 | ~v_3818 | ~v_476 | ~v_3817 | ~v_289 | ~v_475 | ~v_3816 | ~v_474 | ~v_3815 | ~v_286 | ~v_649 | ~v_648 | ~v_647 | ~v_646 | v_3875;
assign x_7252 = v_55 | v_61 | v_51 | v_60 | v_59 | v_58 | v_57 | v_143 | v_142 | v_167 | v_166 | v_183 | ~v_698 | ~v_697 | ~v_3381 | ~v_3380 | ~v_468 | ~v_467 | ~v_696 | ~v_638 | ~v_695 | ~v_637 | ~v_3303 | ~v_3379 | ~v_3378 | ~v_3300 | ~v_3333 | ~v_3332 | ~v_3331 | ~v_3330 | ~v_462 | ~v_3813 | ~v_461 | ~v_3812 | ~v_256 | ~v_460 | ~v_3811 | ~v_459 | ~v_3810 | ~v_253 | ~v_634 | ~v_633 | ~v_632 | ~v_631 | v_3874;
assign x_7253 = v_18 | v_17 | v_16 | v_8 | v_15 | v_14 | v_12 | ~v_453 | ~v_452 | v_135 | v_134 | v_163 | v_162 | v_182 | ~v_693 | ~v_692 | ~v_691 | ~v_623 | ~v_690 | ~v_622 | ~v_3376 | ~v_3375 | ~v_3288 | ~v_3374 | ~v_3373 | ~v_3285 | ~v_3328 | ~v_3327 | ~v_3326 | ~v_3325 | ~v_447 | ~v_3808 | ~v_446 | ~v_3807 | ~v_223 | ~v_445 | ~v_3806 | ~v_444 | ~v_3805 | ~v_220 | ~v_619 | ~v_618 | ~v_617 | ~v_616 | v_3873;
assign x_7254 = v_3872 | ~v_3869;
assign x_7255 = v_3872 | ~v_3870;
assign x_7256 = v_3872 | ~v_3871;
assign x_7257 = v_103 | v_101 | v_96 | v_100 | v_95 | v_93 | v_102 | v_171 | v_170 | v_150 | v_149 | v_184 | ~v_3322 | ~v_3321 | ~v_435 | ~v_434 | ~v_653 | ~v_652 | ~v_687 | ~v_686 | ~v_685 | ~v_684 | ~v_3318 | ~v_3315 | ~v_3314 | ~v_3313 | ~v_3338 | ~v_3337 | ~v_3336 | ~v_3335 | ~v_3818 | ~v_3817 | ~v_289 | ~v_3816 | ~v_3815 | ~v_286 | ~v_649 | ~v_648 | ~v_647 | ~v_646 | ~v_431 | ~v_430 | ~v_429 | ~v_428 | v_3871;
assign x_7258 = v_54 | v_53 | v_61 | v_51 | v_60 | v_59 | v_58 | v_144 | v_145 | v_167 | v_166 | v_183 | ~v_3307 | ~v_3306 | ~v_420 | ~v_419 | ~v_638 | ~v_637 | ~v_682 | ~v_681 | ~v_680 | ~v_679 | ~v_3303 | ~v_3300 | ~v_3299 | ~v_3298 | ~v_3333 | ~v_3332 | ~v_3331 | ~v_3330 | ~v_3813 | ~v_3812 | ~v_256 | ~v_3811 | ~v_3810 | ~v_253 | ~v_634 | ~v_633 | ~v_632 | ~v_631 | ~v_416 | ~v_415 | ~v_414 | ~v_413 | v_3870;
assign x_7259 = v_18 | v_17 | v_16 | v_8 | v_15 | v_11 | v_10 | v_136 | v_137 | v_163 | v_162 | v_182 | ~v_3291 | ~v_3290 | ~v_405 | ~v_404 | ~v_623 | ~v_622 | ~v_677 | ~v_676 | ~v_675 | ~v_674 | ~v_3288 | ~v_3285 | ~v_3284 | ~v_3283 | ~v_3328 | ~v_3327 | ~v_3326 | ~v_3325 | ~v_3808 | ~v_3807 | ~v_223 | ~v_3806 | ~v_3805 | ~v_220 | ~v_619 | ~v_618 | ~v_617 | ~v_616 | ~v_401 | ~v_400 | ~v_399 | ~v_398 | v_3869;
assign x_7260 = v_3868 | ~v_3865;
assign x_7261 = v_3868 | ~v_3866;
assign x_7262 = v_3868 | ~v_3867;
assign x_7263 = v_101 | v_100 | v_93 | v_102 | v_172 | v_171 | v_170 | v_150 | v_149 | v_148 | v_147 | v_184 | ~v_671 | ~v_670 | ~v_387 | ~v_386 | ~v_653 | ~v_652 | ~v_669 | ~v_668 | ~v_3318 | ~v_3315 | ~v_3354 | ~v_3353 | ~v_3352 | ~v_3351 | ~v_3338 | ~v_3337 | ~v_3336 | ~v_3335 | ~v_3818 | ~v_3817 | ~v_289 | ~v_3816 | ~v_3815 | ~v_286 | ~v_649 | ~v_648 | ~v_647 | ~v_646 | ~v_383 | ~v_382 | ~v_381 | ~v_380 | v_3867;
assign x_7264 = v_51 | v_60 | v_59 | v_58 | v_144 | v_145 | v_143 | v_142 | v_168 | v_167 | v_166 | v_183 | ~v_666 | ~v_665 | ~v_372 | ~v_371 | ~v_638 | ~v_637 | ~v_664 | ~v_663 | ~v_3303 | ~v_3300 | ~v_3349 | ~v_3348 | ~v_3347 | ~v_3346 | ~v_3333 | ~v_3332 | ~v_3331 | ~v_3330 | ~v_3813 | ~v_3812 | ~v_256 | ~v_3811 | ~v_3810 | ~v_253 | ~v_634 | ~v_633 | ~v_632 | ~v_631 | ~v_368 | ~v_367 | ~v_366 | ~v_365 | v_3866;
assign x_7265 = v_17 | v_16 | v_8 | v_15 | v_136 | v_135 | v_134 | v_137 | v_164 | v_163 | v_162 | v_182 | ~v_661 | ~v_660 | ~v_357 | ~v_356 | ~v_623 | ~v_622 | ~v_659 | ~v_658 | ~v_3288 | ~v_3285 | ~v_3344 | ~v_3343 | ~v_3342 | ~v_3341 | ~v_3328 | ~v_3327 | ~v_3326 | ~v_3325 | ~v_3808 | ~v_3807 | ~v_223 | ~v_3806 | ~v_3805 | ~v_220 | ~v_619 | ~v_618 | ~v_617 | ~v_616 | ~v_353 | ~v_352 | ~v_351 | ~v_350 | v_3865;
assign x_7266 = v_3864 | ~v_3861;
assign x_7267 = v_3864 | ~v_3862;
assign x_7268 = v_3864 | ~v_3863;
assign x_7269 = v_103 | v_100 | v_93 | v_151 | v_171 | v_170 | v_160 | v_150 | v_149 | v_148 | v_147 | v_184 | ~v_655 | ~v_654 | ~v_297 | ~v_296 | ~v_653 | ~v_652 | ~v_651 | ~v_650 | ~v_3318 | ~v_3315 | ~v_3370 | ~v_3369 | ~v_3368 | ~v_3367 | ~v_3338 | ~v_3337 | ~v_3336 | ~v_3335 | ~v_3818 | ~v_3817 | ~v_289 | ~v_3816 | ~v_3815 | ~v_286 | ~v_649 | ~v_648 | ~v_647 | ~v_646 | ~v_285 | ~v_284 | ~v_283 | ~v_282 | v_3863;
assign x_7270 = v_61 | v_51 | v_58 | v_144 | v_159 | v_145 | v_143 | v_142 | v_167 | v_166 | v_146 | v_183 | ~v_640 | ~v_639 | ~v_264 | ~v_263 | ~v_638 | ~v_637 | ~v_636 | ~v_635 | ~v_3303 | ~v_3300 | ~v_3365 | ~v_3364 | ~v_3363 | ~v_3362 | ~v_3333 | ~v_3332 | ~v_3331 | ~v_3330 | ~v_3813 | ~v_3812 | ~v_256 | ~v_3811 | ~v_3810 | ~v_253 | ~v_634 | ~v_633 | ~v_632 | ~v_631 | ~v_252 | ~v_251 | ~v_250 | ~v_249 | v_3862;
assign x_7271 = v_18 | v_8 | v_15 | v_136 | v_135 | v_134 | v_137 | v_138 | v_163 | v_162 | v_155 | v_182 | ~v_625 | ~v_624 | ~v_231 | ~v_230 | ~v_623 | ~v_622 | ~v_621 | ~v_620 | ~v_3288 | ~v_3285 | ~v_3360 | ~v_3359 | ~v_3358 | ~v_3357 | ~v_3328 | ~v_3327 | ~v_3326 | ~v_3325 | ~v_3808 | ~v_3807 | ~v_223 | ~v_3806 | ~v_3805 | ~v_220 | ~v_619 | ~v_618 | ~v_617 | ~v_616 | ~v_219 | ~v_218 | ~v_217 | ~v_216 | v_3861;
assign x_7272 = v_3860 | ~v_3857;
assign x_7273 = v_3860 | ~v_3858;
assign x_7274 = v_3860 | ~v_3859;
assign x_7275 = v_98 | v_103 | v_101 | v_96 | v_100 | v_94 | v_102 | v_169 | v_150 | v_149 | v_147 | v_184 | ~v_609 | ~v_608 | ~v_3322 | ~v_3321 | ~v_299 | ~v_298 | ~v_435 | ~v_434 | ~v_607 | ~v_606 | ~v_3320 | ~v_3319 | ~v_3318 | ~v_3317 | ~v_3316 | ~v_3315 | ~v_3314 | ~v_3313 | ~v_291 | ~v_3818 | ~v_290 | ~v_3817 | ~v_289 | ~v_288 | ~v_3816 | ~v_287 | ~v_3815 | ~v_286 | ~v_431 | ~v_430 | ~v_429 | ~v_428 | v_3859;
assign x_7276 = v_54 | v_56 | v_61 | v_52 | v_60 | v_59 | v_58 | v_144 | v_145 | v_142 | v_165 | v_183 | ~v_604 | ~v_603 | ~v_3307 | ~v_3306 | ~v_3305 | ~v_266 | ~v_265 | ~v_420 | ~v_419 | ~v_602 | ~v_601 | ~v_3304 | ~v_3303 | ~v_3302 | ~v_3301 | ~v_3300 | ~v_3299 | ~v_3298 | ~v_258 | ~v_3813 | ~v_257 | ~v_3812 | ~v_256 | ~v_255 | ~v_3811 | ~v_254 | ~v_3810 | ~v_253 | ~v_416 | ~v_415 | ~v_414 | ~v_413 | v_3858;
assign x_7277 = v_13 | v_9 | v_18 | v_17 | v_16 | v_15 | v_11 | v_136 | v_134 | ~v_3292 | v_137 | v_161 | v_182 | ~v_599 | ~v_598 | ~v_3291 | ~v_3290 | ~v_233 | ~v_232 | ~v_405 | ~v_404 | ~v_597 | ~v_596 | ~v_3289 | ~v_3288 | ~v_3287 | ~v_3286 | ~v_3285 | ~v_3284 | ~v_3283 | ~v_225 | ~v_3808 | ~v_224 | ~v_3807 | ~v_223 | ~v_222 | ~v_3806 | ~v_221 | ~v_3805 | ~v_220 | ~v_401 | ~v_400 | ~v_399 | ~v_398 | v_3857;
assign x_7278 = v_3856 | ~v_3853;
assign x_7279 = v_3856 | ~v_3854;
assign x_7280 = v_3856 | ~v_3855;
assign x_7281 = v_101 | v_97 | v_100 | v_99 | v_102 | v_172 | v_171 | v_170 | v_169 | v_148 | v_147 | v_184 | ~v_483 | ~v_482 | ~v_593 | ~v_592 | ~v_545 | ~v_591 | ~v_590 | ~v_544 | ~v_3386 | ~v_3385 | ~v_3318 | ~v_3384 | ~v_3383 | ~v_3315 | ~v_3406 | ~v_3405 | ~v_3404 | ~v_3403 | ~v_477 | ~v_3818 | ~v_476 | ~v_3817 | ~v_289 | ~v_475 | ~v_3816 | ~v_474 | ~v_3815 | ~v_286 | ~v_539 | ~v_538 | ~v_537 | ~v_536 | v_3855;
assign x_7282 = v_55 | v_60 | v_59 | v_58 | v_57 | v_143 | v_142 | v_168 | v_167 | v_166 | v_165 | v_183 | ~v_3381 | ~v_3380 | ~v_468 | ~v_467 | ~v_588 | ~v_587 | ~v_530 | ~v_586 | ~v_585 | ~v_529 | ~v_3303 | ~v_3379 | ~v_3378 | ~v_3300 | ~v_3401 | ~v_3400 | ~v_3399 | ~v_3398 | ~v_462 | ~v_3813 | ~v_461 | ~v_3812 | ~v_256 | ~v_460 | ~v_3811 | ~v_459 | ~v_3810 | ~v_253 | ~v_524 | ~v_523 | ~v_522 | ~v_521 | v_3854;
assign x_7283 = v_17 | v_16 | v_15 | v_14 | v_12 | ~v_453 | ~v_452 | v_135 | v_134 | v_164 | v_163 | v_162 | v_161 | v_182 | ~v_583 | ~v_582 | ~v_515 | ~v_581 | ~v_580 | ~v_514 | ~v_3376 | ~v_3375 | ~v_3288 | ~v_3374 | ~v_3373 | ~v_3285 | ~v_3396 | ~v_3395 | ~v_3394 | ~v_3393 | ~v_447 | ~v_3808 | ~v_446 | ~v_3807 | ~v_223 | ~v_445 | ~v_3806 | ~v_444 | ~v_3805 | ~v_220 | ~v_509 | ~v_508 | ~v_507 | ~v_506 | v_3853;
assign x_7284 = v_3852 | ~v_3849;
assign x_7285 = v_3852 | ~v_3850;
assign x_7286 = v_3852 | ~v_3851;
assign x_7287 = v_103 | v_101 | v_96 | v_100 | v_151 | v_171 | v_170 | v_169 | v_150 | v_149 | v_147 | v_184 | ~v_3322 | ~v_3321 | ~v_577 | ~v_576 | ~v_545 | ~v_544 | ~v_575 | ~v_574 | ~v_435 | ~v_434 | ~v_3318 | ~v_3315 | ~v_3406 | ~v_3405 | ~v_3404 | ~v_3403 | ~v_3314 | ~v_3313 | ~v_3818 | ~v_3817 | ~v_289 | ~v_3816 | ~v_3815 | ~v_286 | ~v_431 | ~v_430 | ~v_429 | ~v_428 | ~v_539 | ~v_538 | ~v_537 | ~v_536 | v_3851;
assign x_7288 = v_54 | v_61 | v_59 | v_58 | v_144 | v_145 | v_142 | v_167 | v_166 | v_165 | v_146 | v_183 | ~v_3307 | ~v_3306 | ~v_572 | ~v_571 | ~v_530 | ~v_529 | ~v_570 | ~v_569 | ~v_420 | ~v_419 | ~v_3303 | ~v_3300 | ~v_3401 | ~v_3400 | ~v_3399 | ~v_3398 | ~v_3299 | ~v_3298 | ~v_3813 | ~v_3812 | ~v_256 | ~v_3811 | ~v_3810 | ~v_253 | ~v_416 | ~v_415 | ~v_414 | ~v_413 | ~v_524 | ~v_523 | ~v_522 | ~v_521 | v_3850;
assign x_7289 = v_18 | v_16 | v_15 | v_11 | v_136 | v_134 | v_137 | v_138 | v_163 | v_162 | v_161 | v_182 | ~v_3291 | ~v_3290 | ~v_567 | ~v_566 | ~v_515 | ~v_514 | ~v_565 | ~v_564 | ~v_405 | ~v_404 | ~v_3288 | ~v_3285 | ~v_3396 | ~v_3395 | ~v_3394 | ~v_3393 | ~v_3284 | ~v_3283 | ~v_3808 | ~v_3807 | ~v_223 | ~v_3806 | ~v_3805 | ~v_220 | ~v_401 | ~v_400 | ~v_399 | ~v_398 | ~v_509 | ~v_508 | ~v_507 | ~v_506 | v_3849;
assign x_7290 = v_3848 | ~v_3845;
assign x_7291 = v_3848 | ~v_3846;
assign x_7292 = v_3848 | ~v_3847;
assign x_7293 = v_103 | v_101 | v_100 | v_95 | v_102 | v_171 | v_170 | v_169 | v_150 | v_149 | v_148 | v_184 | ~v_545 | ~v_544 | ~v_561 | ~v_560 | ~v_559 | ~v_558 | ~v_387 | ~v_386 | ~v_3318 | ~v_3315 | ~v_3406 | ~v_3405 | ~v_3404 | ~v_3403 | ~v_3354 | ~v_3353 | ~v_3352 | ~v_3351 | ~v_3818 | ~v_3817 | ~v_289 | ~v_3816 | ~v_3815 | ~v_286 | ~v_383 | ~v_382 | ~v_381 | ~v_380 | ~v_539 | ~v_538 | ~v_537 | ~v_536 | v_3847;
assign x_7294 = v_53 | v_61 | v_60 | v_59 | v_58 | v_144 | v_145 | v_143 | v_167 | v_166 | v_165 | v_183 | ~v_530 | ~v_529 | ~v_556 | ~v_555 | ~v_554 | ~v_553 | ~v_372 | ~v_371 | ~v_3303 | ~v_3300 | ~v_3401 | ~v_3400 | ~v_3399 | ~v_3398 | ~v_3349 | ~v_3348 | ~v_3347 | ~v_3346 | ~v_3813 | ~v_3812 | ~v_256 | ~v_3811 | ~v_3810 | ~v_253 | ~v_368 | ~v_367 | ~v_366 | ~v_365 | ~v_524 | ~v_523 | ~v_522 | ~v_521 | v_3846;
assign x_7295 = v_18 | v_17 | v_16 | v_15 | v_10 | v_136 | v_135 | v_137 | v_163 | v_162 | v_161 | v_182 | ~v_515 | ~v_514 | ~v_551 | ~v_550 | ~v_549 | ~v_548 | ~v_357 | ~v_356 | ~v_3288 | ~v_3285 | ~v_3396 | ~v_3395 | ~v_3394 | ~v_3393 | ~v_3344 | ~v_3343 | ~v_3342 | ~v_3341 | ~v_3808 | ~v_3807 | ~v_223 | ~v_3806 | ~v_3805 | ~v_220 | ~v_353 | ~v_352 | ~v_351 | ~v_350 | ~v_509 | ~v_508 | ~v_507 | ~v_506 | v_3845;
assign x_7296 = v_3844 | ~v_3841;
assign x_7297 = v_3844 | ~v_3842;
assign x_7298 = v_3844 | ~v_3843;
assign x_7299 = v_103 | v_100 | v_102 | v_171 | v_170 | v_169 | v_160 | v_150 | v_149 | v_148 | v_147 | v_184 | ~v_545 | ~v_544 | ~v_543 | ~v_542 | ~v_541 | ~v_540 | ~v_297 | ~v_296 | ~v_3318 | ~v_3315 | ~v_3406 | ~v_3405 | ~v_3404 | ~v_3403 | ~v_3370 | ~v_3369 | ~v_3368 | ~v_3367 | ~v_3818 | ~v_3817 | ~v_289 | ~v_3816 | ~v_3815 | ~v_286 | ~v_285 | ~v_284 | ~v_283 | ~v_282 | ~v_539 | ~v_538 | ~v_537 | ~v_536 | v_3843;
assign x_7300 = v_61 | v_60 | v_58 | v_144 | v_159 | v_145 | v_143 | v_142 | v_167 | v_166 | v_165 | v_183 | ~v_530 | ~v_529 | ~v_528 | ~v_527 | ~v_526 | ~v_525 | ~v_264 | ~v_263 | ~v_3303 | ~v_3300 | ~v_3401 | ~v_3400 | ~v_3399 | ~v_3398 | ~v_3365 | ~v_3364 | ~v_3363 | ~v_3362 | ~v_3813 | ~v_3812 | ~v_256 | ~v_3811 | ~v_3810 | ~v_253 | ~v_252 | ~v_251 | ~v_250 | ~v_249 | ~v_524 | ~v_523 | ~v_522 | ~v_521 | v_3842;
assign x_7301 = v_18 | v_17 | v_15 | v_136 | v_135 | v_134 | v_137 | v_163 | v_162 | v_161 | v_155 | v_182 | ~v_515 | ~v_514 | ~v_513 | ~v_512 | ~v_511 | ~v_510 | ~v_231 | ~v_230 | ~v_3288 | ~v_3285 | ~v_3396 | ~v_3395 | ~v_3394 | ~v_3393 | ~v_3360 | ~v_3359 | ~v_3358 | ~v_3357 | ~v_3808 | ~v_3807 | ~v_223 | ~v_3806 | ~v_3805 | ~v_220 | ~v_219 | ~v_218 | ~v_217 | ~v_216 | ~v_509 | ~v_508 | ~v_507 | ~v_506 | v_3841;
assign x_7302 = v_3840 | ~v_3837;
assign x_7303 = v_3840 | ~v_3838;
assign x_7304 = v_3840 | ~v_3839;
assign x_7305 = v_98 | v_103 | v_101 | v_100 | v_94 | v_151 | v_169 | v_150 | v_149 | v_148 | v_147 | v_184 | ~v_299 | ~v_298 | ~v_387 | ~v_386 | ~v_499 | ~v_498 | ~v_497 | ~v_496 | ~v_3320 | ~v_3319 | ~v_3318 | ~v_3317 | ~v_3316 | ~v_3315 | ~v_3354 | ~v_3353 | ~v_3352 | ~v_3351 | ~v_291 | ~v_3818 | ~v_290 | ~v_3817 | ~v_289 | ~v_288 | ~v_3816 | ~v_287 | ~v_3815 | ~v_286 | ~v_383 | ~v_382 | ~v_381 | ~v_380 | v_3839;
assign x_7306 = v_56 | v_61 | v_52 | v_59 | v_58 | v_144 | v_145 | v_143 | v_142 | v_165 | v_146 | v_183 | ~v_3305 | ~v_266 | ~v_265 | ~v_372 | ~v_371 | ~v_494 | ~v_493 | ~v_492 | ~v_491 | ~v_3304 | ~v_3303 | ~v_3302 | ~v_3301 | ~v_3300 | ~v_3349 | ~v_3348 | ~v_3347 | ~v_3346 | ~v_258 | ~v_3813 | ~v_257 | ~v_3812 | ~v_256 | ~v_255 | ~v_3811 | ~v_254 | ~v_3810 | ~v_253 | ~v_368 | ~v_367 | ~v_366 | ~v_365 | v_3838;
assign x_7307 = v_13 | v_9 | v_18 | v_16 | v_15 | v_136 | v_135 | v_134 | ~v_3292 | v_137 | v_138 | v_161 | v_182 | ~v_233 | ~v_232 | ~v_357 | ~v_356 | ~v_489 | ~v_488 | ~v_487 | ~v_486 | ~v_3289 | ~v_3288 | ~v_3287 | ~v_3286 | ~v_3285 | ~v_3344 | ~v_3343 | ~v_3342 | ~v_3341 | ~v_225 | ~v_3808 | ~v_224 | ~v_3807 | ~v_223 | ~v_222 | ~v_3806 | ~v_221 | ~v_3805 | ~v_220 | ~v_353 | ~v_352 | ~v_351 | ~v_350 | v_3837;
assign x_7308 = v_3836 | ~v_3833;
assign x_7309 = v_3836 | ~v_3834;
assign x_7310 = v_3836 | ~v_3835;
assign x_7311 = v_103 | v_101 | v_97 | v_99 | v_102 | v_171 | v_170 | v_169 | v_148 | v_147 | v_184 | v_181 | ~v_483 | ~v_482 | ~v_481 | ~v_480 | ~v_345 | ~v_479 | ~v_478 | ~v_344 | ~v_3386 | ~v_3385 | ~v_3318 | ~v_3384 | ~v_3383 | ~v_3315 | ~v_3438 | ~v_3437 | ~v_3436 | ~v_3435 | ~v_477 | ~v_3818 | ~v_476 | ~v_3817 | ~v_289 | ~v_475 | ~v_3816 | ~v_474 | ~v_3815 | ~v_286 | ~v_339 | ~v_338 | ~v_337 | ~v_336 | v_3835;
assign x_7312 = v_55 | v_61 | v_60 | v_59 | v_57 | v_180 | v_143 | v_142 | v_167 | v_166 | v_165 | v_183 | ~v_3381 | ~v_3380 | ~v_468 | ~v_467 | ~v_466 | ~v_465 | ~v_330 | ~v_464 | ~v_463 | ~v_329 | ~v_3303 | ~v_3379 | ~v_3378 | ~v_3300 | ~v_3433 | ~v_3432 | ~v_3431 | ~v_3430 | ~v_462 | ~v_3813 | ~v_461 | ~v_3812 | ~v_256 | ~v_460 | ~v_3811 | ~v_459 | ~v_3810 | ~v_253 | ~v_324 | ~v_323 | ~v_322 | ~v_321 | v_3834;
assign x_7313 = v_18 | v_17 | v_16 | v_14 | v_12 | ~v_453 | ~v_452 | v_135 | v_134 | v_179 | v_163 | v_162 | v_161 | v_182 | ~v_451 | ~v_450 | ~v_315 | ~v_449 | ~v_448 | ~v_314 | ~v_3376 | ~v_3375 | ~v_3288 | ~v_3374 | ~v_3373 | ~v_3285 | ~v_3428 | ~v_3427 | ~v_3426 | ~v_3425 | ~v_447 | ~v_3808 | ~v_446 | ~v_3807 | ~v_223 | ~v_445 | ~v_3806 | ~v_444 | ~v_3805 | ~v_220 | ~v_309 | ~v_308 | ~v_307 | ~v_306 | v_3833;
assign x_7314 = v_3832 | ~v_3829;
assign x_7315 = v_3832 | ~v_3830;
assign x_7316 = v_3832 | ~v_3831;
assign x_7317 = v_101 | v_96 | v_102 | v_172 | v_171 | v_170 | v_169 | v_150 | v_149 | v_147 | v_184 | v_181 | ~v_3322 | ~v_3321 | ~v_437 | ~v_436 | ~v_435 | ~v_434 | ~v_345 | ~v_344 | ~v_433 | ~v_432 | ~v_3318 | ~v_3315 | ~v_3314 | ~v_3313 | ~v_3438 | ~v_3437 | ~v_3436 | ~v_3435 | ~v_3818 | ~v_3817 | ~v_289 | ~v_3816 | ~v_3815 | ~v_286 | ~v_431 | ~v_430 | ~v_429 | ~v_428 | ~v_339 | ~v_338 | ~v_337 | ~v_336 | v_3831;
assign x_7318 = v_54 | v_60 | v_59 | v_144 | v_180 | v_145 | v_142 | v_168 | v_167 | v_166 | v_165 | v_183 | ~v_3307 | ~v_3306 | ~v_422 | ~v_421 | ~v_420 | ~v_419 | ~v_330 | ~v_329 | ~v_418 | ~v_417 | ~v_3303 | ~v_3300 | ~v_3299 | ~v_3298 | ~v_3433 | ~v_3432 | ~v_3431 | ~v_3430 | ~v_3813 | ~v_3812 | ~v_256 | ~v_3811 | ~v_3810 | ~v_253 | ~v_416 | ~v_415 | ~v_414 | ~v_413 | ~v_324 | ~v_323 | ~v_322 | ~v_321 | v_3830;
assign x_7319 = v_17 | v_16 | v_11 | v_136 | v_134 | v_137 | v_179 | v_164 | v_163 | v_162 | v_161 | v_182 | ~v_3291 | ~v_3290 | ~v_407 | ~v_406 | ~v_405 | ~v_404 | ~v_315 | ~v_314 | ~v_403 | ~v_402 | ~v_3288 | ~v_3285 | ~v_3284 | ~v_3283 | ~v_3428 | ~v_3427 | ~v_3426 | ~v_3425 | ~v_3808 | ~v_3807 | ~v_223 | ~v_3806 | ~v_3805 | ~v_220 | ~v_401 | ~v_400 | ~v_399 | ~v_398 | ~v_309 | ~v_308 | ~v_307 | ~v_306 | v_3829;
assign x_7320 = v_3828 | ~v_3825;
assign x_7321 = v_3828 | ~v_3826;
assign x_7322 = v_3828 | ~v_3827;
assign x_7323 = v_103 | v_101 | v_102 | v_171 | v_170 | v_169 | v_150 | v_149 | v_148 | v_147 | v_184 | v_181 | ~v_391 | ~v_390 | ~v_387 | ~v_386 | ~v_345 | ~v_344 | ~v_385 | ~v_384 | ~v_3318 | ~v_3315 | ~v_3354 | ~v_3353 | ~v_3352 | ~v_3351 | ~v_3438 | ~v_3437 | ~v_3436 | ~v_3435 | ~v_3818 | ~v_3817 | ~v_289 | ~v_3816 | ~v_3815 | ~v_286 | ~v_383 | ~v_382 | ~v_381 | ~v_380 | ~v_339 | ~v_338 | ~v_337 | ~v_336 | v_3827;
assign x_7324 = v_61 | v_60 | v_59 | v_144 | v_180 | v_145 | v_143 | v_142 | v_167 | v_166 | v_165 | v_183 | ~v_376 | ~v_375 | ~v_372 | ~v_371 | ~v_330 | ~v_329 | ~v_370 | ~v_369 | ~v_3303 | ~v_3300 | ~v_3349 | ~v_3348 | ~v_3347 | ~v_3346 | ~v_3433 | ~v_3432 | ~v_3431 | ~v_3430 | ~v_3813 | ~v_3812 | ~v_256 | ~v_3811 | ~v_3810 | ~v_253 | ~v_368 | ~v_367 | ~v_366 | ~v_365 | ~v_324 | ~v_323 | ~v_322 | ~v_321 | v_3826;
assign x_7325 = v_18 | v_17 | v_16 | v_136 | v_135 | v_134 | v_137 | v_179 | v_163 | v_162 | v_161 | v_182 | ~v_361 | ~v_360 | ~v_357 | ~v_356 | ~v_315 | ~v_314 | ~v_355 | ~v_354 | ~v_3288 | ~v_3285 | ~v_3344 | ~v_3343 | ~v_3342 | ~v_3341 | ~v_3428 | ~v_3427 | ~v_3426 | ~v_3425 | ~v_3808 | ~v_3807 | ~v_223 | ~v_3806 | ~v_3805 | ~v_220 | ~v_353 | ~v_352 | ~v_351 | ~v_350 | ~v_309 | ~v_308 | ~v_307 | ~v_306 | v_3825;
assign x_7326 = v_3824 | ~v_3821;
assign x_7327 = v_3824 | ~v_3822;
assign x_7328 = v_3824 | ~v_3823;
assign x_7329 = v_103 | v_95 | v_102 | v_171 | v_170 | v_169 | v_160 | v_150 | v_149 | v_148 | v_184 | v_181 | ~v_297 | ~v_296 | ~v_345 | ~v_344 | ~v_343 | ~v_342 | ~v_341 | ~v_340 | ~v_3318 | ~v_3315 | ~v_3370 | ~v_3369 | ~v_3368 | ~v_3367 | ~v_3438 | ~v_3437 | ~v_3436 | ~v_3435 | ~v_3818 | ~v_3817 | ~v_289 | ~v_3816 | ~v_3815 | ~v_286 | ~v_285 | ~v_284 | ~v_283 | ~v_282 | ~v_339 | ~v_338 | ~v_337 | ~v_336 | v_3823;
assign x_7330 = v_53 | v_61 | v_60 | v_144 | v_180 | v_159 | v_145 | v_143 | v_167 | v_166 | v_165 | v_183 | ~v_264 | ~v_263 | ~v_330 | ~v_329 | ~v_328 | ~v_327 | ~v_326 | ~v_325 | ~v_3303 | ~v_3300 | ~v_3365 | ~v_3364 | ~v_3363 | ~v_3362 | ~v_3433 | ~v_3432 | ~v_3431 | ~v_3430 | ~v_3813 | ~v_3812 | ~v_256 | ~v_3811 | ~v_3810 | ~v_253 | ~v_252 | ~v_251 | ~v_250 | ~v_249 | ~v_324 | ~v_323 | ~v_322 | ~v_321 | v_3822;
assign x_7331 = v_18 | v_17 | v_10 | v_136 | v_135 | v_137 | v_179 | v_163 | v_162 | v_161 | v_155 | v_182 | ~v_231 | ~v_230 | ~v_315 | ~v_314 | ~v_313 | ~v_312 | ~v_311 | ~v_310 | ~v_3288 | ~v_3285 | ~v_3360 | ~v_3359 | ~v_3358 | ~v_3357 | ~v_3428 | ~v_3427 | ~v_3426 | ~v_3425 | ~v_3808 | ~v_3807 | ~v_223 | ~v_3806 | ~v_3805 | ~v_220 | ~v_219 | ~v_218 | ~v_217 | ~v_216 | ~v_309 | ~v_308 | ~v_307 | ~v_306 | v_3821;
assign x_7332 = v_3820 | ~v_3809;
assign x_7333 = v_3820 | ~v_3814;
assign x_7334 = v_3820 | ~v_3819;
assign x_7335 = v_98 | v_103 | v_100 | v_94 | v_102 | v_169 | v_160 | v_150 | v_149 | v_148 | v_147 | v_184 | ~v_299 | ~v_298 | ~v_297 | ~v_296 | ~v_295 | ~v_294 | ~v_293 | ~v_292 | ~v_3320 | ~v_3319 | ~v_3318 | ~v_3317 | ~v_3316 | ~v_3315 | ~v_3370 | ~v_3369 | ~v_3368 | ~v_3367 | ~v_291 | ~v_3818 | ~v_290 | ~v_3817 | ~v_289 | ~v_288 | ~v_3816 | ~v_287 | ~v_3815 | ~v_286 | ~v_285 | ~v_284 | ~v_283 | ~v_282 | v_3819;
assign x_7336 = v_3818 | v_152;
assign x_7337 = v_3818 | v_123;
assign x_7338 = v_3817 | v_153;
assign x_7339 = v_3817 | v_120;
assign x_7340 = v_3816 | ~v_152;
assign x_7341 = v_3816 | v_108;
assign x_7342 = v_3815 | ~v_153;
assign x_7343 = v_3815 | v_105;
assign x_7344 = v_56 | v_61 | v_52 | v_60 | v_58 | v_144 | v_159 | v_145 | v_143 | v_142 | v_165 | v_183 | ~v_3305 | ~v_266 | ~v_265 | ~v_264 | ~v_263 | ~v_262 | ~v_261 | ~v_260 | ~v_259 | ~v_3304 | ~v_3303 | ~v_3302 | ~v_3301 | ~v_3300 | ~v_3365 | ~v_3364 | ~v_3363 | ~v_3362 | ~v_258 | ~v_3813 | ~v_257 | ~v_3812 | ~v_256 | ~v_255 | ~v_3811 | ~v_254 | ~v_3810 | ~v_253 | ~v_252 | ~v_251 | ~v_250 | ~v_249 | v_3814;
assign x_7345 = v_3813 | v_152;
assign x_7346 = v_3813 | v_81;
assign x_7347 = v_3812 | v_153;
assign x_7348 = v_3812 | v_78;
assign x_7349 = v_3811 | ~v_152;
assign x_7350 = v_3811 | v_66;
assign x_7351 = v_3810 | ~v_153;
assign x_7352 = v_3810 | v_63;
assign x_7353 = v_13 | v_9 | v_18 | v_17 | v_15 | v_136 | v_135 | v_134 | ~v_3292 | v_137 | v_161 | v_155 | v_182 | ~v_233 | ~v_232 | ~v_231 | ~v_230 | ~v_229 | ~v_228 | ~v_227 | ~v_226 | ~v_3289 | ~v_3288 | ~v_3287 | ~v_3286 | ~v_3285 | ~v_3360 | ~v_3359 | ~v_3358 | ~v_3357 | ~v_225 | ~v_3808 | ~v_224 | ~v_3807 | ~v_223 | ~v_222 | ~v_3806 | ~v_221 | ~v_3805 | ~v_220 | ~v_219 | ~v_218 | ~v_217 | ~v_216 | v_3809;
assign x_7354 = v_3808 | v_152;
assign x_7355 = v_3808 | v_39;
assign x_7356 = v_3807 | v_153;
assign x_7357 = v_3807 | v_36;
assign x_7358 = v_3806 | ~v_152;
assign x_7359 = v_3806 | v_24;
assign x_7360 = v_3805 | ~v_153;
assign x_7361 = v_3805 | v_21;
assign x_7362 = v_3804 | ~v_3802;
assign x_7363 = v_3804 | ~v_3803;
assign x_7364 = v_3804 | ~v_1274;
assign x_7365 = v_3804 | ~v_1275;
assign x_7366 = v_3804 | ~v_153;
assign x_7367 = v_3804 | ~v_152;
assign x_7368 = ~v_189 | ~v_2221 | v_3803;
assign x_7369 = ~v_188 | ~v_197 | v_3802;
assign x_7370 = v_3801 | ~v_3720;
assign x_7371 = v_3801 | ~v_3800;
assign x_7372 = v_152 | v_153 | ~v_3799 | ~v_1565 | ~v_1564 | ~v_3722 | ~v_3721 | v_3800;
assign x_7373 = v_3799 | ~v_3738;
assign x_7374 = v_3799 | ~v_3742;
assign x_7375 = v_3799 | ~v_3746;
assign x_7376 = v_3799 | ~v_3750;
assign x_7377 = v_3799 | ~v_3754;
assign x_7378 = v_3799 | ~v_3758;
assign x_7379 = v_3799 | ~v_3762;
assign x_7380 = v_3799 | ~v_3766;
assign x_7381 = v_3799 | ~v_3770;
assign x_7382 = v_3799 | ~v_3774;
assign x_7383 = v_3799 | ~v_3778;
assign x_7384 = v_3799 | ~v_3782;
assign x_7385 = v_3799 | ~v_3786;
assign x_7386 = v_3799 | ~v_3790;
assign x_7387 = v_3799 | ~v_3794;
assign x_7388 = v_3799 | ~v_3798;
assign x_7389 = v_3799 | ~v_1263;
assign x_7390 = v_3799 | ~v_1264;
assign x_7391 = v_3799 | ~v_1265;
assign x_7392 = v_3799 | ~v_1266;
assign x_7393 = ~v_3797 | ~v_3796 | ~v_3795 | v_3798;
assign x_7394 = v_3797 | ~v_3733;
assign x_7395 = v_3797 | ~v_3734;
assign x_7396 = v_3797 | ~v_1636;
assign x_7397 = v_3797 | ~v_1637;
assign x_7398 = v_3797 | ~v_1750;
assign x_7399 = v_3797 | ~v_1638;
assign x_7400 = v_3797 | ~v_1751;
assign x_7401 = v_3797 | ~v_3735;
assign x_7402 = v_3797 | ~v_3736;
assign x_7403 = v_3797 | ~v_1639;
assign x_7404 = v_3797 | ~v_1640;
assign x_7405 = v_3797 | ~v_1752;
assign x_7406 = v_3797 | ~v_1641;
assign x_7407 = v_3797 | ~v_1753;
assign x_7408 = v_3797 | ~v_3133;
assign x_7409 = v_3797 | ~v_3134;
assign x_7410 = v_3797 | ~v_3199;
assign x_7411 = v_3797 | ~v_3135;
assign x_7412 = v_3797 | ~v_839;
assign x_7413 = v_3797 | ~v_3200;
assign x_7414 = v_3797 | ~v_1257;
assign x_7415 = v_3797 | ~v_1023;
assign x_7416 = v_3797 | ~v_3136;
assign x_7417 = v_3797 | ~v_3137;
assign x_7418 = v_3797 | ~v_3201;
assign x_7419 = v_3797 | ~v_3138;
assign x_7420 = v_3797 | ~v_840;
assign x_7421 = v_3797 | ~v_3202;
assign x_7422 = v_3797 | ~v_1258;
assign x_7423 = v_3797 | ~v_1024;
assign x_7424 = v_3797 | ~v_184;
assign x_7425 = v_3797 | ~v_170;
assign x_7426 = v_3797 | ~v_149;
assign x_7427 = v_3797 | ~v_1259;
assign x_7428 = v_3797 | ~v_1260;
assign x_7429 = v_3797 | ~v_103;
assign x_7430 = v_3797 | ~v_102;
assign x_7431 = v_3797 | ~v_101;
assign x_7432 = v_3797 | ~v_100;
assign x_7433 = v_3797 | ~v_99;
assign x_7434 = v_3797 | ~v_98;
assign x_7435 = v_3797 | ~v_96;
assign x_7436 = v_3797 | ~v_95;
assign x_7437 = v_3797 | ~v_93;
assign x_7438 = v_3796 | ~v_3728;
assign x_7439 = v_3796 | ~v_3729;
assign x_7440 = v_3796 | ~v_1611;
assign x_7441 = v_3796 | ~v_1612;
assign x_7442 = v_3796 | ~v_1741;
assign x_7443 = v_3796 | ~v_1613;
assign x_7444 = v_3796 | ~v_1742;
assign x_7445 = v_3796 | ~v_3730;
assign x_7446 = v_3796 | ~v_3731;
assign x_7447 = v_3796 | ~v_1614;
assign x_7448 = v_3796 | ~v_1615;
assign x_7449 = v_3796 | ~v_1743;
assign x_7450 = v_3796 | ~v_1616;
assign x_7451 = v_3796 | ~v_1744;
assign x_7452 = v_3796 | ~v_3118;
assign x_7453 = v_3796 | ~v_3119;
assign x_7454 = v_3796 | ~v_3194;
assign x_7455 = v_3796 | ~v_3120;
assign x_7456 = v_3796 | ~v_806;
assign x_7457 = v_3796 | ~v_3195;
assign x_7458 = v_3796 | ~v_1252;
assign x_7459 = v_3796 | ~v_1008;
assign x_7460 = v_3796 | ~v_3121;
assign x_7461 = v_3796 | ~v_3122;
assign x_7462 = v_3796 | ~v_1253;
assign x_7463 = v_3796 | ~v_1009;
assign x_7464 = v_3796 | ~v_3123;
assign x_7465 = v_3796 | ~v_807;
assign x_7466 = v_3796 | ~v_3196;
assign x_7467 = v_3796 | ~v_183;
assign x_7468 = v_3796 | ~v_166;
assign x_7469 = v_3796 | ~v_144;
assign x_7470 = v_3796 | ~v_3197;
assign x_7471 = v_3796 | ~v_1254;
assign x_7472 = v_3796 | ~v_1255;
assign x_7473 = v_3796 | ~v_61;
assign x_7474 = v_3796 | ~v_60;
assign x_7475 = v_3796 | ~v_59;
assign x_7476 = v_3796 | ~v_58;
assign x_7477 = v_3796 | ~v_57;
assign x_7478 = v_3796 | ~v_56;
assign x_7479 = v_3796 | ~v_54;
assign x_7480 = v_3796 | ~v_53;
assign x_7481 = v_3796 | ~v_51;
assign x_7482 = v_3795 | ~v_3723;
assign x_7483 = v_3795 | ~v_3724;
assign x_7484 = v_3795 | ~v_1586;
assign x_7485 = v_3795 | ~v_1587;
assign x_7486 = v_3795 | ~v_1732;
assign x_7487 = v_3795 | ~v_1588;
assign x_7488 = v_3795 | ~v_1733;
assign x_7489 = v_3795 | ~v_3725;
assign x_7490 = v_3795 | ~v_3726;
assign x_7491 = v_3795 | ~v_1589;
assign x_7492 = v_3795 | ~v_1590;
assign x_7493 = v_3795 | ~v_1734;
assign x_7494 = v_3795 | ~v_1591;
assign x_7495 = v_3795 | ~v_1735;
assign x_7496 = v_3795 | ~v_3103;
assign x_7497 = v_3795 | ~v_3189;
assign x_7498 = v_3795 | ~v_3104;
assign x_7499 = v_3795 | ~v_773;
assign x_7500 = v_3795 | ~v_3190;
assign x_7501 = v_3795 | ~v_3105;
assign x_7502 = v_3795 | ~v_3191;
assign x_7503 = v_3795 | ~v_3106;
assign x_7504 = v_3795 | ~v_774;
assign x_7505 = v_3795 | ~v_3192;
assign x_7506 = v_3795 | ~v_182;
assign x_7507 = v_3795 | ~v_162;
assign x_7508 = v_3795 | ~v_1247;
assign x_7509 = v_3795 | ~v_1248;
assign x_7510 = v_3795 | ~v_136;
assign x_7511 = v_3795 | ~v_3107;
assign x_7512 = v_3795 | ~v_1249;
assign x_7513 = v_3795 | ~v_993;
assign x_7514 = v_3795 | ~v_3108;
assign x_7515 = v_3795 | ~v_1250;
assign x_7516 = v_3795 | ~v_994;
assign x_7517 = v_3795 | ~v_18;
assign x_7518 = v_3795 | ~v_17;
assign x_7519 = v_3795 | ~v_16;
assign x_7520 = v_3795 | ~v_15;
assign x_7521 = v_3795 | ~v_14;
assign x_7522 = v_3795 | ~v_13;
assign x_7523 = v_3795 | ~v_11;
assign x_7524 = v_3795 | ~v_10;
assign x_7525 = v_3795 | ~v_8;
assign x_7526 = ~v_3793 | ~v_3792 | ~v_3791 | v_3794;
assign x_7527 = v_3793 | ~v_1666;
assign x_7528 = v_3793 | ~v_1667;
assign x_7529 = v_3793 | ~v_1668;
assign x_7530 = v_3793 | ~v_1669;
assign x_7531 = v_3793 | ~v_3733;
assign x_7532 = v_3793 | ~v_3734;
assign x_7533 = v_3793 | ~v_1636;
assign x_7534 = v_3793 | ~v_1750;
assign x_7535 = v_3793 | ~v_1751;
assign x_7536 = v_3793 | ~v_3735;
assign x_7537 = v_3793 | ~v_3736;
assign x_7538 = v_3793 | ~v_1639;
assign x_7539 = v_3793 | ~v_1752;
assign x_7540 = v_3793 | ~v_1753;
assign x_7541 = v_3793 | ~v_3151;
assign x_7542 = v_3793 | ~v_3152;
assign x_7543 = v_3793 | ~v_1193;
assign x_7544 = v_3793 | ~v_1241;
assign x_7545 = v_3793 | ~v_3153;
assign x_7546 = v_3793 | ~v_3154;
assign x_7547 = v_3793 | ~v_1194;
assign x_7548 = v_3793 | ~v_1242;
assign x_7549 = v_3793 | ~v_3133;
assign x_7550 = v_3793 | ~v_3199;
assign x_7551 = v_3793 | ~v_3200;
assign x_7552 = v_3793 | ~v_1023;
assign x_7553 = v_3793 | ~v_3136;
assign x_7554 = v_3793 | ~v_3201;
assign x_7555 = v_3793 | ~v_3202;
assign x_7556 = v_3793 | ~v_1024;
assign x_7557 = v_3793 | ~v_1243;
assign x_7558 = v_3793 | ~v_1244;
assign x_7559 = v_3793 | ~v_184;
assign x_7560 = v_3793 | ~v_171;
assign x_7561 = v_3793 | ~v_169;
assign x_7562 = v_3793 | ~v_149;
assign x_7563 = v_3793 | ~v_147;
assign x_7564 = v_3793 | ~v_103;
assign x_7565 = v_3793 | ~v_102;
assign x_7566 = v_3793 | ~v_101;
assign x_7567 = v_3793 | ~v_100;
assign x_7568 = v_3793 | ~v_99;
assign x_7569 = v_3793 | ~v_96;
assign x_7570 = v_3793 | ~v_94;
assign x_7571 = v_3792 | ~v_1657;
assign x_7572 = v_3792 | ~v_1658;
assign x_7573 = v_3792 | ~v_1659;
assign x_7574 = v_3792 | ~v_1660;
assign x_7575 = v_3792 | ~v_3728;
assign x_7576 = v_3792 | ~v_3729;
assign x_7577 = v_3792 | ~v_1611;
assign x_7578 = v_3792 | ~v_1741;
assign x_7579 = v_3792 | ~v_1742;
assign x_7580 = v_3792 | ~v_3730;
assign x_7581 = v_3792 | ~v_3731;
assign x_7582 = v_3792 | ~v_1614;
assign x_7583 = v_3792 | ~v_1743;
assign x_7584 = v_3792 | ~v_1744;
assign x_7585 = v_3792 | ~v_3146;
assign x_7586 = v_3792 | ~v_3147;
assign x_7587 = v_3792 | ~v_1178;
assign x_7588 = v_3792 | ~v_1236;
assign x_7589 = v_3792 | ~v_3148;
assign x_7590 = v_3792 | ~v_3149;
assign x_7591 = v_3792 | ~v_1179;
assign x_7592 = v_3792 | ~v_1237;
assign x_7593 = v_3792 | ~v_3118;
assign x_7594 = v_3792 | ~v_3194;
assign x_7595 = v_3792 | ~v_3195;
assign x_7596 = v_3792 | ~v_1008;
assign x_7597 = v_3792 | ~v_3121;
assign x_7598 = v_3792 | ~v_1009;
assign x_7599 = v_3792 | ~v_3196;
assign x_7600 = v_3792 | ~v_1238;
assign x_7601 = v_3792 | ~v_1239;
assign x_7602 = v_3792 | ~v_183;
assign x_7603 = v_3792 | ~v_167;
assign x_7604 = v_3792 | ~v_165;
assign x_7605 = v_3792 | ~v_144;
assign x_7606 = v_3792 | ~v_142;
assign x_7607 = v_3792 | ~v_3197;
assign x_7608 = v_3792 | ~v_61;
assign x_7609 = v_3792 | ~v_60;
assign x_7610 = v_3792 | ~v_59;
assign x_7611 = v_3792 | ~v_58;
assign x_7612 = v_3792 | ~v_57;
assign x_7613 = v_3792 | ~v_54;
assign x_7614 = v_3792 | ~v_52;
assign x_7615 = v_3791 | ~v_1648;
assign x_7616 = v_3791 | ~v_1649;
assign x_7617 = v_3791 | ~v_1650;
assign x_7618 = v_3791 | ~v_1651;
assign x_7619 = v_3791 | ~v_3723;
assign x_7620 = v_3791 | ~v_3724;
assign x_7621 = v_3791 | ~v_1586;
assign x_7622 = v_3791 | ~v_1732;
assign x_7623 = v_3791 | ~v_1733;
assign x_7624 = v_3791 | ~v_3725;
assign x_7625 = v_3791 | ~v_3726;
assign x_7626 = v_3791 | ~v_1589;
assign x_7627 = v_3791 | ~v_1734;
assign x_7628 = v_3791 | ~v_1735;
assign x_7629 = v_3791 | ~v_3141;
assign x_7630 = v_3791 | ~v_3142;
assign x_7631 = v_3791 | ~v_1163;
assign x_7632 = v_3791 | ~v_1231;
assign x_7633 = v_3791 | ~v_3143;
assign x_7634 = v_3791 | ~v_3144;
assign x_7635 = v_3791 | ~v_1164;
assign x_7636 = v_3791 | ~v_1232;
assign x_7637 = v_3791 | ~v_3189;
assign x_7638 = v_3791 | ~v_3190;
assign x_7639 = v_3791 | ~v_3191;
assign x_7640 = v_3791 | ~v_3192;
assign x_7641 = v_3791 | ~v_1233;
assign x_7642 = v_3791 | ~v_1234;
assign x_7643 = v_3791 | ~v_182;
assign x_7644 = v_3791 | ~v_163;
assign x_7645 = v_3791 | ~v_161;
assign x_7646 = v_3791 | ~v_136;
assign x_7647 = v_3791 | ~v_134;
assign x_7648 = v_3791 | ~v_3107;
assign x_7649 = v_3791 | ~v_993;
assign x_7650 = v_3791 | ~v_3108;
assign x_7651 = v_3791 | ~v_994;
assign x_7652 = v_3791 | ~v_18;
assign x_7653 = v_3791 | ~v_17;
assign x_7654 = v_3791 | ~v_16;
assign x_7655 = v_3791 | ~v_15;
assign x_7656 = v_3791 | ~v_14;
assign x_7657 = v_3791 | ~v_11;
assign x_7658 = v_3791 | ~v_9;
assign x_7659 = ~v_3789 | ~v_3788 | ~v_3787 | v_3790;
assign x_7660 = v_3789 | ~v_1632;
assign x_7661 = v_3789 | ~v_1633;
assign x_7662 = v_3789 | ~v_1634;
assign x_7663 = v_3789 | ~v_1635;
assign x_7664 = v_3789 | ~v_1666;
assign x_7665 = v_3789 | ~v_1667;
assign x_7666 = v_3789 | ~v_1668;
assign x_7667 = v_3789 | ~v_1669;
assign x_7668 = v_3789 | ~v_3733;
assign x_7669 = v_3789 | ~v_3734;
assign x_7670 = v_3789 | ~v_1636;
assign x_7671 = v_3789 | ~v_3735;
assign x_7672 = v_3789 | ~v_3736;
assign x_7673 = v_3789 | ~v_1639;
assign x_7674 = v_3789 | ~v_1225;
assign x_7675 = v_3789 | ~v_1226;
assign x_7676 = v_3789 | ~v_1227;
assign x_7677 = v_3789 | ~v_1228;
assign x_7678 = v_3789 | ~v_3151;
assign x_7679 = v_3789 | ~v_3152;
assign x_7680 = v_3789 | ~v_1193;
assign x_7681 = v_3789 | ~v_3153;
assign x_7682 = v_3789 | ~v_3154;
assign x_7683 = v_3789 | ~v_1194;
assign x_7684 = v_3789 | ~v_3129;
assign x_7685 = v_3789 | ~v_3130;
assign x_7686 = v_3789 | ~v_975;
assign x_7687 = v_3789 | ~v_3131;
assign x_7688 = v_3789 | ~v_3132;
assign x_7689 = v_3789 | ~v_976;
assign x_7690 = v_3789 | ~v_3133;
assign x_7691 = v_3789 | ~v_3136;
assign x_7692 = v_3789 | ~v_184;
assign x_7693 = v_3789 | ~v_171;
assign x_7694 = v_3789 | ~v_169;
assign x_7695 = v_3789 | ~v_150;
assign x_7696 = v_3789 | ~v_148;
assign x_7697 = v_3789 | ~v_103;
assign x_7698 = v_3789 | ~v_102;
assign x_7699 = v_3789 | ~v_101;
assign x_7700 = v_3789 | ~v_100;
assign x_7701 = v_3789 | ~v_97;
assign x_7702 = v_3789 | ~v_95;
assign x_7703 = v_3789 | ~v_94;
assign x_7704 = v_3788 | ~v_1607;
assign x_7705 = v_3788 | ~v_1608;
assign x_7706 = v_3788 | ~v_1609;
assign x_7707 = v_3788 | ~v_1610;
assign x_7708 = v_3788 | ~v_1657;
assign x_7709 = v_3788 | ~v_1658;
assign x_7710 = v_3788 | ~v_1659;
assign x_7711 = v_3788 | ~v_1660;
assign x_7712 = v_3788 | ~v_3728;
assign x_7713 = v_3788 | ~v_3729;
assign x_7714 = v_3788 | ~v_1611;
assign x_7715 = v_3788 | ~v_3730;
assign x_7716 = v_3788 | ~v_3731;
assign x_7717 = v_3788 | ~v_1614;
assign x_7718 = v_3788 | ~v_1220;
assign x_7719 = v_3788 | ~v_1221;
assign x_7720 = v_3788 | ~v_1222;
assign x_7721 = v_3788 | ~v_1223;
assign x_7722 = v_3788 | ~v_3146;
assign x_7723 = v_3788 | ~v_3147;
assign x_7724 = v_3788 | ~v_1178;
assign x_7725 = v_3788 | ~v_3148;
assign x_7726 = v_3788 | ~v_3149;
assign x_7727 = v_3788 | ~v_1179;
assign x_7728 = v_3788 | ~v_3114;
assign x_7729 = v_3788 | ~v_3115;
assign x_7730 = v_3788 | ~v_960;
assign x_7731 = v_3788 | ~v_3116;
assign x_7732 = v_3788 | ~v_3117;
assign x_7733 = v_3788 | ~v_961;
assign x_7734 = v_3788 | ~v_3118;
assign x_7735 = v_3788 | ~v_3121;
assign x_7736 = v_3788 | ~v_183;
assign x_7737 = v_3788 | ~v_167;
assign x_7738 = v_3788 | ~v_165;
assign x_7739 = v_3788 | ~v_145;
assign x_7740 = v_3788 | ~v_143;
assign x_7741 = v_3788 | ~v_61;
assign x_7742 = v_3788 | ~v_60;
assign x_7743 = v_3788 | ~v_59;
assign x_7744 = v_3788 | ~v_58;
assign x_7745 = v_3788 | ~v_55;
assign x_7746 = v_3788 | ~v_53;
assign x_7747 = v_3788 | ~v_52;
assign x_7748 = v_3787 | ~v_1582;
assign x_7749 = v_3787 | ~v_1583;
assign x_7750 = v_3787 | ~v_1584;
assign x_7751 = v_3787 | ~v_1585;
assign x_7752 = v_3787 | ~v_1648;
assign x_7753 = v_3787 | ~v_1649;
assign x_7754 = v_3787 | ~v_1650;
assign x_7755 = v_3787 | ~v_1651;
assign x_7756 = v_3787 | ~v_3723;
assign x_7757 = v_3787 | ~v_3724;
assign x_7758 = v_3787 | ~v_1586;
assign x_7759 = v_3787 | ~v_3725;
assign x_7760 = v_3787 | ~v_3726;
assign x_7761 = v_3787 | ~v_1589;
assign x_7762 = v_3787 | ~v_1215;
assign x_7763 = v_3787 | ~v_1216;
assign x_7764 = v_3787 | ~v_1217;
assign x_7765 = v_3787 | ~v_1218;
assign x_7766 = v_3787 | ~v_3141;
assign x_7767 = v_3787 | ~v_3142;
assign x_7768 = v_3787 | ~v_1163;
assign x_7769 = v_3787 | ~v_3143;
assign x_7770 = v_3787 | ~v_3144;
assign x_7771 = v_3787 | ~v_1164;
assign x_7772 = v_3787 | ~v_3099;
assign x_7773 = v_3787 | ~v_3100;
assign x_7774 = v_3787 | ~v_945;
assign x_7775 = v_3787 | ~v_3101;
assign x_7776 = v_3787 | ~v_3102;
assign x_7777 = v_3787 | ~v_946;
assign x_7778 = v_3787 | ~v_182;
assign x_7779 = v_3787 | ~v_163;
assign x_7780 = v_3787 | ~v_161;
assign x_7781 = v_3787 | ~v_137;
assign x_7782 = v_3787 | ~v_135;
assign x_7783 = v_3787 | ~v_3107;
assign x_7784 = v_3787 | ~v_3108;
assign x_7785 = v_3787 | ~v_18;
assign x_7786 = v_3787 | ~v_17;
assign x_7787 = v_3787 | ~v_16;
assign x_7788 = v_3787 | ~v_15;
assign x_7789 = v_3787 | ~v_12;
assign x_7790 = v_3787 | ~v_10;
assign x_7791 = v_3787 | ~v_9;
assign x_7792 = ~v_3785 | ~v_3784 | ~v_3783 | v_3786;
assign x_7793 = v_3785 | ~v_1694;
assign x_7794 = v_3785 | ~v_1695;
assign x_7795 = v_3785 | ~v_1696;
assign x_7796 = v_3785 | ~v_1697;
assign x_7797 = v_3785 | ~v_1666;
assign x_7798 = v_3785 | ~v_1667;
assign x_7799 = v_3785 | ~v_1668;
assign x_7800 = v_3785 | ~v_1669;
assign x_7801 = v_3785 | ~v_3733;
assign x_7802 = v_3785 | ~v_3734;
assign x_7803 = v_3785 | ~v_1636;
assign x_7804 = v_3785 | ~v_3735;
assign x_7805 = v_3785 | ~v_3736;
assign x_7806 = v_3785 | ~v_1639;
assign x_7807 = v_3785 | ~v_1209;
assign x_7808 = v_3785 | ~v_1210;
assign x_7809 = v_3785 | ~v_3151;
assign x_7810 = v_3785 | ~v_3152;
assign x_7811 = v_3785 | ~v_1193;
assign x_7812 = v_3785 | ~v_3153;
assign x_7813 = v_3785 | ~v_3154;
assign x_7814 = v_3785 | ~v_1194;
assign x_7815 = v_3785 | ~v_3167;
assign x_7816 = v_3785 | ~v_3168;
assign x_7817 = v_3785 | ~v_927;
assign x_7818 = v_3785 | ~v_3169;
assign x_7819 = v_3785 | ~v_3170;
assign x_7820 = v_3785 | ~v_928;
assign x_7821 = v_3785 | ~v_3133;
assign x_7822 = v_3785 | ~v_3136;
assign x_7823 = v_3785 | ~v_1211;
assign x_7824 = v_3785 | ~v_1212;
assign x_7825 = v_3785 | ~v_184;
assign x_7826 = v_3785 | ~v_172;
assign x_7827 = v_3785 | ~v_171;
assign x_7828 = v_3785 | ~v_169;
assign x_7829 = v_3785 | ~v_150;
assign x_7830 = v_3785 | ~v_149;
assign x_7831 = v_3785 | ~v_148;
assign x_7832 = v_3785 | ~v_147;
assign x_7833 = v_3785 | ~v_102;
assign x_7834 = v_3785 | ~v_101;
assign x_7835 = v_3785 | ~v_100;
assign x_7836 = v_3785 | ~v_94;
assign x_7837 = v_3784 | ~v_1685;
assign x_7838 = v_3784 | ~v_1686;
assign x_7839 = v_3784 | ~v_1687;
assign x_7840 = v_3784 | ~v_1688;
assign x_7841 = v_3784 | ~v_1657;
assign x_7842 = v_3784 | ~v_1658;
assign x_7843 = v_3784 | ~v_1659;
assign x_7844 = v_3784 | ~v_1660;
assign x_7845 = v_3784 | ~v_3728;
assign x_7846 = v_3784 | ~v_3729;
assign x_7847 = v_3784 | ~v_1611;
assign x_7848 = v_3784 | ~v_3730;
assign x_7849 = v_3784 | ~v_3731;
assign x_7850 = v_3784 | ~v_1614;
assign x_7851 = v_3784 | ~v_1204;
assign x_7852 = v_3784 | ~v_1205;
assign x_7853 = v_3784 | ~v_3146;
assign x_7854 = v_3784 | ~v_3147;
assign x_7855 = v_3784 | ~v_1178;
assign x_7856 = v_3784 | ~v_3148;
assign x_7857 = v_3784 | ~v_3149;
assign x_7858 = v_3784 | ~v_1179;
assign x_7859 = v_3784 | ~v_3162;
assign x_7860 = v_3784 | ~v_3163;
assign x_7861 = v_3784 | ~v_912;
assign x_7862 = v_3784 | ~v_3164;
assign x_7863 = v_3784 | ~v_3165;
assign x_7864 = v_3784 | ~v_913;
assign x_7865 = v_3784 | ~v_3118;
assign x_7866 = v_3784 | ~v_3121;
assign x_7867 = v_3784 | ~v_1206;
assign x_7868 = v_3784 | ~v_1207;
assign x_7869 = v_3784 | ~v_183;
assign x_7870 = v_3784 | ~v_168;
assign x_7871 = v_3784 | ~v_167;
assign x_7872 = v_3784 | ~v_165;
assign x_7873 = v_3784 | ~v_145;
assign x_7874 = v_3784 | ~v_144;
assign x_7875 = v_3784 | ~v_143;
assign x_7876 = v_3784 | ~v_142;
assign x_7877 = v_3784 | ~v_60;
assign x_7878 = v_3784 | ~v_59;
assign x_7879 = v_3784 | ~v_58;
assign x_7880 = v_3784 | ~v_52;
assign x_7881 = v_3783 | ~v_1676;
assign x_7882 = v_3783 | ~v_1677;
assign x_7883 = v_3783 | ~v_1678;
assign x_7884 = v_3783 | ~v_1679;
assign x_7885 = v_3783 | ~v_1648;
assign x_7886 = v_3783 | ~v_1649;
assign x_7887 = v_3783 | ~v_1650;
assign x_7888 = v_3783 | ~v_1651;
assign x_7889 = v_3783 | ~v_3723;
assign x_7890 = v_3783 | ~v_3724;
assign x_7891 = v_3783 | ~v_1586;
assign x_7892 = v_3783 | ~v_3725;
assign x_7893 = v_3783 | ~v_3726;
assign x_7894 = v_3783 | ~v_1589;
assign x_7895 = v_3783 | ~v_1199;
assign x_7896 = v_3783 | ~v_1200;
assign x_7897 = v_3783 | ~v_3141;
assign x_7898 = v_3783 | ~v_3142;
assign x_7899 = v_3783 | ~v_1163;
assign x_7900 = v_3783 | ~v_3143;
assign x_7901 = v_3783 | ~v_3144;
assign x_7902 = v_3783 | ~v_1164;
assign x_7903 = v_3783 | ~v_3157;
assign x_7904 = v_3783 | ~v_3158;
assign x_7905 = v_3783 | ~v_897;
assign x_7906 = v_3783 | ~v_3159;
assign x_7907 = v_3783 | ~v_3160;
assign x_7908 = v_3783 | ~v_898;
assign x_7909 = v_3783 | ~v_1201;
assign x_7910 = v_3783 | ~v_1202;
assign x_7911 = v_3783 | ~v_182;
assign x_7912 = v_3783 | ~v_164;
assign x_7913 = v_3783 | ~v_163;
assign x_7914 = v_3783 | ~v_161;
assign x_7915 = v_3783 | ~v_137;
assign x_7916 = v_3783 | ~v_136;
assign x_7917 = v_3783 | ~v_135;
assign x_7918 = v_3783 | ~v_134;
assign x_7919 = v_3783 | ~v_3107;
assign x_7920 = v_3783 | ~v_3108;
assign x_7921 = v_3783 | ~v_17;
assign x_7922 = v_3783 | ~v_16;
assign x_7923 = v_3783 | ~v_15;
assign x_7924 = v_3783 | ~v_9;
assign x_7925 = ~v_3781 | ~v_3780 | ~v_3779 | v_3782;
assign x_7926 = v_3781 | ~v_1722;
assign x_7927 = v_3781 | ~v_1723;
assign x_7928 = v_3781 | ~v_1724;
assign x_7929 = v_3781 | ~v_1725;
assign x_7930 = v_3781 | ~v_1666;
assign x_7931 = v_3781 | ~v_1667;
assign x_7932 = v_3781 | ~v_1668;
assign x_7933 = v_3781 | ~v_1669;
assign x_7934 = v_3781 | ~v_3733;
assign x_7935 = v_3781 | ~v_3734;
assign x_7936 = v_3781 | ~v_1636;
assign x_7937 = v_3781 | ~v_3735;
assign x_7938 = v_3781 | ~v_3736;
assign x_7939 = v_3781 | ~v_1639;
assign x_7940 = v_3781 | ~v_1191;
assign x_7941 = v_3781 | ~v_1192;
assign x_7942 = v_3781 | ~v_3151;
assign x_7943 = v_3781 | ~v_3152;
assign x_7944 = v_3781 | ~v_1193;
assign x_7945 = v_3781 | ~v_3153;
assign x_7946 = v_3781 | ~v_3154;
assign x_7947 = v_3781 | ~v_1194;
assign x_7948 = v_3781 | ~v_3183;
assign x_7949 = v_3781 | ~v_3184;
assign x_7950 = v_3781 | ~v_837;
assign x_7951 = v_3781 | ~v_3185;
assign x_7952 = v_3781 | ~v_3186;
assign x_7953 = v_3781 | ~v_838;
assign x_7954 = v_3781 | ~v_3133;
assign x_7955 = v_3781 | ~v_3136;
assign x_7956 = v_3781 | ~v_1195;
assign x_7957 = v_3781 | ~v_1196;
assign x_7958 = v_3781 | ~v_184;
assign x_7959 = v_3781 | ~v_171;
assign x_7960 = v_3781 | ~v_169;
assign x_7961 = v_3781 | ~v_160;
assign x_7962 = v_3781 | ~v_151;
assign x_7963 = v_3781 | ~v_150;
assign x_7964 = v_3781 | ~v_149;
assign x_7965 = v_3781 | ~v_148;
assign x_7966 = v_3781 | ~v_147;
assign x_7967 = v_3781 | ~v_103;
assign x_7968 = v_3781 | ~v_100;
assign x_7969 = v_3781 | ~v_94;
assign x_7970 = v_3780 | ~v_1713;
assign x_7971 = v_3780 | ~v_1714;
assign x_7972 = v_3780 | ~v_1715;
assign x_7973 = v_3780 | ~v_1716;
assign x_7974 = v_3780 | ~v_1657;
assign x_7975 = v_3780 | ~v_1658;
assign x_7976 = v_3780 | ~v_1659;
assign x_7977 = v_3780 | ~v_1660;
assign x_7978 = v_3780 | ~v_3728;
assign x_7979 = v_3780 | ~v_3729;
assign x_7980 = v_3780 | ~v_1611;
assign x_7981 = v_3780 | ~v_3730;
assign x_7982 = v_3780 | ~v_3731;
assign x_7983 = v_3780 | ~v_1614;
assign x_7984 = v_3780 | ~v_1176;
assign x_7985 = v_3780 | ~v_1177;
assign x_7986 = v_3780 | ~v_3146;
assign x_7987 = v_3780 | ~v_3147;
assign x_7988 = v_3780 | ~v_1178;
assign x_7989 = v_3780 | ~v_3148;
assign x_7990 = v_3780 | ~v_3149;
assign x_7991 = v_3780 | ~v_1179;
assign x_7992 = v_3780 | ~v_3178;
assign x_7993 = v_3780 | ~v_3179;
assign x_7994 = v_3780 | ~v_804;
assign x_7995 = v_3780 | ~v_3180;
assign x_7996 = v_3780 | ~v_3181;
assign x_7997 = v_3780 | ~v_805;
assign x_7998 = v_3780 | ~v_3118;
assign x_7999 = v_3780 | ~v_3121;
assign x_8000 = v_3780 | ~v_1180;
assign x_8001 = v_3780 | ~v_1181;
assign x_8002 = v_3780 | ~v_183;
assign x_8003 = v_3780 | ~v_167;
assign x_8004 = v_3780 | ~v_165;
assign x_8005 = v_3780 | ~v_159;
assign x_8006 = v_3780 | ~v_146;
assign x_8007 = v_3780 | ~v_145;
assign x_8008 = v_3780 | ~v_144;
assign x_8009 = v_3780 | ~v_143;
assign x_8010 = v_3780 | ~v_142;
assign x_8011 = v_3780 | ~v_61;
assign x_8012 = v_3780 | ~v_58;
assign x_8013 = v_3780 | ~v_52;
assign x_8014 = v_3779 | ~v_1704;
assign x_8015 = v_3779 | ~v_1705;
assign x_8016 = v_3779 | ~v_1706;
assign x_8017 = v_3779 | ~v_1707;
assign x_8018 = v_3779 | ~v_1648;
assign x_8019 = v_3779 | ~v_1649;
assign x_8020 = v_3779 | ~v_1650;
assign x_8021 = v_3779 | ~v_1651;
assign x_8022 = v_3779 | ~v_3723;
assign x_8023 = v_3779 | ~v_3724;
assign x_8024 = v_3779 | ~v_1586;
assign x_8025 = v_3779 | ~v_3725;
assign x_8026 = v_3779 | ~v_3726;
assign x_8027 = v_3779 | ~v_1589;
assign x_8028 = v_3779 | ~v_1161;
assign x_8029 = v_3779 | ~v_1162;
assign x_8030 = v_3779 | ~v_3141;
assign x_8031 = v_3779 | ~v_3142;
assign x_8032 = v_3779 | ~v_1163;
assign x_8033 = v_3779 | ~v_3143;
assign x_8034 = v_3779 | ~v_3144;
assign x_8035 = v_3779 | ~v_1164;
assign x_8036 = v_3779 | ~v_3173;
assign x_8037 = v_3779 | ~v_3174;
assign x_8038 = v_3779 | ~v_771;
assign x_8039 = v_3779 | ~v_3175;
assign x_8040 = v_3779 | ~v_3176;
assign x_8041 = v_3779 | ~v_772;
assign x_8042 = v_3779 | ~v_1165;
assign x_8043 = v_3779 | ~v_1166;
assign x_8044 = v_3779 | ~v_182;
assign x_8045 = v_3779 | ~v_163;
assign x_8046 = v_3779 | ~v_161;
assign x_8047 = v_3779 | ~v_155;
assign x_8048 = v_3779 | ~v_138;
assign x_8049 = v_3779 | ~v_137;
assign x_8050 = v_3779 | ~v_136;
assign x_8051 = v_3779 | ~v_135;
assign x_8052 = v_3779 | ~v_134;
assign x_8053 = v_3779 | ~v_3107;
assign x_8054 = v_3779 | ~v_3108;
assign x_8055 = v_3779 | ~v_18;
assign x_8056 = v_3779 | ~v_15;
assign x_8057 = v_3779 | ~v_9;
assign x_8058 = ~v_3777 | ~v_3776 | ~v_3775 | v_3778;
assign x_8059 = v_3777 | ~v_1632;
assign x_8060 = v_3777 | ~v_1633;
assign x_8061 = v_3777 | ~v_1634;
assign x_8062 = v_3777 | ~v_1635;
assign x_8063 = v_3777 | ~v_3733;
assign x_8064 = v_3777 | ~v_3734;
assign x_8065 = v_3777 | ~v_1636;
assign x_8066 = v_3777 | ~v_1637;
assign x_8067 = v_3777 | ~v_1638;
assign x_8068 = v_3777 | ~v_3735;
assign x_8069 = v_3777 | ~v_3736;
assign x_8070 = v_3777 | ~v_1639;
assign x_8071 = v_3777 | ~v_1640;
assign x_8072 = v_3777 | ~v_1641;
assign x_8073 = v_3777 | ~v_1147;
assign x_8074 = v_3777 | ~v_1148;
assign x_8075 = v_3777 | ~v_3129;
assign x_8076 = v_3777 | ~v_3130;
assign x_8077 = v_3777 | ~v_975;
assign x_8078 = v_3777 | ~v_3131;
assign x_8079 = v_3777 | ~v_3132;
assign x_8080 = v_3777 | ~v_976;
assign x_8081 = v_3777 | ~v_3133;
assign x_8082 = v_3777 | ~v_3134;
assign x_8083 = v_3777 | ~v_3135;
assign x_8084 = v_3777 | ~v_839;
assign x_8085 = v_3777 | ~v_3136;
assign x_8086 = v_3777 | ~v_3137;
assign x_8087 = v_3777 | ~v_3138;
assign x_8088 = v_3777 | ~v_840;
assign x_8089 = v_3777 | ~v_1149;
assign x_8090 = v_3777 | ~v_1150;
assign x_8091 = v_3777 | ~v_184;
assign x_8092 = v_3777 | ~v_170;
assign x_8093 = v_3777 | ~v_150;
assign x_8094 = v_3777 | ~v_148;
assign x_8095 = v_3777 | ~v_147;
assign x_8096 = v_3777 | ~v_103;
assign x_8097 = v_3777 | ~v_102;
assign x_8098 = v_3777 | ~v_101;
assign x_8099 = v_3777 | ~v_100;
assign x_8100 = v_3777 | ~v_98;
assign x_8101 = v_3777 | ~v_97;
assign x_8102 = v_3777 | ~v_93;
assign x_8103 = v_3776 | ~v_1607;
assign x_8104 = v_3776 | ~v_1608;
assign x_8105 = v_3776 | ~v_1609;
assign x_8106 = v_3776 | ~v_1610;
assign x_8107 = v_3776 | ~v_3728;
assign x_8108 = v_3776 | ~v_3729;
assign x_8109 = v_3776 | ~v_1611;
assign x_8110 = v_3776 | ~v_1612;
assign x_8111 = v_3776 | ~v_1613;
assign x_8112 = v_3776 | ~v_3730;
assign x_8113 = v_3776 | ~v_3731;
assign x_8114 = v_3776 | ~v_1614;
assign x_8115 = v_3776 | ~v_1615;
assign x_8116 = v_3776 | ~v_1616;
assign x_8117 = v_3776 | ~v_1142;
assign x_8118 = v_3776 | ~v_1143;
assign x_8119 = v_3776 | ~v_3114;
assign x_8120 = v_3776 | ~v_3115;
assign x_8121 = v_3776 | ~v_960;
assign x_8122 = v_3776 | ~v_3116;
assign x_8123 = v_3776 | ~v_3117;
assign x_8124 = v_3776 | ~v_961;
assign x_8125 = v_3776 | ~v_3118;
assign x_8126 = v_3776 | ~v_3119;
assign x_8127 = v_3776 | ~v_3120;
assign x_8128 = v_3776 | ~v_806;
assign x_8129 = v_3776 | ~v_3121;
assign x_8130 = v_3776 | ~v_3122;
assign x_8131 = v_3776 | ~v_3123;
assign x_8132 = v_3776 | ~v_807;
assign x_8133 = v_3776 | ~v_1144;
assign x_8134 = v_3776 | ~v_1145;
assign x_8135 = v_3776 | ~v_183;
assign x_8136 = v_3776 | ~v_166;
assign x_8137 = v_3776 | ~v_145;
assign x_8138 = v_3776 | ~v_143;
assign x_8139 = v_3776 | ~v_142;
assign x_8140 = v_3776 | ~v_61;
assign x_8141 = v_3776 | ~v_60;
assign x_8142 = v_3776 | ~v_59;
assign x_8143 = v_3776 | ~v_58;
assign x_8144 = v_3776 | ~v_56;
assign x_8145 = v_3776 | ~v_55;
assign x_8146 = v_3776 | ~v_51;
assign x_8147 = v_3775 | ~v_1582;
assign x_8148 = v_3775 | ~v_1583;
assign x_8149 = v_3775 | ~v_1584;
assign x_8150 = v_3775 | ~v_1585;
assign x_8151 = v_3775 | ~v_3723;
assign x_8152 = v_3775 | ~v_3724;
assign x_8153 = v_3775 | ~v_1586;
assign x_8154 = v_3775 | ~v_1587;
assign x_8155 = v_3775 | ~v_1588;
assign x_8156 = v_3775 | ~v_3725;
assign x_8157 = v_3775 | ~v_3726;
assign x_8158 = v_3775 | ~v_1589;
assign x_8159 = v_3775 | ~v_1590;
assign x_8160 = v_3775 | ~v_1591;
assign x_8161 = v_3775 | ~v_1137;
assign x_8162 = v_3775 | ~v_1138;
assign x_8163 = v_3775 | ~v_3099;
assign x_8164 = v_3775 | ~v_3100;
assign x_8165 = v_3775 | ~v_945;
assign x_8166 = v_3775 | ~v_3101;
assign x_8167 = v_3775 | ~v_3102;
assign x_8168 = v_3775 | ~v_946;
assign x_8169 = v_3775 | ~v_3103;
assign x_8170 = v_3775 | ~v_3104;
assign x_8171 = v_3775 | ~v_773;
assign x_8172 = v_3775 | ~v_3105;
assign x_8173 = v_3775 | ~v_3106;
assign x_8174 = v_3775 | ~v_774;
assign x_8175 = v_3775 | ~v_1139;
assign x_8176 = v_3775 | ~v_1140;
assign x_8177 = v_3775 | ~v_182;
assign x_8178 = v_3775 | ~v_162;
assign x_8179 = v_3775 | ~v_137;
assign x_8180 = v_3775 | ~v_135;
assign x_8181 = v_3775 | ~v_134;
assign x_8182 = v_3775 | ~v_3107;
assign x_8183 = v_3775 | ~v_3108;
assign x_8184 = v_3775 | ~v_18;
assign x_8185 = v_3775 | ~v_17;
assign x_8186 = v_3775 | ~v_16;
assign x_8187 = v_3775 | ~v_15;
assign x_8188 = v_3775 | ~v_13;
assign x_8189 = v_3775 | ~v_12;
assign x_8190 = v_3775 | ~v_8;
assign x_8191 = ~v_3773 | ~v_3772 | ~v_3771 | v_3774;
assign x_8192 = v_3773 | ~v_1782;
assign x_8193 = v_3773 | ~v_1783;
assign x_8194 = v_3773 | ~v_1784;
assign x_8195 = v_3773 | ~v_1785;
assign x_8196 = v_3773 | ~v_3733;
assign x_8197 = v_3773 | ~v_3734;
assign x_8198 = v_3773 | ~v_1636;
assign x_8199 = v_3773 | ~v_1750;
assign x_8200 = v_3773 | ~v_1751;
assign x_8201 = v_3773 | ~v_3735;
assign x_8202 = v_3773 | ~v_3736;
assign x_8203 = v_3773 | ~v_1639;
assign x_8204 = v_3773 | ~v_1752;
assign x_8205 = v_3773 | ~v_1753;
assign x_8206 = v_3773 | ~v_3219;
assign x_8207 = v_3773 | ~v_3220;
assign x_8208 = v_3773 | ~v_1085;
assign x_8209 = v_3773 | ~v_1131;
assign x_8210 = v_3773 | ~v_1132;
assign x_8211 = v_3773 | ~v_3221;
assign x_8212 = v_3773 | ~v_3222;
assign x_8213 = v_3773 | ~v_1086;
assign x_8214 = v_3773 | ~v_1133;
assign x_8215 = v_3773 | ~v_1134;
assign x_8216 = v_3773 | ~v_3133;
assign x_8217 = v_3773 | ~v_3199;
assign x_8218 = v_3773 | ~v_3200;
assign x_8219 = v_3773 | ~v_1023;
assign x_8220 = v_3773 | ~v_3136;
assign x_8221 = v_3773 | ~v_3201;
assign x_8222 = v_3773 | ~v_3202;
assign x_8223 = v_3773 | ~v_1024;
assign x_8224 = v_3773 | ~v_184;
assign x_8225 = v_3773 | ~v_172;
assign x_8226 = v_3773 | ~v_171;
assign x_8227 = v_3773 | ~v_170;
assign x_8228 = v_3773 | ~v_169;
assign x_8229 = v_3773 | ~v_149;
assign x_8230 = v_3773 | ~v_147;
assign x_8231 = v_3773 | ~v_102;
assign x_8232 = v_3773 | ~v_101;
assign x_8233 = v_3773 | ~v_100;
assign x_8234 = v_3773 | ~v_99;
assign x_8235 = v_3773 | ~v_96;
assign x_8236 = v_3772 | ~v_1773;
assign x_8237 = v_3772 | ~v_1774;
assign x_8238 = v_3772 | ~v_1775;
assign x_8239 = v_3772 | ~v_1776;
assign x_8240 = v_3772 | ~v_3728;
assign x_8241 = v_3772 | ~v_3729;
assign x_8242 = v_3772 | ~v_1611;
assign x_8243 = v_3772 | ~v_1741;
assign x_8244 = v_3772 | ~v_1742;
assign x_8245 = v_3772 | ~v_3730;
assign x_8246 = v_3772 | ~v_3731;
assign x_8247 = v_3772 | ~v_1614;
assign x_8248 = v_3772 | ~v_1743;
assign x_8249 = v_3772 | ~v_1744;
assign x_8250 = v_3772 | ~v_3214;
assign x_8251 = v_3772 | ~v_3215;
assign x_8252 = v_3772 | ~v_1070;
assign x_8253 = v_3772 | ~v_1126;
assign x_8254 = v_3772 | ~v_1127;
assign x_8255 = v_3772 | ~v_3216;
assign x_8256 = v_3772 | ~v_3217;
assign x_8257 = v_3772 | ~v_1071;
assign x_8258 = v_3772 | ~v_1128;
assign x_8259 = v_3772 | ~v_1129;
assign x_8260 = v_3772 | ~v_3118;
assign x_8261 = v_3772 | ~v_3194;
assign x_8262 = v_3772 | ~v_3195;
assign x_8263 = v_3772 | ~v_1008;
assign x_8264 = v_3772 | ~v_3121;
assign x_8265 = v_3772 | ~v_1009;
assign x_8266 = v_3772 | ~v_3196;
assign x_8267 = v_3772 | ~v_183;
assign x_8268 = v_3772 | ~v_168;
assign x_8269 = v_3772 | ~v_167;
assign x_8270 = v_3772 | ~v_166;
assign x_8271 = v_3772 | ~v_165;
assign x_8272 = v_3772 | ~v_144;
assign x_8273 = v_3772 | ~v_142;
assign x_8274 = v_3772 | ~v_3197;
assign x_8275 = v_3772 | ~v_60;
assign x_8276 = v_3772 | ~v_59;
assign x_8277 = v_3772 | ~v_58;
assign x_8278 = v_3772 | ~v_57;
assign x_8279 = v_3772 | ~v_54;
assign x_8280 = v_3771 | ~v_1764;
assign x_8281 = v_3771 | ~v_1765;
assign x_8282 = v_3771 | ~v_1766;
assign x_8283 = v_3771 | ~v_1767;
assign x_8284 = v_3771 | ~v_3723;
assign x_8285 = v_3771 | ~v_3724;
assign x_8286 = v_3771 | ~v_1586;
assign x_8287 = v_3771 | ~v_1732;
assign x_8288 = v_3771 | ~v_1733;
assign x_8289 = v_3771 | ~v_3725;
assign x_8290 = v_3771 | ~v_3726;
assign x_8291 = v_3771 | ~v_1589;
assign x_8292 = v_3771 | ~v_1734;
assign x_8293 = v_3771 | ~v_1735;
assign x_8294 = v_3771 | ~v_3209;
assign x_8295 = v_3771 | ~v_3210;
assign x_8296 = v_3771 | ~v_1055;
assign x_8297 = v_3771 | ~v_1121;
assign x_8298 = v_3771 | ~v_1122;
assign x_8299 = v_3771 | ~v_3211;
assign x_8300 = v_3771 | ~v_3212;
assign x_8301 = v_3771 | ~v_1056;
assign x_8302 = v_3771 | ~v_1123;
assign x_8303 = v_3771 | ~v_1124;
assign x_8304 = v_3771 | ~v_3189;
assign x_8305 = v_3771 | ~v_3190;
assign x_8306 = v_3771 | ~v_3191;
assign x_8307 = v_3771 | ~v_3192;
assign x_8308 = v_3771 | ~v_182;
assign x_8309 = v_3771 | ~v_164;
assign x_8310 = v_3771 | ~v_163;
assign x_8311 = v_3771 | ~v_162;
assign x_8312 = v_3771 | ~v_161;
assign x_8313 = v_3771 | ~v_136;
assign x_8314 = v_3771 | ~v_134;
assign x_8315 = v_3771 | ~v_3107;
assign x_8316 = v_3771 | ~v_993;
assign x_8317 = v_3771 | ~v_3108;
assign x_8318 = v_3771 | ~v_994;
assign x_8319 = v_3771 | ~v_17;
assign x_8320 = v_3771 | ~v_16;
assign x_8321 = v_3771 | ~v_15;
assign x_8322 = v_3771 | ~v_14;
assign x_8323 = v_3771 | ~v_11;
assign x_8324 = ~v_3769 | ~v_3768 | ~v_3767 | v_3770;
assign x_8325 = v_3769 | ~v_1782;
assign x_8326 = v_3769 | ~v_1783;
assign x_8327 = v_3769 | ~v_1784;
assign x_8328 = v_3769 | ~v_1785;
assign x_8329 = v_3769 | ~v_1632;
assign x_8330 = v_3769 | ~v_1633;
assign x_8331 = v_3769 | ~v_1634;
assign x_8332 = v_3769 | ~v_1635;
assign x_8333 = v_3769 | ~v_3733;
assign x_8334 = v_3769 | ~v_3734;
assign x_8335 = v_3769 | ~v_1636;
assign x_8336 = v_3769 | ~v_3735;
assign x_8337 = v_3769 | ~v_3736;
assign x_8338 = v_3769 | ~v_1639;
assign x_8339 = v_3769 | ~v_3129;
assign x_8340 = v_3769 | ~v_3130;
assign x_8341 = v_3769 | ~v_975;
assign x_8342 = v_3769 | ~v_3131;
assign x_8343 = v_3769 | ~v_3132;
assign x_8344 = v_3769 | ~v_976;
assign x_8345 = v_3769 | ~v_1115;
assign x_8346 = v_3769 | ~v_1116;
assign x_8347 = v_3769 | ~v_3219;
assign x_8348 = v_3769 | ~v_3220;
assign x_8349 = v_3769 | ~v_1085;
assign x_8350 = v_3769 | ~v_3221;
assign x_8351 = v_3769 | ~v_3222;
assign x_8352 = v_3769 | ~v_1086;
assign x_8353 = v_3769 | ~v_3133;
assign x_8354 = v_3769 | ~v_3136;
assign x_8355 = v_3769 | ~v_1117;
assign x_8356 = v_3769 | ~v_1118;
assign x_8357 = v_3769 | ~v_184;
assign x_8358 = v_3769 | ~v_171;
assign x_8359 = v_3769 | ~v_170;
assign x_8360 = v_3769 | ~v_169;
assign x_8361 = v_3769 | ~v_151;
assign x_8362 = v_3769 | ~v_150;
assign x_8363 = v_3769 | ~v_148;
assign x_8364 = v_3769 | ~v_147;
assign x_8365 = v_3769 | ~v_103;
assign x_8366 = v_3769 | ~v_101;
assign x_8367 = v_3769 | ~v_100;
assign x_8368 = v_3769 | ~v_97;
assign x_8369 = v_3768 | ~v_1773;
assign x_8370 = v_3768 | ~v_1774;
assign x_8371 = v_3768 | ~v_1775;
assign x_8372 = v_3768 | ~v_1776;
assign x_8373 = v_3768 | ~v_1607;
assign x_8374 = v_3768 | ~v_1608;
assign x_8375 = v_3768 | ~v_1609;
assign x_8376 = v_3768 | ~v_1610;
assign x_8377 = v_3768 | ~v_3728;
assign x_8378 = v_3768 | ~v_3729;
assign x_8379 = v_3768 | ~v_1611;
assign x_8380 = v_3768 | ~v_3730;
assign x_8381 = v_3768 | ~v_3731;
assign x_8382 = v_3768 | ~v_1614;
assign x_8383 = v_3768 | ~v_3114;
assign x_8384 = v_3768 | ~v_3115;
assign x_8385 = v_3768 | ~v_960;
assign x_8386 = v_3768 | ~v_3116;
assign x_8387 = v_3768 | ~v_3117;
assign x_8388 = v_3768 | ~v_961;
assign x_8389 = v_3768 | ~v_1110;
assign x_8390 = v_3768 | ~v_1111;
assign x_8391 = v_3768 | ~v_3214;
assign x_8392 = v_3768 | ~v_3215;
assign x_8393 = v_3768 | ~v_1070;
assign x_8394 = v_3768 | ~v_3216;
assign x_8395 = v_3768 | ~v_3217;
assign x_8396 = v_3768 | ~v_1071;
assign x_8397 = v_3768 | ~v_3118;
assign x_8398 = v_3768 | ~v_3121;
assign x_8399 = v_3768 | ~v_1112;
assign x_8400 = v_3768 | ~v_1113;
assign x_8401 = v_3768 | ~v_183;
assign x_8402 = v_3768 | ~v_167;
assign x_8403 = v_3768 | ~v_166;
assign x_8404 = v_3768 | ~v_165;
assign x_8405 = v_3768 | ~v_146;
assign x_8406 = v_3768 | ~v_145;
assign x_8407 = v_3768 | ~v_143;
assign x_8408 = v_3768 | ~v_142;
assign x_8409 = v_3768 | ~v_61;
assign x_8410 = v_3768 | ~v_59;
assign x_8411 = v_3768 | ~v_58;
assign x_8412 = v_3768 | ~v_55;
assign x_8413 = v_3767 | ~v_1764;
assign x_8414 = v_3767 | ~v_1765;
assign x_8415 = v_3767 | ~v_1766;
assign x_8416 = v_3767 | ~v_1767;
assign x_8417 = v_3767 | ~v_1582;
assign x_8418 = v_3767 | ~v_1583;
assign x_8419 = v_3767 | ~v_1584;
assign x_8420 = v_3767 | ~v_1585;
assign x_8421 = v_3767 | ~v_3723;
assign x_8422 = v_3767 | ~v_3724;
assign x_8423 = v_3767 | ~v_1586;
assign x_8424 = v_3767 | ~v_3725;
assign x_8425 = v_3767 | ~v_3726;
assign x_8426 = v_3767 | ~v_1589;
assign x_8427 = v_3767 | ~v_3099;
assign x_8428 = v_3767 | ~v_3100;
assign x_8429 = v_3767 | ~v_945;
assign x_8430 = v_3767 | ~v_3101;
assign x_8431 = v_3767 | ~v_3102;
assign x_8432 = v_3767 | ~v_946;
assign x_8433 = v_3767 | ~v_1105;
assign x_8434 = v_3767 | ~v_1106;
assign x_8435 = v_3767 | ~v_3209;
assign x_8436 = v_3767 | ~v_3210;
assign x_8437 = v_3767 | ~v_1055;
assign x_8438 = v_3767 | ~v_3211;
assign x_8439 = v_3767 | ~v_3212;
assign x_8440 = v_3767 | ~v_1056;
assign x_8441 = v_3767 | ~v_1107;
assign x_8442 = v_3767 | ~v_1108;
assign x_8443 = v_3767 | ~v_182;
assign x_8444 = v_3767 | ~v_163;
assign x_8445 = v_3767 | ~v_162;
assign x_8446 = v_3767 | ~v_161;
assign x_8447 = v_3767 | ~v_138;
assign x_8448 = v_3767 | ~v_137;
assign x_8449 = v_3767 | ~v_135;
assign x_8450 = v_3767 | ~v_134;
assign x_8451 = v_3767 | ~v_3107;
assign x_8452 = v_3767 | ~v_3108;
assign x_8453 = v_3767 | ~v_18;
assign x_8454 = v_3767 | ~v_16;
assign x_8455 = v_3767 | ~v_15;
assign x_8456 = v_3767 | ~v_12;
assign x_8457 = ~v_3765 | ~v_3764 | ~v_3763 | v_3766;
assign x_8458 = v_3765 | ~v_1782;
assign x_8459 = v_3765 | ~v_1783;
assign x_8460 = v_3765 | ~v_1784;
assign x_8461 = v_3765 | ~v_1785;
assign x_8462 = v_3765 | ~v_1694;
assign x_8463 = v_3765 | ~v_1695;
assign x_8464 = v_3765 | ~v_1696;
assign x_8465 = v_3765 | ~v_1697;
assign x_8466 = v_3765 | ~v_3733;
assign x_8467 = v_3765 | ~v_3734;
assign x_8468 = v_3765 | ~v_1636;
assign x_8469 = v_3765 | ~v_3735;
assign x_8470 = v_3765 | ~v_3736;
assign x_8471 = v_3765 | ~v_1639;
assign x_8472 = v_3765 | ~v_3167;
assign x_8473 = v_3765 | ~v_3168;
assign x_8474 = v_3765 | ~v_927;
assign x_8475 = v_3765 | ~v_3169;
assign x_8476 = v_3765 | ~v_3170;
assign x_8477 = v_3765 | ~v_928;
assign x_8478 = v_3765 | ~v_1099;
assign x_8479 = v_3765 | ~v_1100;
assign x_8480 = v_3765 | ~v_1101;
assign x_8481 = v_3765 | ~v_1102;
assign x_8482 = v_3765 | ~v_3219;
assign x_8483 = v_3765 | ~v_3220;
assign x_8484 = v_3765 | ~v_1085;
assign x_8485 = v_3765 | ~v_3221;
assign x_8486 = v_3765 | ~v_3222;
assign x_8487 = v_3765 | ~v_1086;
assign x_8488 = v_3765 | ~v_3133;
assign x_8489 = v_3765 | ~v_3136;
assign x_8490 = v_3765 | ~v_184;
assign x_8491 = v_3765 | ~v_171;
assign x_8492 = v_3765 | ~v_170;
assign x_8493 = v_3765 | ~v_169;
assign x_8494 = v_3765 | ~v_150;
assign x_8495 = v_3765 | ~v_149;
assign x_8496 = v_3765 | ~v_148;
assign x_8497 = v_3765 | ~v_103;
assign x_8498 = v_3765 | ~v_102;
assign x_8499 = v_3765 | ~v_101;
assign x_8500 = v_3765 | ~v_100;
assign x_8501 = v_3765 | ~v_95;
assign x_8502 = v_3764 | ~v_1773;
assign x_8503 = v_3764 | ~v_1774;
assign x_8504 = v_3764 | ~v_1775;
assign x_8505 = v_3764 | ~v_1776;
assign x_8506 = v_3764 | ~v_1685;
assign x_8507 = v_3764 | ~v_1686;
assign x_8508 = v_3764 | ~v_1687;
assign x_8509 = v_3764 | ~v_1688;
assign x_8510 = v_3764 | ~v_3728;
assign x_8511 = v_3764 | ~v_3729;
assign x_8512 = v_3764 | ~v_1611;
assign x_8513 = v_3764 | ~v_3730;
assign x_8514 = v_3764 | ~v_3731;
assign x_8515 = v_3764 | ~v_1614;
assign x_8516 = v_3764 | ~v_3162;
assign x_8517 = v_3764 | ~v_3163;
assign x_8518 = v_3764 | ~v_912;
assign x_8519 = v_3764 | ~v_3164;
assign x_8520 = v_3764 | ~v_3165;
assign x_8521 = v_3764 | ~v_913;
assign x_8522 = v_3764 | ~v_1094;
assign x_8523 = v_3764 | ~v_1095;
assign x_8524 = v_3764 | ~v_1096;
assign x_8525 = v_3764 | ~v_1097;
assign x_8526 = v_3764 | ~v_3214;
assign x_8527 = v_3764 | ~v_3215;
assign x_8528 = v_3764 | ~v_1070;
assign x_8529 = v_3764 | ~v_3216;
assign x_8530 = v_3764 | ~v_3217;
assign x_8531 = v_3764 | ~v_1071;
assign x_8532 = v_3764 | ~v_3118;
assign x_8533 = v_3764 | ~v_3121;
assign x_8534 = v_3764 | ~v_183;
assign x_8535 = v_3764 | ~v_167;
assign x_8536 = v_3764 | ~v_166;
assign x_8537 = v_3764 | ~v_165;
assign x_8538 = v_3764 | ~v_145;
assign x_8539 = v_3764 | ~v_144;
assign x_8540 = v_3764 | ~v_143;
assign x_8541 = v_3764 | ~v_61;
assign x_8542 = v_3764 | ~v_60;
assign x_8543 = v_3764 | ~v_59;
assign x_8544 = v_3764 | ~v_58;
assign x_8545 = v_3764 | ~v_53;
assign x_8546 = v_3763 | ~v_1764;
assign x_8547 = v_3763 | ~v_1765;
assign x_8548 = v_3763 | ~v_1766;
assign x_8549 = v_3763 | ~v_1767;
assign x_8550 = v_3763 | ~v_1676;
assign x_8551 = v_3763 | ~v_1677;
assign x_8552 = v_3763 | ~v_1678;
assign x_8553 = v_3763 | ~v_1679;
assign x_8554 = v_3763 | ~v_3723;
assign x_8555 = v_3763 | ~v_3724;
assign x_8556 = v_3763 | ~v_1586;
assign x_8557 = v_3763 | ~v_3725;
assign x_8558 = v_3763 | ~v_3726;
assign x_8559 = v_3763 | ~v_1589;
assign x_8560 = v_3763 | ~v_3157;
assign x_8561 = v_3763 | ~v_3158;
assign x_8562 = v_3763 | ~v_897;
assign x_8563 = v_3763 | ~v_3159;
assign x_8564 = v_3763 | ~v_3160;
assign x_8565 = v_3763 | ~v_898;
assign x_8566 = v_3763 | ~v_1089;
assign x_8567 = v_3763 | ~v_1090;
assign x_8568 = v_3763 | ~v_1091;
assign x_8569 = v_3763 | ~v_1092;
assign x_8570 = v_3763 | ~v_3209;
assign x_8571 = v_3763 | ~v_3210;
assign x_8572 = v_3763 | ~v_1055;
assign x_8573 = v_3763 | ~v_3211;
assign x_8574 = v_3763 | ~v_3212;
assign x_8575 = v_3763 | ~v_1056;
assign x_8576 = v_3763 | ~v_182;
assign x_8577 = v_3763 | ~v_163;
assign x_8578 = v_3763 | ~v_162;
assign x_8579 = v_3763 | ~v_161;
assign x_8580 = v_3763 | ~v_137;
assign x_8581 = v_3763 | ~v_136;
assign x_8582 = v_3763 | ~v_135;
assign x_8583 = v_3763 | ~v_3107;
assign x_8584 = v_3763 | ~v_3108;
assign x_8585 = v_3763 | ~v_18;
assign x_8586 = v_3763 | ~v_17;
assign x_8587 = v_3763 | ~v_16;
assign x_8588 = v_3763 | ~v_15;
assign x_8589 = v_3763 | ~v_10;
assign x_8590 = ~v_3761 | ~v_3760 | ~v_3759 | v_3762;
assign x_8591 = v_3761 | ~v_1782;
assign x_8592 = v_3761 | ~v_1783;
assign x_8593 = v_3761 | ~v_1784;
assign x_8594 = v_3761 | ~v_1785;
assign x_8595 = v_3761 | ~v_1722;
assign x_8596 = v_3761 | ~v_1723;
assign x_8597 = v_3761 | ~v_1724;
assign x_8598 = v_3761 | ~v_1725;
assign x_8599 = v_3761 | ~v_3733;
assign x_8600 = v_3761 | ~v_3734;
assign x_8601 = v_3761 | ~v_1636;
assign x_8602 = v_3761 | ~v_3735;
assign x_8603 = v_3761 | ~v_3736;
assign x_8604 = v_3761 | ~v_1639;
assign x_8605 = v_3761 | ~v_3183;
assign x_8606 = v_3761 | ~v_3184;
assign x_8607 = v_3761 | ~v_837;
assign x_8608 = v_3761 | ~v_3185;
assign x_8609 = v_3761 | ~v_3186;
assign x_8610 = v_3761 | ~v_838;
assign x_8611 = v_3761 | ~v_1081;
assign x_8612 = v_3761 | ~v_1082;
assign x_8613 = v_3761 | ~v_1083;
assign x_8614 = v_3761 | ~v_1084;
assign x_8615 = v_3761 | ~v_3219;
assign x_8616 = v_3761 | ~v_3220;
assign x_8617 = v_3761 | ~v_1085;
assign x_8618 = v_3761 | ~v_3221;
assign x_8619 = v_3761 | ~v_3222;
assign x_8620 = v_3761 | ~v_1086;
assign x_8621 = v_3761 | ~v_3133;
assign x_8622 = v_3761 | ~v_3136;
assign x_8623 = v_3761 | ~v_184;
assign x_8624 = v_3761 | ~v_171;
assign x_8625 = v_3761 | ~v_170;
assign x_8626 = v_3761 | ~v_169;
assign x_8627 = v_3761 | ~v_160;
assign x_8628 = v_3761 | ~v_150;
assign x_8629 = v_3761 | ~v_149;
assign x_8630 = v_3761 | ~v_148;
assign x_8631 = v_3761 | ~v_147;
assign x_8632 = v_3761 | ~v_103;
assign x_8633 = v_3761 | ~v_102;
assign x_8634 = v_3761 | ~v_100;
assign x_8635 = v_3760 | ~v_1773;
assign x_8636 = v_3760 | ~v_1774;
assign x_8637 = v_3760 | ~v_1775;
assign x_8638 = v_3760 | ~v_1776;
assign x_8639 = v_3760 | ~v_1713;
assign x_8640 = v_3760 | ~v_1714;
assign x_8641 = v_3760 | ~v_1715;
assign x_8642 = v_3760 | ~v_1716;
assign x_8643 = v_3760 | ~v_3728;
assign x_8644 = v_3760 | ~v_3729;
assign x_8645 = v_3760 | ~v_1611;
assign x_8646 = v_3760 | ~v_3730;
assign x_8647 = v_3760 | ~v_3731;
assign x_8648 = v_3760 | ~v_1614;
assign x_8649 = v_3760 | ~v_3178;
assign x_8650 = v_3760 | ~v_3179;
assign x_8651 = v_3760 | ~v_804;
assign x_8652 = v_3760 | ~v_3180;
assign x_8653 = v_3760 | ~v_3181;
assign x_8654 = v_3760 | ~v_805;
assign x_8655 = v_3760 | ~v_1066;
assign x_8656 = v_3760 | ~v_1067;
assign x_8657 = v_3760 | ~v_1068;
assign x_8658 = v_3760 | ~v_1069;
assign x_8659 = v_3760 | ~v_3214;
assign x_8660 = v_3760 | ~v_3215;
assign x_8661 = v_3760 | ~v_1070;
assign x_8662 = v_3760 | ~v_3216;
assign x_8663 = v_3760 | ~v_3217;
assign x_8664 = v_3760 | ~v_1071;
assign x_8665 = v_3760 | ~v_3118;
assign x_8666 = v_3760 | ~v_3121;
assign x_8667 = v_3760 | ~v_183;
assign x_8668 = v_3760 | ~v_167;
assign x_8669 = v_3760 | ~v_166;
assign x_8670 = v_3760 | ~v_165;
assign x_8671 = v_3760 | ~v_159;
assign x_8672 = v_3760 | ~v_145;
assign x_8673 = v_3760 | ~v_144;
assign x_8674 = v_3760 | ~v_143;
assign x_8675 = v_3760 | ~v_142;
assign x_8676 = v_3760 | ~v_61;
assign x_8677 = v_3760 | ~v_60;
assign x_8678 = v_3760 | ~v_58;
assign x_8679 = v_3759 | ~v_1764;
assign x_8680 = v_3759 | ~v_1765;
assign x_8681 = v_3759 | ~v_1766;
assign x_8682 = v_3759 | ~v_1767;
assign x_8683 = v_3759 | ~v_1704;
assign x_8684 = v_3759 | ~v_1705;
assign x_8685 = v_3759 | ~v_1706;
assign x_8686 = v_3759 | ~v_1707;
assign x_8687 = v_3759 | ~v_3723;
assign x_8688 = v_3759 | ~v_3724;
assign x_8689 = v_3759 | ~v_1586;
assign x_8690 = v_3759 | ~v_3725;
assign x_8691 = v_3759 | ~v_3726;
assign x_8692 = v_3759 | ~v_1589;
assign x_8693 = v_3759 | ~v_3173;
assign x_8694 = v_3759 | ~v_3174;
assign x_8695 = v_3759 | ~v_771;
assign x_8696 = v_3759 | ~v_3175;
assign x_8697 = v_3759 | ~v_3176;
assign x_8698 = v_3759 | ~v_772;
assign x_8699 = v_3759 | ~v_1051;
assign x_8700 = v_3759 | ~v_1052;
assign x_8701 = v_3759 | ~v_1053;
assign x_8702 = v_3759 | ~v_1054;
assign x_8703 = v_3759 | ~v_3209;
assign x_8704 = v_3759 | ~v_3210;
assign x_8705 = v_3759 | ~v_1055;
assign x_8706 = v_3759 | ~v_3211;
assign x_8707 = v_3759 | ~v_3212;
assign x_8708 = v_3759 | ~v_1056;
assign x_8709 = v_3759 | ~v_182;
assign x_8710 = v_3759 | ~v_163;
assign x_8711 = v_3759 | ~v_162;
assign x_8712 = v_3759 | ~v_161;
assign x_8713 = v_3759 | ~v_155;
assign x_8714 = v_3759 | ~v_137;
assign x_8715 = v_3759 | ~v_136;
assign x_8716 = v_3759 | ~v_135;
assign x_8717 = v_3759 | ~v_134;
assign x_8718 = v_3759 | ~v_3107;
assign x_8719 = v_3759 | ~v_3108;
assign x_8720 = v_3759 | ~v_18;
assign x_8721 = v_3759 | ~v_17;
assign x_8722 = v_3759 | ~v_15;
assign x_8723 = ~v_3757 | ~v_3756 | ~v_3755 | v_3758;
assign x_8724 = v_3757 | ~v_1694;
assign x_8725 = v_3757 | ~v_1695;
assign x_8726 = v_3757 | ~v_1696;
assign x_8727 = v_3757 | ~v_1697;
assign x_8728 = v_3757 | ~v_3733;
assign x_8729 = v_3757 | ~v_3734;
assign x_8730 = v_3757 | ~v_1636;
assign x_8731 = v_3757 | ~v_1637;
assign x_8732 = v_3757 | ~v_1638;
assign x_8733 = v_3757 | ~v_3735;
assign x_8734 = v_3757 | ~v_3736;
assign x_8735 = v_3757 | ~v_1639;
assign x_8736 = v_3757 | ~v_1640;
assign x_8737 = v_3757 | ~v_1641;
assign x_8738 = v_3757 | ~v_1037;
assign x_8739 = v_3757 | ~v_1038;
assign x_8740 = v_3757 | ~v_1039;
assign x_8741 = v_3757 | ~v_1040;
assign x_8742 = v_3757 | ~v_3167;
assign x_8743 = v_3757 | ~v_3168;
assign x_8744 = v_3757 | ~v_927;
assign x_8745 = v_3757 | ~v_3169;
assign x_8746 = v_3757 | ~v_3170;
assign x_8747 = v_3757 | ~v_928;
assign x_8748 = v_3757 | ~v_3133;
assign x_8749 = v_3757 | ~v_3134;
assign x_8750 = v_3757 | ~v_3135;
assign x_8751 = v_3757 | ~v_839;
assign x_8752 = v_3757 | ~v_3136;
assign x_8753 = v_3757 | ~v_3137;
assign x_8754 = v_3757 | ~v_3138;
assign x_8755 = v_3757 | ~v_840;
assign x_8756 = v_3757 | ~v_184;
assign x_8757 = v_3757 | ~v_170;
assign x_8758 = v_3757 | ~v_151;
assign x_8759 = v_3757 | ~v_150;
assign x_8760 = v_3757 | ~v_149;
assign x_8761 = v_3757 | ~v_148;
assign x_8762 = v_3757 | ~v_147;
assign x_8763 = v_3757 | ~v_103;
assign x_8764 = v_3757 | ~v_101;
assign x_8765 = v_3757 | ~v_100;
assign x_8766 = v_3757 | ~v_98;
assign x_8767 = v_3757 | ~v_93;
assign x_8768 = v_3756 | ~v_1685;
assign x_8769 = v_3756 | ~v_1686;
assign x_8770 = v_3756 | ~v_1687;
assign x_8771 = v_3756 | ~v_1688;
assign x_8772 = v_3756 | ~v_3728;
assign x_8773 = v_3756 | ~v_3729;
assign x_8774 = v_3756 | ~v_1611;
assign x_8775 = v_3756 | ~v_1612;
assign x_8776 = v_3756 | ~v_1613;
assign x_8777 = v_3756 | ~v_3730;
assign x_8778 = v_3756 | ~v_3731;
assign x_8779 = v_3756 | ~v_1614;
assign x_8780 = v_3756 | ~v_1615;
assign x_8781 = v_3756 | ~v_1616;
assign x_8782 = v_3756 | ~v_1032;
assign x_8783 = v_3756 | ~v_1033;
assign x_8784 = v_3756 | ~v_1034;
assign x_8785 = v_3756 | ~v_1035;
assign x_8786 = v_3756 | ~v_3162;
assign x_8787 = v_3756 | ~v_3163;
assign x_8788 = v_3756 | ~v_912;
assign x_8789 = v_3756 | ~v_3164;
assign x_8790 = v_3756 | ~v_3165;
assign x_8791 = v_3756 | ~v_913;
assign x_8792 = v_3756 | ~v_3118;
assign x_8793 = v_3756 | ~v_3119;
assign x_8794 = v_3756 | ~v_3120;
assign x_8795 = v_3756 | ~v_806;
assign x_8796 = v_3756 | ~v_3121;
assign x_8797 = v_3756 | ~v_3122;
assign x_8798 = v_3756 | ~v_3123;
assign x_8799 = v_3756 | ~v_807;
assign x_8800 = v_3756 | ~v_183;
assign x_8801 = v_3756 | ~v_166;
assign x_8802 = v_3756 | ~v_146;
assign x_8803 = v_3756 | ~v_145;
assign x_8804 = v_3756 | ~v_144;
assign x_8805 = v_3756 | ~v_143;
assign x_8806 = v_3756 | ~v_142;
assign x_8807 = v_3756 | ~v_61;
assign x_8808 = v_3756 | ~v_59;
assign x_8809 = v_3756 | ~v_58;
assign x_8810 = v_3756 | ~v_56;
assign x_8811 = v_3756 | ~v_51;
assign x_8812 = v_3755 | ~v_1676;
assign x_8813 = v_3755 | ~v_1677;
assign x_8814 = v_3755 | ~v_1678;
assign x_8815 = v_3755 | ~v_1679;
assign x_8816 = v_3755 | ~v_3723;
assign x_8817 = v_3755 | ~v_3724;
assign x_8818 = v_3755 | ~v_1586;
assign x_8819 = v_3755 | ~v_1587;
assign x_8820 = v_3755 | ~v_1588;
assign x_8821 = v_3755 | ~v_3725;
assign x_8822 = v_3755 | ~v_3726;
assign x_8823 = v_3755 | ~v_1589;
assign x_8824 = v_3755 | ~v_1590;
assign x_8825 = v_3755 | ~v_1591;
assign x_8826 = v_3755 | ~v_1027;
assign x_8827 = v_3755 | ~v_1028;
assign x_8828 = v_3755 | ~v_1029;
assign x_8829 = v_3755 | ~v_1030;
assign x_8830 = v_3755 | ~v_3157;
assign x_8831 = v_3755 | ~v_3158;
assign x_8832 = v_3755 | ~v_897;
assign x_8833 = v_3755 | ~v_3159;
assign x_8834 = v_3755 | ~v_3160;
assign x_8835 = v_3755 | ~v_898;
assign x_8836 = v_3755 | ~v_3103;
assign x_8837 = v_3755 | ~v_3104;
assign x_8838 = v_3755 | ~v_773;
assign x_8839 = v_3755 | ~v_3105;
assign x_8840 = v_3755 | ~v_3106;
assign x_8841 = v_3755 | ~v_774;
assign x_8842 = v_3755 | ~v_182;
assign x_8843 = v_3755 | ~v_162;
assign x_8844 = v_3755 | ~v_138;
assign x_8845 = v_3755 | ~v_137;
assign x_8846 = v_3755 | ~v_136;
assign x_8847 = v_3755 | ~v_135;
assign x_8848 = v_3755 | ~v_134;
assign x_8849 = v_3755 | ~v_3107;
assign x_8850 = v_3755 | ~v_3108;
assign x_8851 = v_3755 | ~v_18;
assign x_8852 = v_3755 | ~v_16;
assign x_8853 = v_3755 | ~v_15;
assign x_8854 = v_3755 | ~v_13;
assign x_8855 = v_3755 | ~v_8;
assign x_8856 = ~v_3753 | ~v_3752 | ~v_3751 | v_3754;
assign x_8857 = v_3753 | ~v_1826;
assign x_8858 = v_3753 | ~v_1827;
assign x_8859 = v_3753 | ~v_1828;
assign x_8860 = v_3753 | ~v_1829;
assign x_8861 = v_3753 | ~v_3733;
assign x_8862 = v_3753 | ~v_3734;
assign x_8863 = v_3753 | ~v_1636;
assign x_8864 = v_3753 | ~v_1750;
assign x_8865 = v_3753 | ~v_1751;
assign x_8866 = v_3753 | ~v_3735;
assign x_8867 = v_3753 | ~v_3736;
assign x_8868 = v_3753 | ~v_1639;
assign x_8869 = v_3753 | ~v_1752;
assign x_8870 = v_3753 | ~v_1753;
assign x_8871 = v_3753 | ~v_3251;
assign x_8872 = v_3753 | ~v_3252;
assign x_8873 = v_3753 | ~v_885;
assign x_8874 = v_3753 | ~v_1019;
assign x_8875 = v_3753 | ~v_1020;
assign x_8876 = v_3753 | ~v_3253;
assign x_8877 = v_3753 | ~v_3254;
assign x_8878 = v_3753 | ~v_886;
assign x_8879 = v_3753 | ~v_1021;
assign x_8880 = v_3753 | ~v_1022;
assign x_8881 = v_3753 | ~v_3133;
assign x_8882 = v_3753 | ~v_3199;
assign x_8883 = v_3753 | ~v_3200;
assign x_8884 = v_3753 | ~v_1023;
assign x_8885 = v_3753 | ~v_3136;
assign x_8886 = v_3753 | ~v_3201;
assign x_8887 = v_3753 | ~v_3202;
assign x_8888 = v_3753 | ~v_1024;
assign x_8889 = v_3753 | ~v_184;
assign x_8890 = v_3753 | ~v_181;
assign x_8891 = v_3753 | ~v_171;
assign x_8892 = v_3753 | ~v_170;
assign x_8893 = v_3753 | ~v_169;
assign x_8894 = v_3753 | ~v_149;
assign x_8895 = v_3753 | ~v_147;
assign x_8896 = v_3753 | ~v_103;
assign x_8897 = v_3753 | ~v_102;
assign x_8898 = v_3753 | ~v_101;
assign x_8899 = v_3753 | ~v_99;
assign x_8900 = v_3753 | ~v_96;
assign x_8901 = v_3752 | ~v_1817;
assign x_8902 = v_3752 | ~v_1818;
assign x_8903 = v_3752 | ~v_1819;
assign x_8904 = v_3752 | ~v_1820;
assign x_8905 = v_3752 | ~v_3728;
assign x_8906 = v_3752 | ~v_3729;
assign x_8907 = v_3752 | ~v_1611;
assign x_8908 = v_3752 | ~v_1741;
assign x_8909 = v_3752 | ~v_1742;
assign x_8910 = v_3752 | ~v_3730;
assign x_8911 = v_3752 | ~v_3731;
assign x_8912 = v_3752 | ~v_1614;
assign x_8913 = v_3752 | ~v_1743;
assign x_8914 = v_3752 | ~v_1744;
assign x_8915 = v_3752 | ~v_3246;
assign x_8916 = v_3752 | ~v_3247;
assign x_8917 = v_3752 | ~v_870;
assign x_8918 = v_3752 | ~v_1004;
assign x_8919 = v_3752 | ~v_1005;
assign x_8920 = v_3752 | ~v_3248;
assign x_8921 = v_3752 | ~v_3249;
assign x_8922 = v_3752 | ~v_871;
assign x_8923 = v_3752 | ~v_1006;
assign x_8924 = v_3752 | ~v_1007;
assign x_8925 = v_3752 | ~v_3118;
assign x_8926 = v_3752 | ~v_3194;
assign x_8927 = v_3752 | ~v_3195;
assign x_8928 = v_3752 | ~v_1008;
assign x_8929 = v_3752 | ~v_3121;
assign x_8930 = v_3752 | ~v_1009;
assign x_8931 = v_3752 | ~v_3196;
assign x_8932 = v_3752 | ~v_183;
assign x_8933 = v_3752 | ~v_180;
assign x_8934 = v_3752 | ~v_167;
assign x_8935 = v_3752 | ~v_166;
assign x_8936 = v_3752 | ~v_165;
assign x_8937 = v_3752 | ~v_144;
assign x_8938 = v_3752 | ~v_142;
assign x_8939 = v_3752 | ~v_3197;
assign x_8940 = v_3752 | ~v_61;
assign x_8941 = v_3752 | ~v_60;
assign x_8942 = v_3752 | ~v_59;
assign x_8943 = v_3752 | ~v_57;
assign x_8944 = v_3752 | ~v_54;
assign x_8945 = v_3751 | ~v_1808;
assign x_8946 = v_3751 | ~v_1809;
assign x_8947 = v_3751 | ~v_1810;
assign x_8948 = v_3751 | ~v_1811;
assign x_8949 = v_3751 | ~v_3723;
assign x_8950 = v_3751 | ~v_3724;
assign x_8951 = v_3751 | ~v_1586;
assign x_8952 = v_3751 | ~v_1732;
assign x_8953 = v_3751 | ~v_1733;
assign x_8954 = v_3751 | ~v_3725;
assign x_8955 = v_3751 | ~v_3726;
assign x_8956 = v_3751 | ~v_1589;
assign x_8957 = v_3751 | ~v_1734;
assign x_8958 = v_3751 | ~v_1735;
assign x_8959 = v_3751 | ~v_3241;
assign x_8960 = v_3751 | ~v_3242;
assign x_8961 = v_3751 | ~v_855;
assign x_8962 = v_3751 | ~v_989;
assign x_8963 = v_3751 | ~v_990;
assign x_8964 = v_3751 | ~v_3243;
assign x_8965 = v_3751 | ~v_3244;
assign x_8966 = v_3751 | ~v_856;
assign x_8967 = v_3751 | ~v_991;
assign x_8968 = v_3751 | ~v_992;
assign x_8969 = v_3751 | ~v_3189;
assign x_8970 = v_3751 | ~v_3190;
assign x_8971 = v_3751 | ~v_3191;
assign x_8972 = v_3751 | ~v_3192;
assign x_8973 = v_3751 | ~v_182;
assign x_8974 = v_3751 | ~v_179;
assign x_8975 = v_3751 | ~v_163;
assign x_8976 = v_3751 | ~v_162;
assign x_8977 = v_3751 | ~v_161;
assign x_8978 = v_3751 | ~v_136;
assign x_8979 = v_3751 | ~v_134;
assign x_8980 = v_3751 | ~v_3107;
assign x_8981 = v_3751 | ~v_993;
assign x_8982 = v_3751 | ~v_3108;
assign x_8983 = v_3751 | ~v_994;
assign x_8984 = v_3751 | ~v_18;
assign x_8985 = v_3751 | ~v_17;
assign x_8986 = v_3751 | ~v_16;
assign x_8987 = v_3751 | ~v_14;
assign x_8988 = v_3751 | ~v_11;
assign x_8989 = ~v_3749 | ~v_3748 | ~v_3747 | v_3750;
assign x_8990 = v_3749 | ~v_1826;
assign x_8991 = v_3749 | ~v_1827;
assign x_8992 = v_3749 | ~v_1828;
assign x_8993 = v_3749 | ~v_1829;
assign x_8994 = v_3749 | ~v_1632;
assign x_8995 = v_3749 | ~v_1633;
assign x_8996 = v_3749 | ~v_1634;
assign x_8997 = v_3749 | ~v_1635;
assign x_8998 = v_3749 | ~v_3733;
assign x_8999 = v_3749 | ~v_3734;
assign x_9000 = v_3749 | ~v_1636;
assign x_9001 = v_3749 | ~v_3735;
assign x_9002 = v_3749 | ~v_3736;
assign x_9003 = v_3749 | ~v_1639;
assign x_9004 = v_3749 | ~v_973;
assign x_9005 = v_3749 | ~v_974;
assign x_9006 = v_3749 | ~v_3251;
assign x_9007 = v_3749 | ~v_3252;
assign x_9008 = v_3749 | ~v_885;
assign x_9009 = v_3749 | ~v_3253;
assign x_9010 = v_3749 | ~v_3254;
assign x_9011 = v_3749 | ~v_886;
assign x_9012 = v_3749 | ~v_3129;
assign x_9013 = v_3749 | ~v_3130;
assign x_9014 = v_3749 | ~v_975;
assign x_9015 = v_3749 | ~v_3131;
assign x_9016 = v_3749 | ~v_3132;
assign x_9017 = v_3749 | ~v_976;
assign x_9018 = v_3749 | ~v_3133;
assign x_9019 = v_3749 | ~v_3136;
assign x_9020 = v_3749 | ~v_977;
assign x_9021 = v_3749 | ~v_978;
assign x_9022 = v_3749 | ~v_184;
assign x_9023 = v_3749 | ~v_181;
assign x_9024 = v_3749 | ~v_172;
assign x_9025 = v_3749 | ~v_171;
assign x_9026 = v_3749 | ~v_170;
assign x_9027 = v_3749 | ~v_169;
assign x_9028 = v_3749 | ~v_150;
assign x_9029 = v_3749 | ~v_148;
assign x_9030 = v_3749 | ~v_147;
assign x_9031 = v_3749 | ~v_102;
assign x_9032 = v_3749 | ~v_101;
assign x_9033 = v_3749 | ~v_97;
assign x_9034 = v_3748 | ~v_1817;
assign x_9035 = v_3748 | ~v_1818;
assign x_9036 = v_3748 | ~v_1819;
assign x_9037 = v_3748 | ~v_1820;
assign x_9038 = v_3748 | ~v_1607;
assign x_9039 = v_3748 | ~v_1608;
assign x_9040 = v_3748 | ~v_1609;
assign x_9041 = v_3748 | ~v_1610;
assign x_9042 = v_3748 | ~v_3728;
assign x_9043 = v_3748 | ~v_3729;
assign x_9044 = v_3748 | ~v_1611;
assign x_9045 = v_3748 | ~v_3730;
assign x_9046 = v_3748 | ~v_3731;
assign x_9047 = v_3748 | ~v_1614;
assign x_9048 = v_3748 | ~v_958;
assign x_9049 = v_3748 | ~v_959;
assign x_9050 = v_3748 | ~v_3246;
assign x_9051 = v_3748 | ~v_3247;
assign x_9052 = v_3748 | ~v_870;
assign x_9053 = v_3748 | ~v_3248;
assign x_9054 = v_3748 | ~v_3249;
assign x_9055 = v_3748 | ~v_871;
assign x_9056 = v_3748 | ~v_3114;
assign x_9057 = v_3748 | ~v_3115;
assign x_9058 = v_3748 | ~v_960;
assign x_9059 = v_3748 | ~v_3116;
assign x_9060 = v_3748 | ~v_3117;
assign x_9061 = v_3748 | ~v_961;
assign x_9062 = v_3748 | ~v_3118;
assign x_9063 = v_3748 | ~v_3121;
assign x_9064 = v_3748 | ~v_962;
assign x_9065 = v_3748 | ~v_963;
assign x_9066 = v_3748 | ~v_183;
assign x_9067 = v_3748 | ~v_180;
assign x_9068 = v_3748 | ~v_168;
assign x_9069 = v_3748 | ~v_167;
assign x_9070 = v_3748 | ~v_166;
assign x_9071 = v_3748 | ~v_165;
assign x_9072 = v_3748 | ~v_145;
assign x_9073 = v_3748 | ~v_143;
assign x_9074 = v_3748 | ~v_142;
assign x_9075 = v_3748 | ~v_60;
assign x_9076 = v_3748 | ~v_59;
assign x_9077 = v_3748 | ~v_55;
assign x_9078 = v_3747 | ~v_1808;
assign x_9079 = v_3747 | ~v_1809;
assign x_9080 = v_3747 | ~v_1810;
assign x_9081 = v_3747 | ~v_1811;
assign x_9082 = v_3747 | ~v_1582;
assign x_9083 = v_3747 | ~v_1583;
assign x_9084 = v_3747 | ~v_1584;
assign x_9085 = v_3747 | ~v_1585;
assign x_9086 = v_3747 | ~v_3723;
assign x_9087 = v_3747 | ~v_3724;
assign x_9088 = v_3747 | ~v_1586;
assign x_9089 = v_3747 | ~v_3725;
assign x_9090 = v_3747 | ~v_3726;
assign x_9091 = v_3747 | ~v_1589;
assign x_9092 = v_3747 | ~v_943;
assign x_9093 = v_3747 | ~v_944;
assign x_9094 = v_3747 | ~v_3241;
assign x_9095 = v_3747 | ~v_3242;
assign x_9096 = v_3747 | ~v_855;
assign x_9097 = v_3747 | ~v_3243;
assign x_9098 = v_3747 | ~v_3244;
assign x_9099 = v_3747 | ~v_856;
assign x_9100 = v_3747 | ~v_3099;
assign x_9101 = v_3747 | ~v_3100;
assign x_9102 = v_3747 | ~v_945;
assign x_9103 = v_3747 | ~v_3101;
assign x_9104 = v_3747 | ~v_3102;
assign x_9105 = v_3747 | ~v_946;
assign x_9106 = v_3747 | ~v_947;
assign x_9107 = v_3747 | ~v_948;
assign x_9108 = v_3747 | ~v_182;
assign x_9109 = v_3747 | ~v_179;
assign x_9110 = v_3747 | ~v_164;
assign x_9111 = v_3747 | ~v_163;
assign x_9112 = v_3747 | ~v_162;
assign x_9113 = v_3747 | ~v_161;
assign x_9114 = v_3747 | ~v_137;
assign x_9115 = v_3747 | ~v_135;
assign x_9116 = v_3747 | ~v_134;
assign x_9117 = v_3747 | ~v_3107;
assign x_9118 = v_3747 | ~v_3108;
assign x_9119 = v_3747 | ~v_17;
assign x_9120 = v_3747 | ~v_16;
assign x_9121 = v_3747 | ~v_12;
assign x_9122 = ~v_3745 | ~v_3744 | ~v_3743 | v_3746;
assign x_9123 = v_3745 | ~v_1826;
assign x_9124 = v_3745 | ~v_1827;
assign x_9125 = v_3745 | ~v_1828;
assign x_9126 = v_3745 | ~v_1829;
assign x_9127 = v_3745 | ~v_1694;
assign x_9128 = v_3745 | ~v_1695;
assign x_9129 = v_3745 | ~v_1696;
assign x_9130 = v_3745 | ~v_1697;
assign x_9131 = v_3745 | ~v_3733;
assign x_9132 = v_3745 | ~v_3734;
assign x_9133 = v_3745 | ~v_1636;
assign x_9134 = v_3745 | ~v_3735;
assign x_9135 = v_3745 | ~v_3736;
assign x_9136 = v_3745 | ~v_1639;
assign x_9137 = v_3745 | ~v_925;
assign x_9138 = v_3745 | ~v_926;
assign x_9139 = v_3745 | ~v_3251;
assign x_9140 = v_3745 | ~v_3252;
assign x_9141 = v_3745 | ~v_885;
assign x_9142 = v_3745 | ~v_3253;
assign x_9143 = v_3745 | ~v_3254;
assign x_9144 = v_3745 | ~v_886;
assign x_9145 = v_3745 | ~v_3167;
assign x_9146 = v_3745 | ~v_3168;
assign x_9147 = v_3745 | ~v_927;
assign x_9148 = v_3745 | ~v_3169;
assign x_9149 = v_3745 | ~v_3170;
assign x_9150 = v_3745 | ~v_928;
assign x_9151 = v_3745 | ~v_3133;
assign x_9152 = v_3745 | ~v_3136;
assign x_9153 = v_3745 | ~v_929;
assign x_9154 = v_3745 | ~v_930;
assign x_9155 = v_3745 | ~v_184;
assign x_9156 = v_3745 | ~v_181;
assign x_9157 = v_3745 | ~v_171;
assign x_9158 = v_3745 | ~v_170;
assign x_9159 = v_3745 | ~v_169;
assign x_9160 = v_3745 | ~v_150;
assign x_9161 = v_3745 | ~v_149;
assign x_9162 = v_3745 | ~v_148;
assign x_9163 = v_3745 | ~v_147;
assign x_9164 = v_3745 | ~v_103;
assign x_9165 = v_3745 | ~v_102;
assign x_9166 = v_3745 | ~v_101;
assign x_9167 = v_3744 | ~v_1817;
assign x_9168 = v_3744 | ~v_1818;
assign x_9169 = v_3744 | ~v_1819;
assign x_9170 = v_3744 | ~v_1820;
assign x_9171 = v_3744 | ~v_1685;
assign x_9172 = v_3744 | ~v_1686;
assign x_9173 = v_3744 | ~v_1687;
assign x_9174 = v_3744 | ~v_1688;
assign x_9175 = v_3744 | ~v_3728;
assign x_9176 = v_3744 | ~v_3729;
assign x_9177 = v_3744 | ~v_1611;
assign x_9178 = v_3744 | ~v_3730;
assign x_9179 = v_3744 | ~v_3731;
assign x_9180 = v_3744 | ~v_1614;
assign x_9181 = v_3744 | ~v_910;
assign x_9182 = v_3744 | ~v_911;
assign x_9183 = v_3744 | ~v_3246;
assign x_9184 = v_3744 | ~v_3247;
assign x_9185 = v_3744 | ~v_870;
assign x_9186 = v_3744 | ~v_3248;
assign x_9187 = v_3744 | ~v_3249;
assign x_9188 = v_3744 | ~v_871;
assign x_9189 = v_3744 | ~v_3162;
assign x_9190 = v_3744 | ~v_3163;
assign x_9191 = v_3744 | ~v_912;
assign x_9192 = v_3744 | ~v_3164;
assign x_9193 = v_3744 | ~v_3165;
assign x_9194 = v_3744 | ~v_913;
assign x_9195 = v_3744 | ~v_3118;
assign x_9196 = v_3744 | ~v_3121;
assign x_9197 = v_3744 | ~v_914;
assign x_9198 = v_3744 | ~v_915;
assign x_9199 = v_3744 | ~v_183;
assign x_9200 = v_3744 | ~v_180;
assign x_9201 = v_3744 | ~v_167;
assign x_9202 = v_3744 | ~v_166;
assign x_9203 = v_3744 | ~v_165;
assign x_9204 = v_3744 | ~v_145;
assign x_9205 = v_3744 | ~v_144;
assign x_9206 = v_3744 | ~v_143;
assign x_9207 = v_3744 | ~v_142;
assign x_9208 = v_3744 | ~v_61;
assign x_9209 = v_3744 | ~v_60;
assign x_9210 = v_3744 | ~v_59;
assign x_9211 = v_3743 | ~v_1808;
assign x_9212 = v_3743 | ~v_1809;
assign x_9213 = v_3743 | ~v_1810;
assign x_9214 = v_3743 | ~v_1811;
assign x_9215 = v_3743 | ~v_1676;
assign x_9216 = v_3743 | ~v_1677;
assign x_9217 = v_3743 | ~v_1678;
assign x_9218 = v_3743 | ~v_1679;
assign x_9219 = v_3743 | ~v_3723;
assign x_9220 = v_3743 | ~v_3724;
assign x_9221 = v_3743 | ~v_1586;
assign x_9222 = v_3743 | ~v_3725;
assign x_9223 = v_3743 | ~v_3726;
assign x_9224 = v_3743 | ~v_1589;
assign x_9225 = v_3743 | ~v_895;
assign x_9226 = v_3743 | ~v_896;
assign x_9227 = v_3743 | ~v_3241;
assign x_9228 = v_3743 | ~v_3242;
assign x_9229 = v_3743 | ~v_855;
assign x_9230 = v_3743 | ~v_3243;
assign x_9231 = v_3743 | ~v_3244;
assign x_9232 = v_3743 | ~v_856;
assign x_9233 = v_3743 | ~v_3157;
assign x_9234 = v_3743 | ~v_3158;
assign x_9235 = v_3743 | ~v_897;
assign x_9236 = v_3743 | ~v_3159;
assign x_9237 = v_3743 | ~v_3160;
assign x_9238 = v_3743 | ~v_898;
assign x_9239 = v_3743 | ~v_899;
assign x_9240 = v_3743 | ~v_900;
assign x_9241 = v_3743 | ~v_182;
assign x_9242 = v_3743 | ~v_179;
assign x_9243 = v_3743 | ~v_163;
assign x_9244 = v_3743 | ~v_162;
assign x_9245 = v_3743 | ~v_161;
assign x_9246 = v_3743 | ~v_137;
assign x_9247 = v_3743 | ~v_136;
assign x_9248 = v_3743 | ~v_135;
assign x_9249 = v_3743 | ~v_134;
assign x_9250 = v_3743 | ~v_3107;
assign x_9251 = v_3743 | ~v_3108;
assign x_9252 = v_3743 | ~v_18;
assign x_9253 = v_3743 | ~v_17;
assign x_9254 = v_3743 | ~v_16;
assign x_9255 = ~v_3741 | ~v_3740 | ~v_3739 | v_3742;
assign x_9256 = v_3741 | ~v_1826;
assign x_9257 = v_3741 | ~v_1827;
assign x_9258 = v_3741 | ~v_1828;
assign x_9259 = v_3741 | ~v_1829;
assign x_9260 = v_3741 | ~v_1722;
assign x_9261 = v_3741 | ~v_1723;
assign x_9262 = v_3741 | ~v_1724;
assign x_9263 = v_3741 | ~v_1725;
assign x_9264 = v_3741 | ~v_3733;
assign x_9265 = v_3741 | ~v_3734;
assign x_9266 = v_3741 | ~v_1636;
assign x_9267 = v_3741 | ~v_3735;
assign x_9268 = v_3741 | ~v_3736;
assign x_9269 = v_3741 | ~v_1639;
assign x_9270 = v_3741 | ~v_881;
assign x_9271 = v_3741 | ~v_882;
assign x_9272 = v_3741 | ~v_883;
assign x_9273 = v_3741 | ~v_884;
assign x_9274 = v_3741 | ~v_3251;
assign x_9275 = v_3741 | ~v_3252;
assign x_9276 = v_3741 | ~v_885;
assign x_9277 = v_3741 | ~v_3253;
assign x_9278 = v_3741 | ~v_3254;
assign x_9279 = v_3741 | ~v_886;
assign x_9280 = v_3741 | ~v_3183;
assign x_9281 = v_3741 | ~v_3184;
assign x_9282 = v_3741 | ~v_837;
assign x_9283 = v_3741 | ~v_3185;
assign x_9284 = v_3741 | ~v_3186;
assign x_9285 = v_3741 | ~v_838;
assign x_9286 = v_3741 | ~v_3133;
assign x_9287 = v_3741 | ~v_3136;
assign x_9288 = v_3741 | ~v_184;
assign x_9289 = v_3741 | ~v_181;
assign x_9290 = v_3741 | ~v_171;
assign x_9291 = v_3741 | ~v_170;
assign x_9292 = v_3741 | ~v_169;
assign x_9293 = v_3741 | ~v_160;
assign x_9294 = v_3741 | ~v_150;
assign x_9295 = v_3741 | ~v_149;
assign x_9296 = v_3741 | ~v_148;
assign x_9297 = v_3741 | ~v_103;
assign x_9298 = v_3741 | ~v_102;
assign x_9299 = v_3741 | ~v_95;
assign x_9300 = v_3740 | ~v_1817;
assign x_9301 = v_3740 | ~v_1818;
assign x_9302 = v_3740 | ~v_1819;
assign x_9303 = v_3740 | ~v_1820;
assign x_9304 = v_3740 | ~v_1713;
assign x_9305 = v_3740 | ~v_1714;
assign x_9306 = v_3740 | ~v_1715;
assign x_9307 = v_3740 | ~v_1716;
assign x_9308 = v_3740 | ~v_3728;
assign x_9309 = v_3740 | ~v_3729;
assign x_9310 = v_3740 | ~v_1611;
assign x_9311 = v_3740 | ~v_3730;
assign x_9312 = v_3740 | ~v_3731;
assign x_9313 = v_3740 | ~v_1614;
assign x_9314 = v_3740 | ~v_866;
assign x_9315 = v_3740 | ~v_867;
assign x_9316 = v_3740 | ~v_868;
assign x_9317 = v_3740 | ~v_869;
assign x_9318 = v_3740 | ~v_3246;
assign x_9319 = v_3740 | ~v_3247;
assign x_9320 = v_3740 | ~v_870;
assign x_9321 = v_3740 | ~v_3248;
assign x_9322 = v_3740 | ~v_3249;
assign x_9323 = v_3740 | ~v_871;
assign x_9324 = v_3740 | ~v_3178;
assign x_9325 = v_3740 | ~v_3179;
assign x_9326 = v_3740 | ~v_804;
assign x_9327 = v_3740 | ~v_3180;
assign x_9328 = v_3740 | ~v_3181;
assign x_9329 = v_3740 | ~v_805;
assign x_9330 = v_3740 | ~v_3118;
assign x_9331 = v_3740 | ~v_3121;
assign x_9332 = v_3740 | ~v_183;
assign x_9333 = v_3740 | ~v_180;
assign x_9334 = v_3740 | ~v_167;
assign x_9335 = v_3740 | ~v_166;
assign x_9336 = v_3740 | ~v_165;
assign x_9337 = v_3740 | ~v_159;
assign x_9338 = v_3740 | ~v_145;
assign x_9339 = v_3740 | ~v_144;
assign x_9340 = v_3740 | ~v_143;
assign x_9341 = v_3740 | ~v_61;
assign x_9342 = v_3740 | ~v_60;
assign x_9343 = v_3740 | ~v_53;
assign x_9344 = v_3739 | ~v_1808;
assign x_9345 = v_3739 | ~v_1809;
assign x_9346 = v_3739 | ~v_1810;
assign x_9347 = v_3739 | ~v_1811;
assign x_9348 = v_3739 | ~v_1704;
assign x_9349 = v_3739 | ~v_1705;
assign x_9350 = v_3739 | ~v_1706;
assign x_9351 = v_3739 | ~v_1707;
assign x_9352 = v_3739 | ~v_3723;
assign x_9353 = v_3739 | ~v_3724;
assign x_9354 = v_3739 | ~v_1586;
assign x_9355 = v_3739 | ~v_3725;
assign x_9356 = v_3739 | ~v_3726;
assign x_9357 = v_3739 | ~v_1589;
assign x_9358 = v_3739 | ~v_851;
assign x_9359 = v_3739 | ~v_852;
assign x_9360 = v_3739 | ~v_853;
assign x_9361 = v_3739 | ~v_854;
assign x_9362 = v_3739 | ~v_3241;
assign x_9363 = v_3739 | ~v_3242;
assign x_9364 = v_3739 | ~v_855;
assign x_9365 = v_3739 | ~v_3243;
assign x_9366 = v_3739 | ~v_3244;
assign x_9367 = v_3739 | ~v_856;
assign x_9368 = v_3739 | ~v_3173;
assign x_9369 = v_3739 | ~v_3174;
assign x_9370 = v_3739 | ~v_771;
assign x_9371 = v_3739 | ~v_3175;
assign x_9372 = v_3739 | ~v_3176;
assign x_9373 = v_3739 | ~v_772;
assign x_9374 = v_3739 | ~v_182;
assign x_9375 = v_3739 | ~v_179;
assign x_9376 = v_3739 | ~v_163;
assign x_9377 = v_3739 | ~v_162;
assign x_9378 = v_3739 | ~v_161;
assign x_9379 = v_3739 | ~v_155;
assign x_9380 = v_3739 | ~v_137;
assign x_9381 = v_3739 | ~v_136;
assign x_9382 = v_3739 | ~v_135;
assign x_9383 = v_3739 | ~v_3107;
assign x_9384 = v_3739 | ~v_3108;
assign x_9385 = v_3739 | ~v_18;
assign x_9386 = v_3739 | ~v_17;
assign x_9387 = v_3739 | ~v_10;
assign x_9388 = ~v_3737 | ~v_3732 | ~v_3727 | v_3738;
assign x_9389 = v_3737 | ~v_1722;
assign x_9390 = v_3737 | ~v_1723;
assign x_9391 = v_3737 | ~v_1724;
assign x_9392 = v_3737 | ~v_1725;
assign x_9393 = v_3737 | ~v_3733;
assign x_9394 = v_3737 | ~v_3734;
assign x_9395 = v_3737 | ~v_1636;
assign x_9396 = v_3737 | ~v_1637;
assign x_9397 = v_3737 | ~v_1638;
assign x_9398 = v_3737 | ~v_3735;
assign x_9399 = v_3737 | ~v_3736;
assign x_9400 = v_3737 | ~v_1639;
assign x_9401 = v_3737 | ~v_1640;
assign x_9402 = v_3737 | ~v_1641;
assign x_9403 = v_3737 | ~v_833;
assign x_9404 = v_3737 | ~v_834;
assign x_9405 = v_3737 | ~v_835;
assign x_9406 = v_3737 | ~v_836;
assign x_9407 = v_3737 | ~v_3183;
assign x_9408 = v_3737 | ~v_3184;
assign x_9409 = v_3737 | ~v_837;
assign x_9410 = v_3737 | ~v_3185;
assign x_9411 = v_3737 | ~v_3186;
assign x_9412 = v_3737 | ~v_838;
assign x_9413 = v_3737 | ~v_3133;
assign x_9414 = v_3737 | ~v_3134;
assign x_9415 = v_3737 | ~v_3135;
assign x_9416 = v_3737 | ~v_839;
assign x_9417 = v_3737 | ~v_3136;
assign x_9418 = v_3737 | ~v_3137;
assign x_9419 = v_3737 | ~v_3138;
assign x_9420 = v_3737 | ~v_840;
assign x_9421 = v_3737 | ~v_184;
assign x_9422 = v_3737 | ~v_170;
assign x_9423 = v_3737 | ~v_160;
assign x_9424 = v_3737 | ~v_150;
assign x_9425 = v_3737 | ~v_149;
assign x_9426 = v_3737 | ~v_148;
assign x_9427 = v_3737 | ~v_147;
assign x_9428 = v_3737 | ~v_103;
assign x_9429 = v_3737 | ~v_102;
assign x_9430 = v_3737 | ~v_100;
assign x_9431 = v_3737 | ~v_98;
assign x_9432 = v_3737 | ~v_93;
assign x_9433 = ~v_123 | ~v_153 | v_3736;
assign x_9434 = ~v_120 | ~v_152 | v_3735;
assign x_9435 = ~v_108 | v_153 | v_3734;
assign x_9436 = ~v_105 | v_152 | v_3733;
assign x_9437 = v_3732 | ~v_1713;
assign x_9438 = v_3732 | ~v_1714;
assign x_9439 = v_3732 | ~v_1715;
assign x_9440 = v_3732 | ~v_1716;
assign x_9441 = v_3732 | ~v_3728;
assign x_9442 = v_3732 | ~v_3729;
assign x_9443 = v_3732 | ~v_1611;
assign x_9444 = v_3732 | ~v_1612;
assign x_9445 = v_3732 | ~v_1613;
assign x_9446 = v_3732 | ~v_3730;
assign x_9447 = v_3732 | ~v_3731;
assign x_9448 = v_3732 | ~v_1614;
assign x_9449 = v_3732 | ~v_1615;
assign x_9450 = v_3732 | ~v_1616;
assign x_9451 = v_3732 | ~v_800;
assign x_9452 = v_3732 | ~v_801;
assign x_9453 = v_3732 | ~v_802;
assign x_9454 = v_3732 | ~v_803;
assign x_9455 = v_3732 | ~v_3178;
assign x_9456 = v_3732 | ~v_3179;
assign x_9457 = v_3732 | ~v_804;
assign x_9458 = v_3732 | ~v_3180;
assign x_9459 = v_3732 | ~v_3181;
assign x_9460 = v_3732 | ~v_805;
assign x_9461 = v_3732 | ~v_3118;
assign x_9462 = v_3732 | ~v_3119;
assign x_9463 = v_3732 | ~v_3120;
assign x_9464 = v_3732 | ~v_806;
assign x_9465 = v_3732 | ~v_3121;
assign x_9466 = v_3732 | ~v_3122;
assign x_9467 = v_3732 | ~v_3123;
assign x_9468 = v_3732 | ~v_807;
assign x_9469 = v_3732 | ~v_183;
assign x_9470 = v_3732 | ~v_166;
assign x_9471 = v_3732 | ~v_159;
assign x_9472 = v_3732 | ~v_145;
assign x_9473 = v_3732 | ~v_144;
assign x_9474 = v_3732 | ~v_143;
assign x_9475 = v_3732 | ~v_142;
assign x_9476 = v_3732 | ~v_61;
assign x_9477 = v_3732 | ~v_60;
assign x_9478 = v_3732 | ~v_58;
assign x_9479 = v_3732 | ~v_56;
assign x_9480 = v_3732 | ~v_51;
assign x_9481 = ~v_81 | ~v_153 | v_3731;
assign x_9482 = ~v_78 | ~v_152 | v_3730;
assign x_9483 = ~v_66 | v_153 | v_3729;
assign x_9484 = ~v_63 | v_152 | v_3728;
assign x_9485 = v_3727 | ~v_1704;
assign x_9486 = v_3727 | ~v_1705;
assign x_9487 = v_3727 | ~v_1706;
assign x_9488 = v_3727 | ~v_1707;
assign x_9489 = v_3727 | ~v_3723;
assign x_9490 = v_3727 | ~v_3724;
assign x_9491 = v_3727 | ~v_1586;
assign x_9492 = v_3727 | ~v_1587;
assign x_9493 = v_3727 | ~v_1588;
assign x_9494 = v_3727 | ~v_3725;
assign x_9495 = v_3727 | ~v_3726;
assign x_9496 = v_3727 | ~v_1589;
assign x_9497 = v_3727 | ~v_1590;
assign x_9498 = v_3727 | ~v_1591;
assign x_9499 = v_3727 | ~v_767;
assign x_9500 = v_3727 | ~v_768;
assign x_9501 = v_3727 | ~v_769;
assign x_9502 = v_3727 | ~v_770;
assign x_9503 = v_3727 | ~v_3173;
assign x_9504 = v_3727 | ~v_3174;
assign x_9505 = v_3727 | ~v_771;
assign x_9506 = v_3727 | ~v_3175;
assign x_9507 = v_3727 | ~v_3176;
assign x_9508 = v_3727 | ~v_772;
assign x_9509 = v_3727 | ~v_3103;
assign x_9510 = v_3727 | ~v_3104;
assign x_9511 = v_3727 | ~v_773;
assign x_9512 = v_3727 | ~v_3105;
assign x_9513 = v_3727 | ~v_3106;
assign x_9514 = v_3727 | ~v_774;
assign x_9515 = v_3727 | ~v_182;
assign x_9516 = v_3727 | ~v_162;
assign x_9517 = v_3727 | ~v_155;
assign x_9518 = v_3727 | ~v_137;
assign x_9519 = v_3727 | ~v_136;
assign x_9520 = v_3727 | ~v_135;
assign x_9521 = v_3727 | ~v_134;
assign x_9522 = v_3727 | ~v_3107;
assign x_9523 = v_3727 | ~v_3108;
assign x_9524 = v_3727 | ~v_18;
assign x_9525 = v_3727 | ~v_17;
assign x_9526 = v_3727 | ~v_15;
assign x_9527 = v_3727 | ~v_13;
assign x_9528 = v_3727 | ~v_8;
assign x_9529 = ~v_39 | ~v_153 | v_3726;
assign x_9530 = ~v_36 | ~v_152 | v_3725;
assign x_9531 = ~v_24 | v_153 | v_3724;
assign x_9532 = ~v_21 | v_152 | v_3723;
assign x_9533 = v_3722 | ~v_1562;
assign x_9534 = v_3722 | ~v_728;
assign x_9535 = v_3721 | ~v_2034;
assign x_9536 = v_3721 | ~v_727;
assign x_9537 = ~v_725 | ~v_724 | ~v_723 | ~v_722 | ~v_3719 | ~v_3715 | ~v_3711 | ~v_3707 | ~v_3703 | ~v_3699 | ~v_3695 | ~v_3691 | ~v_3687 | ~v_3683 | ~v_3679 | ~v_3675 | ~v_3671 | ~v_3667 | ~v_3663 | ~v_3659 | ~v_3643 | v_3720;
assign x_9538 = v_3719 | ~v_3716;
assign x_9539 = v_3719 | ~v_3717;
assign x_9540 = v_3719 | ~v_3718;
assign x_9541 = v_98 | v_103 | v_101 | v_96 | v_100 | v_95 | v_99 | v_93 | v_102 | ~v_719 | ~v_718 | v_170 | v_149 | v_184 | ~v_483 | ~v_717 | ~v_3021 | ~v_299 | ~v_2957 | ~v_3020 | ~v_2956 | ~v_2955 | ~v_482 | ~v_716 | ~v_3019 | ~v_298 | ~v_2954 | ~v_3018 | ~v_2953 | ~v_2952 | ~v_1464 | ~v_1352 | ~v_1463 | ~v_1351 | ~v_1350 | ~v_3657 | ~v_3656 | ~v_1462 | ~v_1349 | ~v_1461 | ~v_1348 | ~v_1347 | ~v_3655 | ~v_3654 | v_3718;
assign x_9542 = v_54 | v_53 | v_56 | v_61 | v_51 | v_60 | v_59 | v_58 | v_57 | ~v_714 | ~v_713 | ~v_3016 | v_144 | v_166 | v_183 | ~v_3015 | ~v_266 | ~v_2942 | ~v_468 | ~v_712 | ~v_2941 | ~v_2940 | ~v_467 | ~v_711 | ~v_3014 | ~v_265 | ~v_2939 | ~v_3013 | ~v_2938 | ~v_2937 | ~v_1455 | ~v_1327 | ~v_1454 | ~v_1326 | ~v_1325 | ~v_3652 | ~v_3651 | ~v_1453 | ~v_1324 | ~v_1452 | ~v_1323 | ~v_1322 | ~v_3650 | ~v_3649 | v_3717;
assign x_9543 = v_13 | v_18 | v_17 | v_16 | v_8 | v_15 | v_14 | v_11 | v_10 | ~v_453 | ~v_709 | ~v_2927 | ~v_452 | ~v_708 | ~v_2926 | v_136 | ~v_707 | ~v_706 | v_162 | v_182 | ~v_3011 | ~v_233 | ~v_2925 | ~v_3010 | ~v_2924 | ~v_3009 | ~v_232 | ~v_2923 | ~v_3008 | ~v_2922 | ~v_1446 | ~v_1302 | ~v_1445 | ~v_1301 | ~v_1300 | ~v_3647 | ~v_3646 | ~v_1444 | ~v_1299 | ~v_1443 | ~v_1298 | ~v_1297 | ~v_3645 | ~v_3644 | v_3716;
assign x_9544 = v_3715 | ~v_3712;
assign x_9545 = v_3715 | ~v_3713;
assign x_9546 = v_3715 | ~v_3714;
assign x_9547 = v_103 | v_101 | v_96 | v_100 | v_94 | v_99 | v_102 | v_171 | v_169 | v_149 | v_147 | v_184 | ~v_703 | ~v_702 | ~v_483 | ~v_3021 | ~v_3020 | ~v_2955 | ~v_482 | ~v_3019 | ~v_3018 | ~v_2952 | ~v_701 | ~v_653 | ~v_2973 | ~v_2972 | ~v_700 | ~v_652 | ~v_2971 | ~v_2970 | ~v_1464 | ~v_1463 | ~v_1350 | ~v_3657 | ~v_3656 | ~v_1462 | ~v_1461 | ~v_1347 | ~v_3655 | ~v_3654 | ~v_1380 | ~v_1379 | ~v_1378 | ~v_1377 | v_3714;
assign x_9548 = v_54 | v_61 | v_52 | v_60 | v_59 | v_58 | v_57 | ~v_3016 | v_144 | v_142 | v_167 | v_165 | v_183 | ~v_698 | ~v_697 | ~v_3015 | ~v_468 | ~v_2940 | ~v_467 | ~v_3014 | ~v_3013 | ~v_2937 | ~v_696 | ~v_638 | ~v_2968 | ~v_2967 | ~v_695 | ~v_637 | ~v_2966 | ~v_2965 | ~v_1455 | ~v_1454 | ~v_1325 | ~v_3652 | ~v_3651 | ~v_1453 | ~v_1452 | ~v_1322 | ~v_3650 | ~v_3649 | ~v_1371 | ~v_1370 | ~v_1369 | ~v_1368 | v_3713;
assign x_9549 = v_9 | v_18 | v_17 | v_16 | v_15 | v_14 | v_11 | ~v_453 | ~v_2927 | ~v_452 | ~v_2926 | v_136 | v_134 | v_163 | v_161 | v_182 | ~v_693 | ~v_692 | ~v_3011 | ~v_3010 | ~v_3009 | ~v_3008 | ~v_691 | ~v_623 | ~v_2963 | ~v_2962 | ~v_690 | ~v_622 | ~v_2961 | ~v_2960 | ~v_1446 | ~v_1445 | ~v_1300 | ~v_3647 | ~v_3646 | ~v_1444 | ~v_1443 | ~v_1297 | ~v_3645 | ~v_3644 | ~v_1362 | ~v_1361 | ~v_1360 | ~v_1359 | v_3712;
assign x_9550 = v_3711 | ~v_3708;
assign x_9551 = v_3711 | ~v_3709;
assign x_9552 = v_3711 | ~v_3710;
assign x_9553 = v_103 | v_101 | v_97 | v_100 | v_95 | v_94 | v_102 | v_171 | v_169 | v_150 | v_148 | v_184 | ~v_2955 | ~v_2952 | ~v_435 | ~v_2951 | ~v_2950 | ~v_434 | ~v_2949 | ~v_2948 | ~v_653 | ~v_2973 | ~v_2972 | ~v_652 | ~v_2971 | ~v_2970 | ~v_687 | ~v_686 | ~v_685 | ~v_684 | ~v_1350 | ~v_3657 | ~v_3656 | ~v_1347 | ~v_3655 | ~v_3654 | ~v_1380 | ~v_1379 | ~v_1378 | ~v_1377 | ~v_1346 | ~v_1345 | ~v_1344 | ~v_1343 | v_3710;
assign x_9554 = v_53 | v_55 | v_61 | v_52 | v_60 | v_59 | v_58 | v_145 | v_143 | v_167 | v_165 | v_183 | ~v_2940 | ~v_2937 | ~v_420 | ~v_2936 | ~v_2935 | ~v_419 | ~v_2934 | ~v_2933 | ~v_638 | ~v_2968 | ~v_2967 | ~v_637 | ~v_2966 | ~v_2965 | ~v_682 | ~v_681 | ~v_680 | ~v_679 | ~v_1325 | ~v_3652 | ~v_3651 | ~v_1322 | ~v_3650 | ~v_3649 | ~v_1371 | ~v_1370 | ~v_1369 | ~v_1368 | ~v_1321 | ~v_1320 | ~v_1319 | ~v_1318 | v_3709;
assign x_9555 = v_9 | v_18 | v_17 | v_16 | v_15 | v_12 | v_10 | ~v_2927 | ~v_2926 | v_135 | v_137 | v_163 | v_161 | v_182 | ~v_405 | ~v_2921 | ~v_2920 | ~v_404 | ~v_2919 | ~v_2918 | ~v_623 | ~v_2963 | ~v_2962 | ~v_622 | ~v_2961 | ~v_2960 | ~v_677 | ~v_676 | ~v_675 | ~v_674 | ~v_1300 | ~v_3647 | ~v_3646 | ~v_1297 | ~v_3645 | ~v_3644 | ~v_1362 | ~v_1361 | ~v_1360 | ~v_1359 | ~v_1296 | ~v_1295 | ~v_1294 | ~v_1293 | v_3708;
assign x_9556 = v_3707 | ~v_3704;
assign x_9557 = v_3707 | ~v_3705;
assign x_9558 = v_3707 | ~v_3706;
assign x_9559 = v_101 | v_100 | v_94 | v_102 | v_172 | v_171 | v_169 | v_150 | v_149 | v_148 | v_147 | v_184 | ~v_671 | ~v_670 | ~v_2955 | ~v_2952 | ~v_387 | ~v_2989 | ~v_2988 | ~v_386 | ~v_2987 | ~v_2986 | ~v_653 | ~v_2973 | ~v_2972 | ~v_652 | ~v_2971 | ~v_2970 | ~v_669 | ~v_668 | ~v_1350 | ~v_3657 | ~v_3656 | ~v_1347 | ~v_3655 | ~v_3654 | ~v_1380 | ~v_1379 | ~v_1378 | ~v_1377 | ~v_1408 | ~v_1407 | ~v_1406 | ~v_1405 | v_3706;
assign x_9560 = v_52 | v_60 | v_59 | v_58 | v_144 | v_145 | v_143 | v_142 | v_168 | v_167 | v_165 | v_183 | ~v_666 | ~v_665 | ~v_2940 | ~v_2937 | ~v_372 | ~v_2984 | ~v_2983 | ~v_371 | ~v_2982 | ~v_2981 | ~v_638 | ~v_2968 | ~v_2967 | ~v_637 | ~v_2966 | ~v_2965 | ~v_664 | ~v_663 | ~v_1325 | ~v_3652 | ~v_3651 | ~v_1322 | ~v_3650 | ~v_3649 | ~v_1371 | ~v_1370 | ~v_1369 | ~v_1368 | ~v_1399 | ~v_1398 | ~v_1397 | ~v_1396 | v_3705;
assign x_9561 = v_9 | v_17 | v_16 | v_15 | ~v_2927 | ~v_2926 | v_136 | v_135 | v_134 | v_137 | v_164 | v_163 | v_161 | v_182 | ~v_661 | ~v_660 | ~v_357 | ~v_2979 | ~v_2978 | ~v_356 | ~v_2977 | ~v_2976 | ~v_623 | ~v_2963 | ~v_2962 | ~v_622 | ~v_2961 | ~v_2960 | ~v_659 | ~v_658 | ~v_1300 | ~v_3647 | ~v_3646 | ~v_1297 | ~v_3645 | ~v_3644 | ~v_1362 | ~v_1361 | ~v_1360 | ~v_1359 | ~v_1390 | ~v_1389 | ~v_1388 | ~v_1387 | v_3704;
assign x_9562 = v_3703 | ~v_3700;
assign x_9563 = v_3703 | ~v_3701;
assign x_9564 = v_3703 | ~v_3702;
assign x_9565 = v_103 | v_100 | v_94 | v_151 | v_171 | v_169 | v_160 | v_150 | v_149 | v_148 | v_147 | v_184 | ~v_655 | ~v_654 | ~v_2955 | ~v_2952 | ~v_297 | ~v_3005 | ~v_3004 | ~v_296 | ~v_3003 | ~v_3002 | ~v_653 | ~v_2973 | ~v_2972 | ~v_652 | ~v_2971 | ~v_2970 | ~v_651 | ~v_650 | ~v_1350 | ~v_3657 | ~v_3656 | ~v_1347 | ~v_3655 | ~v_3654 | ~v_1380 | ~v_1379 | ~v_1378 | ~v_1377 | ~v_1436 | ~v_1435 | ~v_1434 | ~v_1433 | v_3702;
assign x_9566 = v_61 | v_52 | v_58 | v_144 | v_159 | v_145 | v_143 | v_142 | v_167 | v_165 | v_146 | v_183 | ~v_640 | ~v_639 | ~v_2940 | ~v_2937 | ~v_264 | ~v_3000 | ~v_2999 | ~v_263 | ~v_2998 | ~v_2997 | ~v_638 | ~v_2968 | ~v_2967 | ~v_637 | ~v_2966 | ~v_2965 | ~v_636 | ~v_635 | ~v_1325 | ~v_3652 | ~v_3651 | ~v_1322 | ~v_3650 | ~v_3649 | ~v_1371 | ~v_1370 | ~v_1369 | ~v_1368 | ~v_1427 | ~v_1426 | ~v_1425 | ~v_1424 | v_3701;
assign x_9567 = v_9 | v_18 | v_15 | ~v_2927 | ~v_2926 | v_136 | v_135 | v_134 | v_137 | v_138 | v_163 | v_161 | v_155 | v_182 | ~v_625 | ~v_624 | ~v_231 | ~v_2995 | ~v_2994 | ~v_230 | ~v_2993 | ~v_2992 | ~v_623 | ~v_2963 | ~v_2962 | ~v_622 | ~v_2961 | ~v_2960 | ~v_621 | ~v_620 | ~v_1300 | ~v_3647 | ~v_3646 | ~v_1297 | ~v_3645 | ~v_3644 | ~v_1362 | ~v_1361 | ~v_1360 | ~v_1359 | ~v_1418 | ~v_1417 | ~v_1416 | ~v_1415 | v_3700;
assign x_9568 = v_3699 | ~v_3696;
assign x_9569 = v_3699 | ~v_3697;
assign x_9570 = v_3699 | ~v_3698;
assign x_9571 = v_98 | v_103 | v_101 | v_97 | v_100 | v_93 | v_102 | v_170 | v_150 | v_148 | v_147 | v_184 | ~v_609 | ~v_608 | ~v_299 | ~v_2957 | ~v_2956 | ~v_2955 | ~v_298 | ~v_2954 | ~v_2953 | ~v_2952 | ~v_435 | ~v_2951 | ~v_2950 | ~v_434 | ~v_2949 | ~v_2948 | ~v_607 | ~v_606 | ~v_1352 | ~v_1351 | ~v_1350 | ~v_3657 | ~v_3656 | ~v_1349 | ~v_1348 | ~v_1347 | ~v_3655 | ~v_3654 | ~v_1346 | ~v_1345 | ~v_1344 | ~v_1343 | v_3698;
assign x_9572 = v_56 | v_55 | v_61 | v_51 | v_60 | v_59 | v_58 | v_145 | v_143 | v_142 | v_166 | v_183 | ~v_604 | ~v_603 | ~v_266 | ~v_2942 | ~v_2941 | ~v_2940 | ~v_265 | ~v_2939 | ~v_2938 | ~v_2937 | ~v_420 | ~v_2936 | ~v_2935 | ~v_419 | ~v_2934 | ~v_2933 | ~v_602 | ~v_601 | ~v_1327 | ~v_1326 | ~v_1325 | ~v_3652 | ~v_3651 | ~v_1324 | ~v_1323 | ~v_1322 | ~v_3650 | ~v_3649 | ~v_1321 | ~v_1320 | ~v_1319 | ~v_1318 | v_3697;
assign x_9573 = v_13 | v_18 | v_17 | v_16 | v_8 | v_15 | v_12 | ~v_2927 | ~v_2926 | v_135 | v_134 | v_137 | v_162 | v_182 | ~v_599 | ~v_598 | ~v_233 | ~v_2925 | ~v_2924 | ~v_232 | ~v_2923 | ~v_2922 | ~v_405 | ~v_2921 | ~v_2920 | ~v_404 | ~v_2919 | ~v_2918 | ~v_597 | ~v_596 | ~v_1302 | ~v_1301 | ~v_1300 | ~v_3647 | ~v_3646 | ~v_1299 | ~v_1298 | ~v_1297 | ~v_3645 | ~v_3644 | ~v_1296 | ~v_1295 | ~v_1294 | ~v_1293 | v_3696;
assign x_9574 = v_3695 | ~v_3692;
assign x_9575 = v_3695 | ~v_3693;
assign x_9576 = v_3695 | ~v_3694;
assign x_9577 = v_101 | v_96 | v_100 | v_99 | v_102 | v_172 | v_171 | v_170 | v_169 | v_149 | v_147 | v_184 | ~v_483 | ~v_3021 | ~v_3020 | ~v_2955 | ~v_482 | ~v_3019 | ~v_3018 | ~v_2952 | ~v_593 | ~v_592 | ~v_545 | ~v_3041 | ~v_3040 | ~v_591 | ~v_590 | ~v_544 | ~v_3039 | ~v_3038 | ~v_1464 | ~v_1463 | ~v_1350 | ~v_3657 | ~v_3656 | ~v_1462 | ~v_1461 | ~v_1347 | ~v_3655 | ~v_3654 | ~v_1496 | ~v_1495 | ~v_1494 | ~v_1493 | v_3694;
assign x_9578 = v_54 | v_60 | v_59 | v_58 | v_57 | ~v_3016 | v_144 | v_142 | v_168 | v_167 | v_166 | v_165 | v_183 | ~v_3015 | ~v_468 | ~v_2940 | ~v_467 | ~v_3014 | ~v_3013 | ~v_2937 | ~v_588 | ~v_587 | ~v_530 | ~v_3036 | ~v_3035 | ~v_586 | ~v_585 | ~v_529 | ~v_3034 | ~v_3033 | ~v_1455 | ~v_1454 | ~v_1325 | ~v_3652 | ~v_3651 | ~v_1453 | ~v_1452 | ~v_1322 | ~v_3650 | ~v_3649 | ~v_1487 | ~v_1486 | ~v_1485 | ~v_1484 | v_3693;
assign x_9579 = v_17 | v_16 | v_15 | v_14 | v_11 | ~v_453 | ~v_2927 | ~v_452 | ~v_2926 | v_136 | v_134 | v_164 | v_163 | v_162 | v_161 | v_182 | ~v_3011 | ~v_3010 | ~v_3009 | ~v_3008 | ~v_583 | ~v_582 | ~v_515 | ~v_3031 | ~v_3030 | ~v_581 | ~v_580 | ~v_514 | ~v_3029 | ~v_3028 | ~v_1446 | ~v_1445 | ~v_1300 | ~v_3647 | ~v_3646 | ~v_1444 | ~v_1443 | ~v_1297 | ~v_3645 | ~v_3644 | ~v_1478 | ~v_1477 | ~v_1476 | ~v_1475 | v_3692;
assign x_9580 = v_3691 | ~v_3688;
assign x_9581 = v_3691 | ~v_3689;
assign x_9582 = v_3691 | ~v_3690;
assign x_9583 = v_103 | v_101 | v_97 | v_100 | v_151 | v_171 | v_170 | v_169 | v_150 | v_148 | v_147 | v_184 | ~v_577 | ~v_576 | ~v_2955 | ~v_2952 | ~v_545 | ~v_3041 | ~v_3040 | ~v_544 | ~v_3039 | ~v_3038 | ~v_575 | ~v_574 | ~v_435 | ~v_2951 | ~v_2950 | ~v_434 | ~v_2949 | ~v_2948 | ~v_1350 | ~v_3657 | ~v_3656 | ~v_1347 | ~v_3655 | ~v_3654 | ~v_1346 | ~v_1345 | ~v_1344 | ~v_1343 | ~v_1496 | ~v_1495 | ~v_1494 | ~v_1493 | v_3690;
assign x_9584 = v_55 | v_61 | v_59 | v_58 | v_145 | v_143 | v_142 | v_167 | v_166 | v_165 | v_146 | v_183 | ~v_572 | ~v_571 | ~v_2940 | ~v_2937 | ~v_530 | ~v_3036 | ~v_3035 | ~v_529 | ~v_3034 | ~v_3033 | ~v_570 | ~v_569 | ~v_420 | ~v_2936 | ~v_2935 | ~v_419 | ~v_2934 | ~v_2933 | ~v_1325 | ~v_3652 | ~v_3651 | ~v_1322 | ~v_3650 | ~v_3649 | ~v_1321 | ~v_1320 | ~v_1319 | ~v_1318 | ~v_1487 | ~v_1486 | ~v_1485 | ~v_1484 | v_3689;
assign x_9585 = v_18 | v_16 | v_15 | v_12 | ~v_2927 | ~v_2926 | v_135 | v_134 | v_137 | v_138 | v_163 | v_162 | v_161 | v_182 | ~v_567 | ~v_566 | ~v_515 | ~v_3031 | ~v_3030 | ~v_514 | ~v_3029 | ~v_3028 | ~v_565 | ~v_564 | ~v_405 | ~v_2921 | ~v_2920 | ~v_404 | ~v_2919 | ~v_2918 | ~v_1300 | ~v_3647 | ~v_3646 | ~v_1297 | ~v_3645 | ~v_3644 | ~v_1296 | ~v_1295 | ~v_1294 | ~v_1293 | ~v_1478 | ~v_1477 | ~v_1476 | ~v_1475 | v_3688;
assign x_9586 = v_3687 | ~v_3684;
assign x_9587 = v_3687 | ~v_3685;
assign x_9588 = v_3687 | ~v_3686;
assign x_9589 = v_103 | v_101 | v_100 | v_95 | v_102 | v_171 | v_170 | v_169 | v_150 | v_149 | v_148 | v_184 | ~v_2955 | ~v_2952 | ~v_545 | ~v_3041 | ~v_3040 | ~v_544 | ~v_3039 | ~v_3038 | ~v_561 | ~v_560 | ~v_559 | ~v_558 | ~v_387 | ~v_2989 | ~v_2988 | ~v_386 | ~v_2987 | ~v_2986 | ~v_1350 | ~v_3657 | ~v_3656 | ~v_1347 | ~v_3655 | ~v_3654 | ~v_1408 | ~v_1407 | ~v_1406 | ~v_1405 | ~v_1496 | ~v_1495 | ~v_1494 | ~v_1493 | v_3686;
assign x_9590 = v_53 | v_61 | v_60 | v_59 | v_58 | v_144 | v_145 | v_143 | v_167 | v_166 | v_165 | v_183 | ~v_2940 | ~v_2937 | ~v_530 | ~v_3036 | ~v_3035 | ~v_529 | ~v_3034 | ~v_3033 | ~v_556 | ~v_555 | ~v_554 | ~v_553 | ~v_372 | ~v_2984 | ~v_2983 | ~v_371 | ~v_2982 | ~v_2981 | ~v_1325 | ~v_3652 | ~v_3651 | ~v_1322 | ~v_3650 | ~v_3649 | ~v_1399 | ~v_1398 | ~v_1397 | ~v_1396 | ~v_1487 | ~v_1486 | ~v_1485 | ~v_1484 | v_3685;
assign x_9591 = v_18 | v_17 | v_16 | v_15 | v_10 | ~v_2927 | ~v_2926 | v_136 | v_135 | v_137 | v_163 | v_162 | v_161 | v_182 | ~v_515 | ~v_3031 | ~v_3030 | ~v_514 | ~v_3029 | ~v_3028 | ~v_551 | ~v_550 | ~v_549 | ~v_548 | ~v_357 | ~v_2979 | ~v_2978 | ~v_356 | ~v_2977 | ~v_2976 | ~v_1300 | ~v_3647 | ~v_3646 | ~v_1297 | ~v_3645 | ~v_3644 | ~v_1390 | ~v_1389 | ~v_1388 | ~v_1387 | ~v_1478 | ~v_1477 | ~v_1476 | ~v_1475 | v_3684;
assign x_9592 = v_3683 | ~v_3680;
assign x_9593 = v_3683 | ~v_3681;
assign x_9594 = v_3683 | ~v_3682;
assign x_9595 = v_103 | v_100 | v_102 | v_171 | v_170 | v_169 | v_160 | v_150 | v_149 | v_148 | v_147 | v_184 | ~v_2955 | ~v_2952 | ~v_545 | ~v_3041 | ~v_3040 | ~v_544 | ~v_3039 | ~v_3038 | ~v_543 | ~v_542 | ~v_541 | ~v_540 | ~v_297 | ~v_3005 | ~v_3004 | ~v_296 | ~v_3003 | ~v_3002 | ~v_1350 | ~v_3657 | ~v_3656 | ~v_1347 | ~v_3655 | ~v_3654 | ~v_1436 | ~v_1435 | ~v_1434 | ~v_1433 | ~v_1496 | ~v_1495 | ~v_1494 | ~v_1493 | v_3682;
assign x_9596 = v_61 | v_60 | v_58 | v_144 | v_159 | v_145 | v_143 | v_142 | v_167 | v_166 | v_165 | v_183 | ~v_2940 | ~v_2937 | ~v_530 | ~v_3036 | ~v_3035 | ~v_529 | ~v_3034 | ~v_3033 | ~v_528 | ~v_527 | ~v_526 | ~v_525 | ~v_264 | ~v_3000 | ~v_2999 | ~v_263 | ~v_2998 | ~v_2997 | ~v_1325 | ~v_3652 | ~v_3651 | ~v_1322 | ~v_3650 | ~v_3649 | ~v_1427 | ~v_1426 | ~v_1425 | ~v_1424 | ~v_1487 | ~v_1486 | ~v_1485 | ~v_1484 | v_3681;
assign x_9597 = v_18 | v_17 | v_15 | ~v_2927 | ~v_2926 | v_136 | v_135 | v_134 | v_137 | v_163 | v_162 | v_161 | v_155 | v_182 | ~v_515 | ~v_3031 | ~v_3030 | ~v_514 | ~v_3029 | ~v_3028 | ~v_513 | ~v_512 | ~v_511 | ~v_510 | ~v_231 | ~v_2995 | ~v_2994 | ~v_230 | ~v_2993 | ~v_2992 | ~v_1300 | ~v_3647 | ~v_3646 | ~v_1297 | ~v_3645 | ~v_3644 | ~v_1418 | ~v_1417 | ~v_1416 | ~v_1415 | ~v_1478 | ~v_1477 | ~v_1476 | ~v_1475 | v_3680;
assign x_9598 = v_3679 | ~v_3676;
assign x_9599 = v_3679 | ~v_3677;
assign x_9600 = v_3679 | ~v_3678;
assign x_9601 = v_98 | v_103 | v_101 | v_100 | v_93 | v_151 | v_170 | v_150 | v_149 | v_148 | v_147 | v_184 | ~v_299 | ~v_2957 | ~v_2956 | ~v_2955 | ~v_298 | ~v_2954 | ~v_2953 | ~v_2952 | ~v_387 | ~v_2989 | ~v_2988 | ~v_386 | ~v_2987 | ~v_2986 | ~v_499 | ~v_498 | ~v_497 | ~v_496 | ~v_1352 | ~v_1351 | ~v_1350 | ~v_3657 | ~v_3656 | ~v_1349 | ~v_1348 | ~v_1347 | ~v_3655 | ~v_3654 | ~v_1408 | ~v_1407 | ~v_1406 | ~v_1405 | v_3678;
assign x_9602 = v_56 | v_61 | v_51 | v_59 | v_58 | v_144 | v_145 | v_143 | v_142 | v_166 | v_146 | v_183 | ~v_266 | ~v_2942 | ~v_2941 | ~v_2940 | ~v_265 | ~v_2939 | ~v_2938 | ~v_2937 | ~v_372 | ~v_2984 | ~v_2983 | ~v_371 | ~v_2982 | ~v_2981 | ~v_494 | ~v_493 | ~v_492 | ~v_491 | ~v_1327 | ~v_1326 | ~v_1325 | ~v_3652 | ~v_3651 | ~v_1324 | ~v_1323 | ~v_1322 | ~v_3650 | ~v_3649 | ~v_1399 | ~v_1398 | ~v_1397 | ~v_1396 | v_3677;
assign x_9603 = v_13 | v_18 | v_16 | v_8 | v_15 | ~v_2927 | ~v_2926 | v_136 | v_135 | v_134 | v_137 | v_138 | v_162 | v_182 | ~v_233 | ~v_2925 | ~v_2924 | ~v_232 | ~v_2923 | ~v_2922 | ~v_357 | ~v_2979 | ~v_2978 | ~v_356 | ~v_2977 | ~v_2976 | ~v_489 | ~v_488 | ~v_487 | ~v_486 | ~v_1302 | ~v_1301 | ~v_1300 | ~v_3647 | ~v_3646 | ~v_1299 | ~v_1298 | ~v_1297 | ~v_3645 | ~v_3644 | ~v_1390 | ~v_1389 | ~v_1388 | ~v_1387 | v_3676;
assign x_9604 = v_3675 | ~v_3672;
assign x_9605 = v_3675 | ~v_3673;
assign x_9606 = v_3675 | ~v_3674;
assign x_9607 = v_103 | v_101 | v_96 | v_99 | v_102 | v_171 | v_170 | v_169 | v_149 | v_147 | v_184 | v_181 | ~v_483 | ~v_3021 | ~v_3020 | ~v_2955 | ~v_482 | ~v_3019 | ~v_3018 | ~v_2952 | ~v_481 | ~v_480 | ~v_345 | ~v_3073 | ~v_3072 | ~v_479 | ~v_478 | ~v_344 | ~v_3071 | ~v_3070 | ~v_1464 | ~v_1463 | ~v_1350 | ~v_3657 | ~v_3656 | ~v_1462 | ~v_1461 | ~v_1347 | ~v_3655 | ~v_3654 | ~v_1540 | ~v_1539 | ~v_1538 | ~v_1537 | v_3674;
assign x_9608 = v_54 | v_61 | v_60 | v_59 | v_57 | ~v_3016 | v_144 | v_180 | v_142 | v_167 | v_166 | v_165 | v_183 | ~v_3015 | ~v_468 | ~v_2940 | ~v_467 | ~v_3014 | ~v_3013 | ~v_2937 | ~v_466 | ~v_465 | ~v_330 | ~v_3068 | ~v_3067 | ~v_464 | ~v_463 | ~v_329 | ~v_3066 | ~v_3065 | ~v_1455 | ~v_1454 | ~v_1325 | ~v_3652 | ~v_3651 | ~v_1453 | ~v_1452 | ~v_1322 | ~v_3650 | ~v_3649 | ~v_1531 | ~v_1530 | ~v_1529 | ~v_1528 | v_3673;
assign x_9609 = v_18 | v_17 | v_16 | v_14 | v_11 | ~v_453 | ~v_2927 | ~v_452 | ~v_2926 | v_136 | v_134 | v_179 | v_163 | v_162 | v_161 | v_182 | ~v_3011 | ~v_3010 | ~v_3009 | ~v_3008 | ~v_451 | ~v_450 | ~v_315 | ~v_3063 | ~v_3062 | ~v_449 | ~v_448 | ~v_314 | ~v_3061 | ~v_3060 | ~v_1446 | ~v_1445 | ~v_1300 | ~v_3647 | ~v_3646 | ~v_1444 | ~v_1443 | ~v_1297 | ~v_3645 | ~v_3644 | ~v_1522 | ~v_1521 | ~v_1520 | ~v_1519 | v_3672;
assign x_9610 = v_3671 | ~v_3668;
assign x_9611 = v_3671 | ~v_3669;
assign x_9612 = v_3671 | ~v_3670;
assign x_9613 = v_101 | v_97 | v_102 | v_172 | v_171 | v_170 | v_169 | v_150 | v_148 | v_147 | v_184 | v_181 | ~v_437 | ~v_436 | ~v_2955 | ~v_2952 | ~v_435 | ~v_2951 | ~v_2950 | ~v_434 | ~v_2949 | ~v_2948 | ~v_345 | ~v_3073 | ~v_3072 | ~v_344 | ~v_3071 | ~v_3070 | ~v_433 | ~v_432 | ~v_1350 | ~v_3657 | ~v_3656 | ~v_1347 | ~v_3655 | ~v_3654 | ~v_1346 | ~v_1345 | ~v_1344 | ~v_1343 | ~v_1540 | ~v_1539 | ~v_1538 | ~v_1537 | v_3670;
assign x_9614 = v_55 | v_60 | v_59 | v_180 | v_145 | v_143 | v_142 | v_168 | v_167 | v_166 | v_165 | v_183 | ~v_422 | ~v_421 | ~v_2940 | ~v_2937 | ~v_420 | ~v_2936 | ~v_2935 | ~v_419 | ~v_2934 | ~v_2933 | ~v_330 | ~v_3068 | ~v_3067 | ~v_329 | ~v_3066 | ~v_3065 | ~v_418 | ~v_417 | ~v_1325 | ~v_3652 | ~v_3651 | ~v_1322 | ~v_3650 | ~v_3649 | ~v_1321 | ~v_1320 | ~v_1319 | ~v_1318 | ~v_1531 | ~v_1530 | ~v_1529 | ~v_1528 | v_3669;
assign x_9615 = v_17 | v_16 | v_12 | ~v_2927 | ~v_2926 | v_135 | v_134 | v_137 | v_179 | v_164 | v_163 | v_162 | v_161 | v_182 | ~v_407 | ~v_406 | ~v_405 | ~v_2921 | ~v_2920 | ~v_404 | ~v_2919 | ~v_2918 | ~v_315 | ~v_3063 | ~v_3062 | ~v_314 | ~v_3061 | ~v_3060 | ~v_403 | ~v_402 | ~v_1300 | ~v_3647 | ~v_3646 | ~v_1297 | ~v_3645 | ~v_3644 | ~v_1296 | ~v_1295 | ~v_1294 | ~v_1293 | ~v_1522 | ~v_1521 | ~v_1520 | ~v_1519 | v_3668;
assign x_9616 = v_3667 | ~v_3664;
assign x_9617 = v_3667 | ~v_3665;
assign x_9618 = v_3667 | ~v_3666;
assign x_9619 = v_103 | v_101 | v_102 | v_171 | v_170 | v_169 | v_150 | v_149 | v_148 | v_147 | v_184 | v_181 | ~v_391 | ~v_390 | ~v_2955 | ~v_2952 | ~v_387 | ~v_2989 | ~v_2988 | ~v_386 | ~v_2987 | ~v_2986 | ~v_345 | ~v_3073 | ~v_3072 | ~v_344 | ~v_3071 | ~v_3070 | ~v_385 | ~v_384 | ~v_1350 | ~v_3657 | ~v_3656 | ~v_1347 | ~v_3655 | ~v_3654 | ~v_1408 | ~v_1407 | ~v_1406 | ~v_1405 | ~v_1540 | ~v_1539 | ~v_1538 | ~v_1537 | v_3666;
assign x_9620 = v_61 | v_60 | v_59 | v_144 | v_180 | v_145 | v_143 | v_142 | v_167 | v_166 | v_165 | v_183 | ~v_376 | ~v_375 | ~v_2940 | ~v_2937 | ~v_372 | ~v_2984 | ~v_2983 | ~v_371 | ~v_2982 | ~v_2981 | ~v_330 | ~v_3068 | ~v_3067 | ~v_329 | ~v_3066 | ~v_3065 | ~v_370 | ~v_369 | ~v_1325 | ~v_3652 | ~v_3651 | ~v_1322 | ~v_3650 | ~v_3649 | ~v_1399 | ~v_1398 | ~v_1397 | ~v_1396 | ~v_1531 | ~v_1530 | ~v_1529 | ~v_1528 | v_3665;
assign x_9621 = v_18 | v_17 | v_16 | ~v_2927 | ~v_2926 | v_136 | v_135 | v_134 | v_137 | v_179 | v_163 | v_162 | v_161 | v_182 | ~v_361 | ~v_360 | ~v_357 | ~v_2979 | ~v_2978 | ~v_356 | ~v_2977 | ~v_2976 | ~v_315 | ~v_3063 | ~v_3062 | ~v_314 | ~v_3061 | ~v_3060 | ~v_355 | ~v_354 | ~v_1300 | ~v_3647 | ~v_3646 | ~v_1297 | ~v_3645 | ~v_3644 | ~v_1390 | ~v_1389 | ~v_1388 | ~v_1387 | ~v_1522 | ~v_1521 | ~v_1520 | ~v_1519 | v_3664;
assign x_9622 = v_3663 | ~v_3660;
assign x_9623 = v_3663 | ~v_3661;
assign x_9624 = v_3663 | ~v_3662;
assign x_9625 = v_103 | v_95 | v_102 | v_171 | v_170 | v_169 | v_160 | v_150 | v_149 | v_148 | v_184 | v_181 | ~v_2955 | ~v_2952 | ~v_297 | ~v_3005 | ~v_3004 | ~v_296 | ~v_3003 | ~v_3002 | ~v_345 | ~v_3073 | ~v_3072 | ~v_344 | ~v_3071 | ~v_3070 | ~v_343 | ~v_342 | ~v_341 | ~v_340 | ~v_1350 | ~v_3657 | ~v_3656 | ~v_1347 | ~v_3655 | ~v_3654 | ~v_1436 | ~v_1435 | ~v_1434 | ~v_1433 | ~v_1540 | ~v_1539 | ~v_1538 | ~v_1537 | v_3662;
assign x_9626 = v_53 | v_61 | v_60 | v_144 | v_180 | v_159 | v_145 | v_143 | v_167 | v_166 | v_165 | v_183 | ~v_2940 | ~v_2937 | ~v_264 | ~v_3000 | ~v_2999 | ~v_263 | ~v_2998 | ~v_2997 | ~v_330 | ~v_3068 | ~v_3067 | ~v_329 | ~v_3066 | ~v_3065 | ~v_328 | ~v_327 | ~v_326 | ~v_325 | ~v_1325 | ~v_3652 | ~v_3651 | ~v_1322 | ~v_3650 | ~v_3649 | ~v_1427 | ~v_1426 | ~v_1425 | ~v_1424 | ~v_1531 | ~v_1530 | ~v_1529 | ~v_1528 | v_3661;
assign x_9627 = v_18 | v_17 | v_10 | ~v_2927 | ~v_2926 | v_136 | v_135 | v_137 | v_179 | v_163 | v_162 | v_161 | v_155 | v_182 | ~v_231 | ~v_2995 | ~v_2994 | ~v_230 | ~v_2993 | ~v_2992 | ~v_315 | ~v_3063 | ~v_3062 | ~v_314 | ~v_3061 | ~v_3060 | ~v_313 | ~v_312 | ~v_311 | ~v_310 | ~v_1300 | ~v_3647 | ~v_3646 | ~v_1297 | ~v_3645 | ~v_3644 | ~v_1418 | ~v_1417 | ~v_1416 | ~v_1415 | ~v_1522 | ~v_1521 | ~v_1520 | ~v_1519 | v_3660;
assign x_9628 = v_3659 | ~v_3648;
assign x_9629 = v_3659 | ~v_3653;
assign x_9630 = v_3659 | ~v_3658;
assign x_9631 = v_98 | v_103 | v_100 | v_93 | v_102 | v_170 | v_160 | v_150 | v_149 | v_148 | v_147 | v_184 | ~v_299 | ~v_2957 | ~v_2956 | ~v_2955 | ~v_298 | ~v_2954 | ~v_2953 | ~v_2952 | ~v_297 | ~v_3005 | ~v_3004 | ~v_296 | ~v_3003 | ~v_3002 | ~v_295 | ~v_294 | ~v_293 | ~v_292 | ~v_1352 | ~v_1351 | ~v_1350 | ~v_3657 | ~v_3656 | ~v_1349 | ~v_1348 | ~v_1347 | ~v_3655 | ~v_3654 | ~v_1436 | ~v_1435 | ~v_1434 | ~v_1433 | v_3658;
assign x_9632 = v_3657 | v_153;
assign x_9633 = v_3657 | v_123;
assign x_9634 = v_3656 | v_152;
assign x_9635 = v_3656 | v_120;
assign x_9636 = v_3655 | ~v_153;
assign x_9637 = v_3655 | v_108;
assign x_9638 = v_3654 | ~v_152;
assign x_9639 = v_3654 | v_105;
assign x_9640 = v_56 | v_61 | v_51 | v_60 | v_58 | v_144 | v_159 | v_145 | v_143 | v_142 | v_166 | v_183 | ~v_266 | ~v_2942 | ~v_2941 | ~v_2940 | ~v_265 | ~v_2939 | ~v_2938 | ~v_2937 | ~v_264 | ~v_3000 | ~v_2999 | ~v_263 | ~v_2998 | ~v_2997 | ~v_262 | ~v_261 | ~v_260 | ~v_259 | ~v_1327 | ~v_1326 | ~v_1325 | ~v_3652 | ~v_3651 | ~v_1324 | ~v_1323 | ~v_1322 | ~v_3650 | ~v_3649 | ~v_1427 | ~v_1426 | ~v_1425 | ~v_1424 | v_3653;
assign x_9641 = v_3652 | v_153;
assign x_9642 = v_3652 | v_81;
assign x_9643 = v_3651 | v_152;
assign x_9644 = v_3651 | v_78;
assign x_9645 = v_3650 | ~v_153;
assign x_9646 = v_3650 | v_66;
assign x_9647 = v_3649 | ~v_152;
assign x_9648 = v_3649 | v_63;
assign x_9649 = v_13 | v_18 | v_17 | v_8 | v_15 | ~v_2927 | ~v_2926 | v_136 | v_135 | v_134 | v_137 | v_162 | v_155 | v_182 | ~v_233 | ~v_2925 | ~v_2924 | ~v_232 | ~v_2923 | ~v_2922 | ~v_231 | ~v_2995 | ~v_2994 | ~v_230 | ~v_2993 | ~v_2992 | ~v_229 | ~v_228 | ~v_227 | ~v_226 | ~v_1302 | ~v_1301 | ~v_1300 | ~v_3647 | ~v_3646 | ~v_1299 | ~v_1298 | ~v_1297 | ~v_3645 | ~v_3644 | ~v_1418 | ~v_1417 | ~v_1416 | ~v_1415 | v_3648;
assign x_9650 = v_3647 | v_153;
assign x_9651 = v_3647 | v_39;
assign x_9652 = v_3646 | v_152;
assign x_9653 = v_3646 | v_36;
assign x_9654 = v_3645 | ~v_153;
assign x_9655 = v_3645 | v_24;
assign x_9656 = v_3644 | ~v_152;
assign x_9657 = v_3644 | v_21;
assign x_9658 = v_3643 | ~v_3641;
assign x_9659 = v_3643 | ~v_3642;
assign x_9660 = v_3643 | ~v_1274;
assign x_9661 = v_3643 | ~v_1275;
assign x_9662 = v_3643 | ~v_153;
assign x_9663 = v_3643 | ~v_152;
assign x_9664 = ~v_186 | ~v_1272 | v_3642;
assign x_9665 = ~v_185 | ~v_1851 | v_3641;
assign x_9666 = v_3640 | ~v_3457;
assign x_9667 = v_3640 | ~v_3639;
assign x_9668 = v_157 | v_156 | ~v_3638 | ~v_738 | ~v_736 | ~v_3459 | ~v_3458 | v_3639;
assign x_9669 = v_3638 | ~v_3505;
assign x_9670 = v_3638 | ~v_3521;
assign x_9671 = v_3638 | ~v_3537;
assign x_9672 = v_3638 | ~v_3553;
assign x_9673 = v_3638 | ~v_3569;
assign x_9674 = v_3638 | ~v_3573;
assign x_9675 = v_3638 | ~v_3589;
assign x_9676 = v_3638 | ~v_3593;
assign x_9677 = v_3638 | ~v_3597;
assign x_9678 = v_3638 | ~v_3601;
assign x_9679 = v_3638 | ~v_3605;
assign x_9680 = v_3638 | ~v_3621;
assign x_9681 = v_3638 | ~v_3625;
assign x_9682 = v_3638 | ~v_3629;
assign x_9683 = v_3638 | ~v_3633;
assign x_9684 = v_3638 | ~v_3637;
assign x_9685 = v_3638 | ~v_1263;
assign x_9686 = v_3638 | ~v_1264;
assign x_9687 = v_3638 | ~v_1265;
assign x_9688 = v_3638 | ~v_1266;
assign x_9689 = ~v_3636 | ~v_3635 | ~v_3634 | v_3637;
assign x_9690 = v_3636 | ~v_1626;
assign x_9691 = v_3636 | ~v_3490;
assign x_9692 = v_3636 | ~v_1627;
assign x_9693 = v_3636 | ~v_1746;
assign x_9694 = v_3636 | ~v_3491;
assign x_9695 = v_3636 | ~v_1628;
assign x_9696 = v_3636 | ~v_1747;
assign x_9697 = v_3636 | ~v_1629;
assign x_9698 = v_3636 | ~v_3492;
assign x_9699 = v_3636 | ~v_1630;
assign x_9700 = v_3636 | ~v_1748;
assign x_9701 = v_3636 | ~v_3493;
assign x_9702 = v_3636 | ~v_1631;
assign x_9703 = v_3636 | ~v_1749;
assign x_9704 = v_3636 | ~v_3496;
assign x_9705 = v_3636 | ~v_3497;
assign x_9706 = v_3636 | ~v_3564;
assign x_9707 = v_3636 | ~v_3498;
assign x_9708 = v_3636 | ~v_3565;
assign x_9709 = v_3636 | ~v_3499;
assign x_9710 = v_3636 | ~v_3500;
assign x_9711 = v_3636 | ~v_3566;
assign x_9712 = v_3636 | ~v_3501;
assign x_9713 = v_3636 | ~v_3567;
assign x_9714 = v_3636 | ~v_839;
assign x_9715 = v_3636 | ~v_1257;
assign x_9716 = v_3636 | ~v_1023;
assign x_9717 = v_3636 | ~v_840;
assign x_9718 = v_3636 | ~v_1258;
assign x_9719 = v_3636 | ~v_1024;
assign x_9720 = v_3636 | ~v_184;
assign x_9721 = v_3636 | ~v_169;
assign x_9722 = v_3636 | ~v_148;
assign x_9723 = v_3636 | ~v_1259;
assign x_9724 = v_3636 | ~v_1260;
assign x_9725 = v_3636 | ~v_103;
assign x_9726 = v_3636 | ~v_102;
assign x_9727 = v_3636 | ~v_101;
assign x_9728 = v_3636 | ~v_100;
assign x_9729 = v_3636 | ~v_99;
assign x_9730 = v_3636 | ~v_98;
assign x_9731 = v_3636 | ~v_97;
assign x_9732 = v_3636 | ~v_95;
assign x_9733 = v_3636 | ~v_94;
assign x_9734 = v_3635 | ~v_1601;
assign x_9735 = v_3635 | ~v_3475;
assign x_9736 = v_3635 | ~v_1602;
assign x_9737 = v_3635 | ~v_1737;
assign x_9738 = v_3635 | ~v_3476;
assign x_9739 = v_3635 | ~v_1603;
assign x_9740 = v_3635 | ~v_1738;
assign x_9741 = v_3635 | ~v_1604;
assign x_9742 = v_3635 | ~v_3477;
assign x_9743 = v_3635 | ~v_1605;
assign x_9744 = v_3635 | ~v_1739;
assign x_9745 = v_3635 | ~v_3478;
assign x_9746 = v_3635 | ~v_1606;
assign x_9747 = v_3635 | ~v_1740;
assign x_9748 = v_3635 | ~v_3481;
assign x_9749 = v_3635 | ~v_3482;
assign x_9750 = v_3635 | ~v_3559;
assign x_9751 = v_3635 | ~v_3483;
assign x_9752 = v_3635 | ~v_3560;
assign x_9753 = v_3635 | ~v_3484;
assign x_9754 = v_3635 | ~v_3485;
assign x_9755 = v_3635 | ~v_806;
assign x_9756 = v_3635 | ~v_1252;
assign x_9757 = v_3635 | ~v_1008;
assign x_9758 = v_3635 | ~v_1253;
assign x_9759 = v_3635 | ~v_1009;
assign x_9760 = v_3635 | ~v_3561;
assign x_9761 = v_3635 | ~v_807;
assign x_9762 = v_3635 | ~v_3486;
assign x_9763 = v_3635 | ~v_3562;
assign x_9764 = v_3635 | ~v_183;
assign x_9765 = v_3635 | ~v_165;
assign x_9766 = v_3635 | ~v_143;
assign x_9767 = v_3635 | ~v_1254;
assign x_9768 = v_3635 | ~v_1255;
assign x_9769 = v_3635 | ~v_61;
assign x_9770 = v_3635 | ~v_60;
assign x_9771 = v_3635 | ~v_59;
assign x_9772 = v_3635 | ~v_58;
assign x_9773 = v_3635 | ~v_57;
assign x_9774 = v_3635 | ~v_56;
assign x_9775 = v_3635 | ~v_55;
assign x_9776 = v_3635 | ~v_53;
assign x_9777 = v_3635 | ~v_52;
assign x_9778 = v_3634 | ~v_1576;
assign x_9779 = v_3634 | ~v_3460;
assign x_9780 = v_3634 | ~v_1577;
assign x_9781 = v_3634 | ~v_1728;
assign x_9782 = v_3634 | ~v_3461;
assign x_9783 = v_3634 | ~v_1578;
assign x_9784 = v_3634 | ~v_1729;
assign x_9785 = v_3634 | ~v_1579;
assign x_9786 = v_3634 | ~v_3462;
assign x_9787 = v_3634 | ~v_1580;
assign x_9788 = v_3634 | ~v_1730;
assign x_9789 = v_3634 | ~v_3463;
assign x_9790 = v_3634 | ~v_1581;
assign x_9791 = v_3634 | ~v_1731;
assign x_9792 = v_3634 | ~v_3466;
assign x_9793 = v_3634 | ~v_3467;
assign x_9794 = v_3634 | ~v_3554;
assign x_9795 = v_3634 | ~v_3468;
assign x_9796 = v_3634 | ~v_3555;
assign x_9797 = v_3634 | ~v_3469;
assign x_9798 = v_3634 | ~v_3556;
assign x_9799 = v_3634 | ~v_3470;
assign x_9800 = v_3634 | ~v_3557;
assign x_9801 = v_3634 | ~v_773;
assign x_9802 = v_3634 | ~v_774;
assign x_9803 = v_3634 | ~v_182;
assign x_9804 = v_3634 | ~v_161;
assign x_9805 = v_3634 | ~v_3473;
assign x_9806 = v_3634 | ~v_1247;
assign x_9807 = v_3634 | ~v_1248;
assign x_9808 = v_3634 | ~v_135;
assign x_9809 = v_3634 | ~v_1249;
assign x_9810 = v_3634 | ~v_993;
assign x_9811 = v_3634 | ~v_1250;
assign x_9812 = v_3634 | ~v_994;
assign x_9813 = v_3634 | ~v_18;
assign x_9814 = v_3634 | ~v_17;
assign x_9815 = v_3634 | ~v_16;
assign x_9816 = v_3634 | ~v_15;
assign x_9817 = v_3634 | ~v_14;
assign x_9818 = v_3634 | ~v_13;
assign x_9819 = v_3634 | ~v_12;
assign x_9820 = v_3634 | ~v_10;
assign x_9821 = v_3634 | ~v_9;
assign x_9822 = ~v_3632 | ~v_3631 | ~v_3630 | v_3633;
assign x_9823 = v_3632 | ~v_1822;
assign x_9824 = v_3632 | ~v_1823;
assign x_9825 = v_3632 | ~v_1824;
assign x_9826 = v_3632 | ~v_1825;
assign x_9827 = v_3632 | ~v_1626;
assign x_9828 = v_3632 | ~v_3490;
assign x_9829 = v_3632 | ~v_1746;
assign x_9830 = v_3632 | ~v_3491;
assign x_9831 = v_3632 | ~v_1747;
assign x_9832 = v_3632 | ~v_1629;
assign x_9833 = v_3632 | ~v_3492;
assign x_9834 = v_3632 | ~v_1748;
assign x_9835 = v_3632 | ~v_3493;
assign x_9836 = v_3632 | ~v_1749;
assign x_9837 = v_3632 | ~v_3616;
assign x_9838 = v_3632 | ~v_3617;
assign x_9839 = v_3632 | ~v_3618;
assign x_9840 = v_3632 | ~v_3619;
assign x_9841 = v_3632 | ~v_3496;
assign x_9842 = v_3632 | ~v_3564;
assign x_9843 = v_3632 | ~v_3565;
assign x_9844 = v_3632 | ~v_3499;
assign x_9845 = v_3632 | ~v_3566;
assign x_9846 = v_3632 | ~v_3567;
assign x_9847 = v_3632 | ~v_885;
assign x_9848 = v_3632 | ~v_1019;
assign x_9849 = v_3632 | ~v_1020;
assign x_9850 = v_3632 | ~v_886;
assign x_9851 = v_3632 | ~v_1021;
assign x_9852 = v_3632 | ~v_1022;
assign x_9853 = v_3632 | ~v_1023;
assign x_9854 = v_3632 | ~v_1024;
assign x_9855 = v_3632 | ~v_184;
assign x_9856 = v_3632 | ~v_181;
assign x_9857 = v_3632 | ~v_171;
assign x_9858 = v_3632 | ~v_170;
assign x_9859 = v_3632 | ~v_148;
assign x_9860 = v_3632 | ~v_147;
assign x_9861 = v_3632 | ~v_103;
assign x_9862 = v_3632 | ~v_102;
assign x_9863 = v_3632 | ~v_101;
assign x_9864 = v_3632 | ~v_99;
assign x_9865 = v_3632 | ~v_97;
assign x_9866 = v_3632 | ~v_93;
assign x_9867 = v_3631 | ~v_1813;
assign x_9868 = v_3631 | ~v_1814;
assign x_9869 = v_3631 | ~v_1815;
assign x_9870 = v_3631 | ~v_1816;
assign x_9871 = v_3631 | ~v_1601;
assign x_9872 = v_3631 | ~v_3475;
assign x_9873 = v_3631 | ~v_1737;
assign x_9874 = v_3631 | ~v_3476;
assign x_9875 = v_3631 | ~v_1738;
assign x_9876 = v_3631 | ~v_1604;
assign x_9877 = v_3631 | ~v_3477;
assign x_9878 = v_3631 | ~v_1739;
assign x_9879 = v_3631 | ~v_3478;
assign x_9880 = v_3631 | ~v_1740;
assign x_9881 = v_3631 | ~v_3611;
assign x_9882 = v_3631 | ~v_3612;
assign x_9883 = v_3631 | ~v_3613;
assign x_9884 = v_3631 | ~v_3614;
assign x_9885 = v_3631 | ~v_3481;
assign x_9886 = v_3631 | ~v_3559;
assign x_9887 = v_3631 | ~v_3560;
assign x_9888 = v_3631 | ~v_3484;
assign x_9889 = v_3631 | ~v_870;
assign x_9890 = v_3631 | ~v_1004;
assign x_9891 = v_3631 | ~v_1005;
assign x_9892 = v_3631 | ~v_871;
assign x_9893 = v_3631 | ~v_1006;
assign x_9894 = v_3631 | ~v_1007;
assign x_9895 = v_3631 | ~v_1008;
assign x_9896 = v_3631 | ~v_1009;
assign x_9897 = v_3631 | ~v_3561;
assign x_9898 = v_3631 | ~v_3562;
assign x_9899 = v_3631 | ~v_183;
assign x_9900 = v_3631 | ~v_180;
assign x_9901 = v_3631 | ~v_167;
assign x_9902 = v_3631 | ~v_166;
assign x_9903 = v_3631 | ~v_143;
assign x_9904 = v_3631 | ~v_142;
assign x_9905 = v_3631 | ~v_61;
assign x_9906 = v_3631 | ~v_60;
assign x_9907 = v_3631 | ~v_59;
assign x_9908 = v_3631 | ~v_57;
assign x_9909 = v_3631 | ~v_55;
assign x_9910 = v_3631 | ~v_51;
assign x_9911 = v_3630 | ~v_1804;
assign x_9912 = v_3630 | ~v_1805;
assign x_9913 = v_3630 | ~v_1806;
assign x_9914 = v_3630 | ~v_1807;
assign x_9915 = v_3630 | ~v_1576;
assign x_9916 = v_3630 | ~v_3460;
assign x_9917 = v_3630 | ~v_1728;
assign x_9918 = v_3630 | ~v_3461;
assign x_9919 = v_3630 | ~v_1729;
assign x_9920 = v_3630 | ~v_1579;
assign x_9921 = v_3630 | ~v_3462;
assign x_9922 = v_3630 | ~v_1730;
assign x_9923 = v_3630 | ~v_3463;
assign x_9924 = v_3630 | ~v_1731;
assign x_9925 = v_3630 | ~v_3606;
assign x_9926 = v_3630 | ~v_3607;
assign x_9927 = v_3630 | ~v_3608;
assign x_9928 = v_3630 | ~v_3609;
assign x_9929 = v_3630 | ~v_3466;
assign x_9930 = v_3630 | ~v_3554;
assign x_9931 = v_3630 | ~v_3555;
assign x_9932 = v_3630 | ~v_3469;
assign x_9933 = v_3630 | ~v_3556;
assign x_9934 = v_3630 | ~v_3557;
assign x_9935 = v_3630 | ~v_855;
assign x_9936 = v_3630 | ~v_989;
assign x_9937 = v_3630 | ~v_990;
assign x_9938 = v_3630 | ~v_856;
assign x_9939 = v_3630 | ~v_991;
assign x_9940 = v_3630 | ~v_992;
assign x_9941 = v_3630 | ~v_182;
assign x_9942 = v_3630 | ~v_179;
assign x_9943 = v_3630 | ~v_163;
assign x_9944 = v_3630 | ~v_162;
assign x_9945 = v_3630 | ~v_135;
assign x_9946 = v_3630 | ~v_134;
assign x_9947 = v_3630 | ~v_993;
assign x_9948 = v_3630 | ~v_994;
assign x_9949 = v_3630 | ~v_18;
assign x_9950 = v_3630 | ~v_17;
assign x_9951 = v_3630 | ~v_16;
assign x_9952 = v_3630 | ~v_14;
assign x_9953 = v_3630 | ~v_12;
assign x_9954 = v_3630 | ~v_8;
assign x_9955 = ~v_3628 | ~v_3627 | ~v_3626 | v_3629;
assign x_9956 = v_3628 | ~v_1718;
assign x_9957 = v_3628 | ~v_1719;
assign x_9958 = v_3628 | ~v_1720;
assign x_9959 = v_3628 | ~v_1721;
assign x_9960 = v_3628 | ~v_1822;
assign x_9961 = v_3628 | ~v_1823;
assign x_9962 = v_3628 | ~v_1824;
assign x_9963 = v_3628 | ~v_1825;
assign x_9964 = v_3628 | ~v_1626;
assign x_9965 = v_3628 | ~v_3490;
assign x_9966 = v_3628 | ~v_3491;
assign x_9967 = v_3628 | ~v_1629;
assign x_9968 = v_3628 | ~v_3492;
assign x_9969 = v_3628 | ~v_3493;
assign x_9970 = v_3628 | ~v_3616;
assign x_9971 = v_3628 | ~v_3617;
assign x_9972 = v_3628 | ~v_3618;
assign x_9973 = v_3628 | ~v_3619;
assign x_9974 = v_3628 | ~v_3548;
assign x_9975 = v_3628 | ~v_3549;
assign x_9976 = v_3628 | ~v_3550;
assign x_9977 = v_3628 | ~v_3551;
assign x_9978 = v_3628 | ~v_3496;
assign x_9979 = v_3628 | ~v_3499;
assign x_9980 = v_3628 | ~v_881;
assign x_9981 = v_3628 | ~v_882;
assign x_9982 = v_3628 | ~v_883;
assign x_9983 = v_3628 | ~v_884;
assign x_9984 = v_3628 | ~v_885;
assign x_9985 = v_3628 | ~v_886;
assign x_9986 = v_3628 | ~v_837;
assign x_9987 = v_3628 | ~v_838;
assign x_9988 = v_3628 | ~v_184;
assign x_9989 = v_3628 | ~v_181;
assign x_9990 = v_3628 | ~v_171;
assign x_9991 = v_3628 | ~v_170;
assign x_9992 = v_3628 | ~v_160;
assign x_9993 = v_3628 | ~v_150;
assign x_9994 = v_3628 | ~v_149;
assign x_9995 = v_3628 | ~v_103;
assign x_9996 = v_3628 | ~v_102;
assign x_9997 = v_3628 | ~v_96;
assign x_9998 = v_3628 | ~v_95;
assign x_9999 = v_3628 | ~v_93;
assign x_10000 = v_3627 | ~v_1709;
assign x_10001 = v_3627 | ~v_1710;
assign x_10002 = v_3627 | ~v_1711;
assign x_10003 = v_3627 | ~v_1712;
assign x_10004 = v_3627 | ~v_1813;
assign x_10005 = v_3627 | ~v_1814;
assign x_10006 = v_3627 | ~v_1815;
assign x_10007 = v_3627 | ~v_1816;
assign x_10008 = v_3627 | ~v_1601;
assign x_10009 = v_3627 | ~v_3475;
assign x_10010 = v_3627 | ~v_3476;
assign x_10011 = v_3627 | ~v_1604;
assign x_10012 = v_3627 | ~v_3477;
assign x_10013 = v_3627 | ~v_3478;
assign x_10014 = v_3627 | ~v_3611;
assign x_10015 = v_3627 | ~v_3612;
assign x_10016 = v_3627 | ~v_3613;
assign x_10017 = v_3627 | ~v_3614;
assign x_10018 = v_3627 | ~v_3543;
assign x_10019 = v_3627 | ~v_3544;
assign x_10020 = v_3627 | ~v_3545;
assign x_10021 = v_3627 | ~v_3546;
assign x_10022 = v_3627 | ~v_3481;
assign x_10023 = v_3627 | ~v_3484;
assign x_10024 = v_3627 | ~v_866;
assign x_10025 = v_3627 | ~v_867;
assign x_10026 = v_3627 | ~v_868;
assign x_10027 = v_3627 | ~v_869;
assign x_10028 = v_3627 | ~v_870;
assign x_10029 = v_3627 | ~v_871;
assign x_10030 = v_3627 | ~v_804;
assign x_10031 = v_3627 | ~v_805;
assign x_10032 = v_3627 | ~v_183;
assign x_10033 = v_3627 | ~v_180;
assign x_10034 = v_3627 | ~v_167;
assign x_10035 = v_3627 | ~v_166;
assign x_10036 = v_3627 | ~v_159;
assign x_10037 = v_3627 | ~v_145;
assign x_10038 = v_3627 | ~v_144;
assign x_10039 = v_3627 | ~v_61;
assign x_10040 = v_3627 | ~v_60;
assign x_10041 = v_3627 | ~v_54;
assign x_10042 = v_3627 | ~v_53;
assign x_10043 = v_3627 | ~v_51;
assign x_10044 = v_3626 | ~v_1700;
assign x_10045 = v_3626 | ~v_1701;
assign x_10046 = v_3626 | ~v_1702;
assign x_10047 = v_3626 | ~v_1703;
assign x_10048 = v_3626 | ~v_1804;
assign x_10049 = v_3626 | ~v_1805;
assign x_10050 = v_3626 | ~v_1806;
assign x_10051 = v_3626 | ~v_1807;
assign x_10052 = v_3626 | ~v_1576;
assign x_10053 = v_3626 | ~v_3460;
assign x_10054 = v_3626 | ~v_3461;
assign x_10055 = v_3626 | ~v_1579;
assign x_10056 = v_3626 | ~v_3462;
assign x_10057 = v_3626 | ~v_3463;
assign x_10058 = v_3626 | ~v_3606;
assign x_10059 = v_3626 | ~v_3607;
assign x_10060 = v_3626 | ~v_3608;
assign x_10061 = v_3626 | ~v_3609;
assign x_10062 = v_3626 | ~v_3538;
assign x_10063 = v_3626 | ~v_3539;
assign x_10064 = v_3626 | ~v_3540;
assign x_10065 = v_3626 | ~v_3541;
assign x_10066 = v_3626 | ~v_3466;
assign x_10067 = v_3626 | ~v_3469;
assign x_10068 = v_3626 | ~v_851;
assign x_10069 = v_3626 | ~v_852;
assign x_10070 = v_3626 | ~v_853;
assign x_10071 = v_3626 | ~v_854;
assign x_10072 = v_3626 | ~v_855;
assign x_10073 = v_3626 | ~v_856;
assign x_10074 = v_3626 | ~v_771;
assign x_10075 = v_3626 | ~v_772;
assign x_10076 = v_3626 | ~v_182;
assign x_10077 = v_3626 | ~v_179;
assign x_10078 = v_3626 | ~v_163;
assign x_10079 = v_3626 | ~v_162;
assign x_10080 = v_3626 | ~v_155;
assign x_10081 = v_3626 | ~v_137;
assign x_10082 = v_3626 | ~v_136;
assign x_10083 = v_3626 | ~v_18;
assign x_10084 = v_3626 | ~v_17;
assign x_10085 = v_3626 | ~v_11;
assign x_10086 = v_3626 | ~v_10;
assign x_10087 = v_3626 | ~v_8;
assign x_10088 = ~v_3624 | ~v_3623 | ~v_3622 | v_3625;
assign x_10089 = v_3624 | ~v_1690;
assign x_10090 = v_3624 | ~v_1691;
assign x_10091 = v_3624 | ~v_1692;
assign x_10092 = v_3624 | ~v_1693;
assign x_10093 = v_3624 | ~v_1822;
assign x_10094 = v_3624 | ~v_1823;
assign x_10095 = v_3624 | ~v_1824;
assign x_10096 = v_3624 | ~v_1825;
assign x_10097 = v_3624 | ~v_1626;
assign x_10098 = v_3624 | ~v_3490;
assign x_10099 = v_3624 | ~v_3491;
assign x_10100 = v_3624 | ~v_1629;
assign x_10101 = v_3624 | ~v_3492;
assign x_10102 = v_3624 | ~v_3493;
assign x_10103 = v_3624 | ~v_3616;
assign x_10104 = v_3624 | ~v_3617;
assign x_10105 = v_3624 | ~v_3618;
assign x_10106 = v_3624 | ~v_3619;
assign x_10107 = v_3624 | ~v_3532;
assign x_10108 = v_3624 | ~v_3533;
assign x_10109 = v_3624 | ~v_3534;
assign x_10110 = v_3624 | ~v_3535;
assign x_10111 = v_3624 | ~v_3496;
assign x_10112 = v_3624 | ~v_3499;
assign x_10113 = v_3624 | ~v_925;
assign x_10114 = v_3624 | ~v_926;
assign x_10115 = v_3624 | ~v_885;
assign x_10116 = v_3624 | ~v_886;
assign x_10117 = v_3624 | ~v_927;
assign x_10118 = v_3624 | ~v_928;
assign x_10119 = v_3624 | ~v_929;
assign x_10120 = v_3624 | ~v_930;
assign x_10121 = v_3624 | ~v_184;
assign x_10122 = v_3624 | ~v_181;
assign x_10123 = v_3624 | ~v_171;
assign x_10124 = v_3624 | ~v_170;
assign x_10125 = v_3624 | ~v_150;
assign x_10126 = v_3624 | ~v_149;
assign x_10127 = v_3624 | ~v_148;
assign x_10128 = v_3624 | ~v_147;
assign x_10129 = v_3624 | ~v_103;
assign x_10130 = v_3624 | ~v_102;
assign x_10131 = v_3624 | ~v_101;
assign x_10132 = v_3624 | ~v_93;
assign x_10133 = v_3623 | ~v_1681;
assign x_10134 = v_3623 | ~v_1682;
assign x_10135 = v_3623 | ~v_1683;
assign x_10136 = v_3623 | ~v_1684;
assign x_10137 = v_3623 | ~v_1813;
assign x_10138 = v_3623 | ~v_1814;
assign x_10139 = v_3623 | ~v_1815;
assign x_10140 = v_3623 | ~v_1816;
assign x_10141 = v_3623 | ~v_1601;
assign x_10142 = v_3623 | ~v_3475;
assign x_10143 = v_3623 | ~v_3476;
assign x_10144 = v_3623 | ~v_1604;
assign x_10145 = v_3623 | ~v_3477;
assign x_10146 = v_3623 | ~v_3478;
assign x_10147 = v_3623 | ~v_3611;
assign x_10148 = v_3623 | ~v_3612;
assign x_10149 = v_3623 | ~v_3613;
assign x_10150 = v_3623 | ~v_3614;
assign x_10151 = v_3623 | ~v_3527;
assign x_10152 = v_3623 | ~v_3528;
assign x_10153 = v_3623 | ~v_3529;
assign x_10154 = v_3623 | ~v_3530;
assign x_10155 = v_3623 | ~v_3481;
assign x_10156 = v_3623 | ~v_3484;
assign x_10157 = v_3623 | ~v_910;
assign x_10158 = v_3623 | ~v_911;
assign x_10159 = v_3623 | ~v_870;
assign x_10160 = v_3623 | ~v_871;
assign x_10161 = v_3623 | ~v_912;
assign x_10162 = v_3623 | ~v_913;
assign x_10163 = v_3623 | ~v_914;
assign x_10164 = v_3623 | ~v_915;
assign x_10165 = v_3623 | ~v_183;
assign x_10166 = v_3623 | ~v_180;
assign x_10167 = v_3623 | ~v_167;
assign x_10168 = v_3623 | ~v_166;
assign x_10169 = v_3623 | ~v_145;
assign x_10170 = v_3623 | ~v_144;
assign x_10171 = v_3623 | ~v_143;
assign x_10172 = v_3623 | ~v_142;
assign x_10173 = v_3623 | ~v_61;
assign x_10174 = v_3623 | ~v_60;
assign x_10175 = v_3623 | ~v_59;
assign x_10176 = v_3623 | ~v_51;
assign x_10177 = v_3622 | ~v_1672;
assign x_10178 = v_3622 | ~v_1673;
assign x_10179 = v_3622 | ~v_1674;
assign x_10180 = v_3622 | ~v_1675;
assign x_10181 = v_3622 | ~v_1804;
assign x_10182 = v_3622 | ~v_1805;
assign x_10183 = v_3622 | ~v_1806;
assign x_10184 = v_3622 | ~v_1807;
assign x_10185 = v_3622 | ~v_1576;
assign x_10186 = v_3622 | ~v_3460;
assign x_10187 = v_3622 | ~v_3461;
assign x_10188 = v_3622 | ~v_1579;
assign x_10189 = v_3622 | ~v_3462;
assign x_10190 = v_3622 | ~v_3463;
assign x_10191 = v_3622 | ~v_3606;
assign x_10192 = v_3622 | ~v_3607;
assign x_10193 = v_3622 | ~v_3608;
assign x_10194 = v_3622 | ~v_3609;
assign x_10195 = v_3622 | ~v_3522;
assign x_10196 = v_3622 | ~v_3523;
assign x_10197 = v_3622 | ~v_3524;
assign x_10198 = v_3622 | ~v_3525;
assign x_10199 = v_3622 | ~v_3466;
assign x_10200 = v_3622 | ~v_3469;
assign x_10201 = v_3622 | ~v_895;
assign x_10202 = v_3622 | ~v_896;
assign x_10203 = v_3622 | ~v_855;
assign x_10204 = v_3622 | ~v_856;
assign x_10205 = v_3622 | ~v_897;
assign x_10206 = v_3622 | ~v_898;
assign x_10207 = v_3622 | ~v_899;
assign x_10208 = v_3622 | ~v_900;
assign x_10209 = v_3622 | ~v_182;
assign x_10210 = v_3622 | ~v_179;
assign x_10211 = v_3622 | ~v_163;
assign x_10212 = v_3622 | ~v_162;
assign x_10213 = v_3622 | ~v_137;
assign x_10214 = v_3622 | ~v_136;
assign x_10215 = v_3622 | ~v_135;
assign x_10216 = v_3622 | ~v_134;
assign x_10217 = v_3622 | ~v_18;
assign x_10218 = v_3622 | ~v_17;
assign x_10219 = v_3622 | ~v_16;
assign x_10220 = v_3622 | ~v_8;
assign x_10221 = ~v_3620 | ~v_3615 | ~v_3610 | v_3621;
assign x_10222 = v_3620 | ~v_1622;
assign x_10223 = v_3620 | ~v_1623;
assign x_10224 = v_3620 | ~v_1624;
assign x_10225 = v_3620 | ~v_1625;
assign x_10226 = v_3620 | ~v_1822;
assign x_10227 = v_3620 | ~v_1823;
assign x_10228 = v_3620 | ~v_1824;
assign x_10229 = v_3620 | ~v_1825;
assign x_10230 = v_3620 | ~v_1626;
assign x_10231 = v_3620 | ~v_3490;
assign x_10232 = v_3620 | ~v_3491;
assign x_10233 = v_3620 | ~v_1629;
assign x_10234 = v_3620 | ~v_3492;
assign x_10235 = v_3620 | ~v_3493;
assign x_10236 = v_3620 | ~v_3616;
assign x_10237 = v_3620 | ~v_3617;
assign x_10238 = v_3620 | ~v_3618;
assign x_10239 = v_3620 | ~v_3619;
assign x_10240 = v_3620 | ~v_3494;
assign x_10241 = v_3620 | ~v_3495;
assign x_10242 = v_3620 | ~v_3496;
assign x_10243 = v_3620 | ~v_3499;
assign x_10244 = v_3620 | ~v_973;
assign x_10245 = v_3620 | ~v_974;
assign x_10246 = v_3620 | ~v_885;
assign x_10247 = v_3620 | ~v_886;
assign x_10248 = v_3620 | ~v_975;
assign x_10249 = v_3620 | ~v_976;
assign x_10250 = v_3620 | ~v_977;
assign x_10251 = v_3620 | ~v_978;
assign x_10252 = v_3620 | ~v_3502;
assign x_10253 = v_3620 | ~v_3503;
assign x_10254 = v_3620 | ~v_184;
assign x_10255 = v_3620 | ~v_181;
assign x_10256 = v_3620 | ~v_172;
assign x_10257 = v_3620 | ~v_171;
assign x_10258 = v_3620 | ~v_170;
assign x_10259 = v_3620 | ~v_150;
assign x_10260 = v_3620 | ~v_149;
assign x_10261 = v_3620 | ~v_148;
assign x_10262 = v_3620 | ~v_147;
assign x_10263 = v_3620 | ~v_102;
assign x_10264 = v_3620 | ~v_101;
assign x_10265 = v_3620 | ~v_93;
assign x_10266 = ~v_128 | ~v_157 | v_3619;
assign x_10267 = ~v_125 | ~v_156 | v_3618;
assign x_10268 = ~v_113 | v_157 | v_3617;
assign x_10269 = ~v_110 | v_156 | v_3616;
assign x_10270 = v_3615 | ~v_1597;
assign x_10271 = v_3615 | ~v_1598;
assign x_10272 = v_3615 | ~v_1599;
assign x_10273 = v_3615 | ~v_1600;
assign x_10274 = v_3615 | ~v_1813;
assign x_10275 = v_3615 | ~v_1814;
assign x_10276 = v_3615 | ~v_1815;
assign x_10277 = v_3615 | ~v_1816;
assign x_10278 = v_3615 | ~v_1601;
assign x_10279 = v_3615 | ~v_3475;
assign x_10280 = v_3615 | ~v_3476;
assign x_10281 = v_3615 | ~v_1604;
assign x_10282 = v_3615 | ~v_3477;
assign x_10283 = v_3615 | ~v_3478;
assign x_10284 = v_3615 | ~v_3611;
assign x_10285 = v_3615 | ~v_3612;
assign x_10286 = v_3615 | ~v_3613;
assign x_10287 = v_3615 | ~v_3614;
assign x_10288 = v_3615 | ~v_3479;
assign x_10289 = v_3615 | ~v_3480;
assign x_10290 = v_3615 | ~v_3481;
assign x_10291 = v_3615 | ~v_3484;
assign x_10292 = v_3615 | ~v_958;
assign x_10293 = v_3615 | ~v_959;
assign x_10294 = v_3615 | ~v_870;
assign x_10295 = v_3615 | ~v_871;
assign x_10296 = v_3615 | ~v_960;
assign x_10297 = v_3615 | ~v_961;
assign x_10298 = v_3615 | ~v_962;
assign x_10299 = v_3615 | ~v_963;
assign x_10300 = v_3615 | ~v_3487;
assign x_10301 = v_3615 | ~v_3488;
assign x_10302 = v_3615 | ~v_183;
assign x_10303 = v_3615 | ~v_180;
assign x_10304 = v_3615 | ~v_168;
assign x_10305 = v_3615 | ~v_167;
assign x_10306 = v_3615 | ~v_166;
assign x_10307 = v_3615 | ~v_145;
assign x_10308 = v_3615 | ~v_144;
assign x_10309 = v_3615 | ~v_143;
assign x_10310 = v_3615 | ~v_142;
assign x_10311 = v_3615 | ~v_60;
assign x_10312 = v_3615 | ~v_59;
assign x_10313 = v_3615 | ~v_51;
assign x_10314 = ~v_86 | ~v_157 | v_3614;
assign x_10315 = ~v_83 | ~v_156 | v_3613;
assign x_10316 = ~v_71 | v_157 | v_3612;
assign x_10317 = ~v_68 | v_156 | v_3611;
assign x_10318 = v_3610 | ~v_1572;
assign x_10319 = v_3610 | ~v_1573;
assign x_10320 = v_3610 | ~v_1574;
assign x_10321 = v_3610 | ~v_1575;
assign x_10322 = v_3610 | ~v_1804;
assign x_10323 = v_3610 | ~v_1805;
assign x_10324 = v_3610 | ~v_1806;
assign x_10325 = v_3610 | ~v_1807;
assign x_10326 = v_3610 | ~v_1576;
assign x_10327 = v_3610 | ~v_3460;
assign x_10328 = v_3610 | ~v_3461;
assign x_10329 = v_3610 | ~v_1579;
assign x_10330 = v_3610 | ~v_3462;
assign x_10331 = v_3610 | ~v_3463;
assign x_10332 = v_3610 | ~v_3606;
assign x_10333 = v_3610 | ~v_3607;
assign x_10334 = v_3610 | ~v_3608;
assign x_10335 = v_3610 | ~v_3609;
assign x_10336 = v_3610 | ~v_3464;
assign x_10337 = v_3610 | ~v_3465;
assign x_10338 = v_3610 | ~v_3466;
assign x_10339 = v_3610 | ~v_3469;
assign x_10340 = v_3610 | ~v_943;
assign x_10341 = v_3610 | ~v_944;
assign x_10342 = v_3610 | ~v_855;
assign x_10343 = v_3610 | ~v_856;
assign x_10344 = v_3610 | ~v_945;
assign x_10345 = v_3610 | ~v_946;
assign x_10346 = v_3610 | ~v_947;
assign x_10347 = v_3610 | ~v_948;
assign x_10348 = v_3610 | ~v_3471;
assign x_10349 = v_3610 | ~v_3472;
assign x_10350 = v_3610 | ~v_182;
assign x_10351 = v_3610 | ~v_179;
assign x_10352 = v_3610 | ~v_164;
assign x_10353 = v_3610 | ~v_163;
assign x_10354 = v_3610 | ~v_162;
assign x_10355 = v_3610 | ~v_137;
assign x_10356 = v_3610 | ~v_136;
assign x_10357 = v_3610 | ~v_135;
assign x_10358 = v_3610 | ~v_134;
assign x_10359 = v_3610 | ~v_17;
assign x_10360 = v_3610 | ~v_16;
assign x_10361 = v_3610 | ~v_8;
assign x_10362 = ~v_44 | ~v_157 | v_3609;
assign x_10363 = ~v_41 | ~v_156 | v_3608;
assign x_10364 = ~v_29 | v_157 | v_3607;
assign x_10365 = ~v_26 | v_156 | v_3606;
assign x_10366 = ~v_3604 | ~v_3603 | ~v_3602 | v_3605;
assign x_10367 = v_3604 | ~v_1718;
assign x_10368 = v_3604 | ~v_1719;
assign x_10369 = v_3604 | ~v_1720;
assign x_10370 = v_3604 | ~v_1721;
assign x_10371 = v_3604 | ~v_1626;
assign x_10372 = v_3604 | ~v_3490;
assign x_10373 = v_3604 | ~v_1627;
assign x_10374 = v_3604 | ~v_3491;
assign x_10375 = v_3604 | ~v_1628;
assign x_10376 = v_3604 | ~v_1629;
assign x_10377 = v_3604 | ~v_3492;
assign x_10378 = v_3604 | ~v_1630;
assign x_10379 = v_3604 | ~v_3493;
assign x_10380 = v_3604 | ~v_1631;
assign x_10381 = v_3604 | ~v_3548;
assign x_10382 = v_3604 | ~v_3549;
assign x_10383 = v_3604 | ~v_3550;
assign x_10384 = v_3604 | ~v_3551;
assign x_10385 = v_3604 | ~v_3496;
assign x_10386 = v_3604 | ~v_3497;
assign x_10387 = v_3604 | ~v_3498;
assign x_10388 = v_3604 | ~v_3499;
assign x_10389 = v_3604 | ~v_3500;
assign x_10390 = v_3604 | ~v_3501;
assign x_10391 = v_3604 | ~v_833;
assign x_10392 = v_3604 | ~v_834;
assign x_10393 = v_3604 | ~v_835;
assign x_10394 = v_3604 | ~v_836;
assign x_10395 = v_3604 | ~v_837;
assign x_10396 = v_3604 | ~v_838;
assign x_10397 = v_3604 | ~v_839;
assign x_10398 = v_3604 | ~v_840;
assign x_10399 = v_3604 | ~v_184;
assign x_10400 = v_3604 | ~v_169;
assign x_10401 = v_3604 | ~v_160;
assign x_10402 = v_3604 | ~v_150;
assign x_10403 = v_3604 | ~v_149;
assign x_10404 = v_3604 | ~v_147;
assign x_10405 = v_3604 | ~v_103;
assign x_10406 = v_3604 | ~v_102;
assign x_10407 = v_3604 | ~v_100;
assign x_10408 = v_3604 | ~v_98;
assign x_10409 = v_3604 | ~v_96;
assign x_10410 = v_3604 | ~v_94;
assign x_10411 = v_3603 | ~v_1709;
assign x_10412 = v_3603 | ~v_1710;
assign x_10413 = v_3603 | ~v_1711;
assign x_10414 = v_3603 | ~v_1712;
assign x_10415 = v_3603 | ~v_1601;
assign x_10416 = v_3603 | ~v_3475;
assign x_10417 = v_3603 | ~v_1602;
assign x_10418 = v_3603 | ~v_3476;
assign x_10419 = v_3603 | ~v_1603;
assign x_10420 = v_3603 | ~v_1604;
assign x_10421 = v_3603 | ~v_3477;
assign x_10422 = v_3603 | ~v_1605;
assign x_10423 = v_3603 | ~v_3478;
assign x_10424 = v_3603 | ~v_1606;
assign x_10425 = v_3603 | ~v_3543;
assign x_10426 = v_3603 | ~v_3544;
assign x_10427 = v_3603 | ~v_3545;
assign x_10428 = v_3603 | ~v_3546;
assign x_10429 = v_3603 | ~v_3481;
assign x_10430 = v_3603 | ~v_3482;
assign x_10431 = v_3603 | ~v_3483;
assign x_10432 = v_3603 | ~v_3484;
assign x_10433 = v_3603 | ~v_3485;
assign x_10434 = v_3603 | ~v_800;
assign x_10435 = v_3603 | ~v_801;
assign x_10436 = v_3603 | ~v_802;
assign x_10437 = v_3603 | ~v_803;
assign x_10438 = v_3603 | ~v_804;
assign x_10439 = v_3603 | ~v_805;
assign x_10440 = v_3603 | ~v_806;
assign x_10441 = v_3603 | ~v_807;
assign x_10442 = v_3603 | ~v_3486;
assign x_10443 = v_3603 | ~v_183;
assign x_10444 = v_3603 | ~v_165;
assign x_10445 = v_3603 | ~v_159;
assign x_10446 = v_3603 | ~v_145;
assign x_10447 = v_3603 | ~v_144;
assign x_10448 = v_3603 | ~v_142;
assign x_10449 = v_3603 | ~v_61;
assign x_10450 = v_3603 | ~v_60;
assign x_10451 = v_3603 | ~v_58;
assign x_10452 = v_3603 | ~v_56;
assign x_10453 = v_3603 | ~v_54;
assign x_10454 = v_3603 | ~v_52;
assign x_10455 = v_3602 | ~v_1700;
assign x_10456 = v_3602 | ~v_1701;
assign x_10457 = v_3602 | ~v_1702;
assign x_10458 = v_3602 | ~v_1703;
assign x_10459 = v_3602 | ~v_1576;
assign x_10460 = v_3602 | ~v_3460;
assign x_10461 = v_3602 | ~v_1577;
assign x_10462 = v_3602 | ~v_3461;
assign x_10463 = v_3602 | ~v_1578;
assign x_10464 = v_3602 | ~v_1579;
assign x_10465 = v_3602 | ~v_3462;
assign x_10466 = v_3602 | ~v_1580;
assign x_10467 = v_3602 | ~v_3463;
assign x_10468 = v_3602 | ~v_1581;
assign x_10469 = v_3602 | ~v_3538;
assign x_10470 = v_3602 | ~v_3539;
assign x_10471 = v_3602 | ~v_3540;
assign x_10472 = v_3602 | ~v_3541;
assign x_10473 = v_3602 | ~v_3466;
assign x_10474 = v_3602 | ~v_3467;
assign x_10475 = v_3602 | ~v_3468;
assign x_10476 = v_3602 | ~v_3469;
assign x_10477 = v_3602 | ~v_3470;
assign x_10478 = v_3602 | ~v_767;
assign x_10479 = v_3602 | ~v_768;
assign x_10480 = v_3602 | ~v_769;
assign x_10481 = v_3602 | ~v_770;
assign x_10482 = v_3602 | ~v_771;
assign x_10483 = v_3602 | ~v_772;
assign x_10484 = v_3602 | ~v_773;
assign x_10485 = v_3602 | ~v_774;
assign x_10486 = v_3602 | ~v_182;
assign x_10487 = v_3602 | ~v_161;
assign x_10488 = v_3602 | ~v_155;
assign x_10489 = v_3602 | ~v_137;
assign x_10490 = v_3602 | ~v_3473;
assign x_10491 = v_3602 | ~v_136;
assign x_10492 = v_3602 | ~v_134;
assign x_10493 = v_3602 | ~v_18;
assign x_10494 = v_3602 | ~v_17;
assign x_10495 = v_3602 | ~v_15;
assign x_10496 = v_3602 | ~v_13;
assign x_10497 = v_3602 | ~v_11;
assign x_10498 = v_3602 | ~v_9;
assign x_10499 = ~v_3600 | ~v_3599 | ~v_3598 | v_3601;
assign x_10500 = v_3600 | ~v_1778;
assign x_10501 = v_3600 | ~v_1779;
assign x_10502 = v_3600 | ~v_1780;
assign x_10503 = v_3600 | ~v_1781;
assign x_10504 = v_3600 | ~v_1626;
assign x_10505 = v_3600 | ~v_3490;
assign x_10506 = v_3600 | ~v_1746;
assign x_10507 = v_3600 | ~v_3491;
assign x_10508 = v_3600 | ~v_1747;
assign x_10509 = v_3600 | ~v_1629;
assign x_10510 = v_3600 | ~v_3492;
assign x_10511 = v_3600 | ~v_1748;
assign x_10512 = v_3600 | ~v_3493;
assign x_10513 = v_3600 | ~v_1749;
assign x_10514 = v_3600 | ~v_3584;
assign x_10515 = v_3600 | ~v_3585;
assign x_10516 = v_3600 | ~v_3586;
assign x_10517 = v_3600 | ~v_3587;
assign x_10518 = v_3600 | ~v_3496;
assign x_10519 = v_3600 | ~v_3564;
assign x_10520 = v_3600 | ~v_3565;
assign x_10521 = v_3600 | ~v_3499;
assign x_10522 = v_3600 | ~v_3566;
assign x_10523 = v_3600 | ~v_3567;
assign x_10524 = v_3600 | ~v_1085;
assign x_10525 = v_3600 | ~v_1131;
assign x_10526 = v_3600 | ~v_1132;
assign x_10527 = v_3600 | ~v_1086;
assign x_10528 = v_3600 | ~v_1133;
assign x_10529 = v_3600 | ~v_1134;
assign x_10530 = v_3600 | ~v_1023;
assign x_10531 = v_3600 | ~v_1024;
assign x_10532 = v_3600 | ~v_184;
assign x_10533 = v_3600 | ~v_172;
assign x_10534 = v_3600 | ~v_171;
assign x_10535 = v_3600 | ~v_170;
assign x_10536 = v_3600 | ~v_169;
assign x_10537 = v_3600 | ~v_148;
assign x_10538 = v_3600 | ~v_147;
assign x_10539 = v_3600 | ~v_102;
assign x_10540 = v_3600 | ~v_101;
assign x_10541 = v_3600 | ~v_100;
assign x_10542 = v_3600 | ~v_99;
assign x_10543 = v_3600 | ~v_97;
assign x_10544 = v_3599 | ~v_1769;
assign x_10545 = v_3599 | ~v_1770;
assign x_10546 = v_3599 | ~v_1771;
assign x_10547 = v_3599 | ~v_1772;
assign x_10548 = v_3599 | ~v_1601;
assign x_10549 = v_3599 | ~v_3475;
assign x_10550 = v_3599 | ~v_1737;
assign x_10551 = v_3599 | ~v_3476;
assign x_10552 = v_3599 | ~v_1738;
assign x_10553 = v_3599 | ~v_1604;
assign x_10554 = v_3599 | ~v_3477;
assign x_10555 = v_3599 | ~v_1739;
assign x_10556 = v_3599 | ~v_3478;
assign x_10557 = v_3599 | ~v_1740;
assign x_10558 = v_3599 | ~v_3579;
assign x_10559 = v_3599 | ~v_3580;
assign x_10560 = v_3599 | ~v_3581;
assign x_10561 = v_3599 | ~v_3582;
assign x_10562 = v_3599 | ~v_3481;
assign x_10563 = v_3599 | ~v_3559;
assign x_10564 = v_3599 | ~v_3560;
assign x_10565 = v_3599 | ~v_3484;
assign x_10566 = v_3599 | ~v_1070;
assign x_10567 = v_3599 | ~v_1126;
assign x_10568 = v_3599 | ~v_1127;
assign x_10569 = v_3599 | ~v_1071;
assign x_10570 = v_3599 | ~v_1128;
assign x_10571 = v_3599 | ~v_1129;
assign x_10572 = v_3599 | ~v_1008;
assign x_10573 = v_3599 | ~v_1009;
assign x_10574 = v_3599 | ~v_3561;
assign x_10575 = v_3599 | ~v_3562;
assign x_10576 = v_3599 | ~v_183;
assign x_10577 = v_3599 | ~v_168;
assign x_10578 = v_3599 | ~v_167;
assign x_10579 = v_3599 | ~v_166;
assign x_10580 = v_3599 | ~v_165;
assign x_10581 = v_3599 | ~v_143;
assign x_10582 = v_3599 | ~v_142;
assign x_10583 = v_3599 | ~v_60;
assign x_10584 = v_3599 | ~v_59;
assign x_10585 = v_3599 | ~v_58;
assign x_10586 = v_3599 | ~v_57;
assign x_10587 = v_3599 | ~v_55;
assign x_10588 = v_3598 | ~v_1760;
assign x_10589 = v_3598 | ~v_1761;
assign x_10590 = v_3598 | ~v_1762;
assign x_10591 = v_3598 | ~v_1763;
assign x_10592 = v_3598 | ~v_1576;
assign x_10593 = v_3598 | ~v_3460;
assign x_10594 = v_3598 | ~v_1728;
assign x_10595 = v_3598 | ~v_3461;
assign x_10596 = v_3598 | ~v_1729;
assign x_10597 = v_3598 | ~v_1579;
assign x_10598 = v_3598 | ~v_3462;
assign x_10599 = v_3598 | ~v_1730;
assign x_10600 = v_3598 | ~v_3463;
assign x_10601 = v_3598 | ~v_1731;
assign x_10602 = v_3598 | ~v_3574;
assign x_10603 = v_3598 | ~v_3575;
assign x_10604 = v_3598 | ~v_3576;
assign x_10605 = v_3598 | ~v_3577;
assign x_10606 = v_3598 | ~v_3466;
assign x_10607 = v_3598 | ~v_3554;
assign x_10608 = v_3598 | ~v_3555;
assign x_10609 = v_3598 | ~v_3469;
assign x_10610 = v_3598 | ~v_3556;
assign x_10611 = v_3598 | ~v_3557;
assign x_10612 = v_3598 | ~v_1055;
assign x_10613 = v_3598 | ~v_1121;
assign x_10614 = v_3598 | ~v_1122;
assign x_10615 = v_3598 | ~v_1056;
assign x_10616 = v_3598 | ~v_1123;
assign x_10617 = v_3598 | ~v_1124;
assign x_10618 = v_3598 | ~v_182;
assign x_10619 = v_3598 | ~v_164;
assign x_10620 = v_3598 | ~v_163;
assign x_10621 = v_3598 | ~v_162;
assign x_10622 = v_3598 | ~v_161;
assign x_10623 = v_3598 | ~v_135;
assign x_10624 = v_3598 | ~v_134;
assign x_10625 = v_3598 | ~v_993;
assign x_10626 = v_3598 | ~v_994;
assign x_10627 = v_3598 | ~v_17;
assign x_10628 = v_3598 | ~v_16;
assign x_10629 = v_3598 | ~v_15;
assign x_10630 = v_3598 | ~v_14;
assign x_10631 = v_3598 | ~v_12;
assign x_10632 = ~v_3596 | ~v_3595 | ~v_3594 | v_3597;
assign x_10633 = v_3596 | ~v_1778;
assign x_10634 = v_3596 | ~v_1779;
assign x_10635 = v_3596 | ~v_1780;
assign x_10636 = v_3596 | ~v_1781;
assign x_10637 = v_3596 | ~v_1718;
assign x_10638 = v_3596 | ~v_1719;
assign x_10639 = v_3596 | ~v_1720;
assign x_10640 = v_3596 | ~v_1721;
assign x_10641 = v_3596 | ~v_1626;
assign x_10642 = v_3596 | ~v_3490;
assign x_10643 = v_3596 | ~v_3491;
assign x_10644 = v_3596 | ~v_1629;
assign x_10645 = v_3596 | ~v_3492;
assign x_10646 = v_3596 | ~v_3493;
assign x_10647 = v_3596 | ~v_3548;
assign x_10648 = v_3596 | ~v_3549;
assign x_10649 = v_3596 | ~v_3550;
assign x_10650 = v_3596 | ~v_3551;
assign x_10651 = v_3596 | ~v_3584;
assign x_10652 = v_3596 | ~v_3585;
assign x_10653 = v_3596 | ~v_3586;
assign x_10654 = v_3596 | ~v_3587;
assign x_10655 = v_3596 | ~v_3496;
assign x_10656 = v_3596 | ~v_3499;
assign x_10657 = v_3596 | ~v_837;
assign x_10658 = v_3596 | ~v_838;
assign x_10659 = v_3596 | ~v_1081;
assign x_10660 = v_3596 | ~v_1082;
assign x_10661 = v_3596 | ~v_1083;
assign x_10662 = v_3596 | ~v_1084;
assign x_10663 = v_3596 | ~v_1085;
assign x_10664 = v_3596 | ~v_1086;
assign x_10665 = v_3596 | ~v_184;
assign x_10666 = v_3596 | ~v_171;
assign x_10667 = v_3596 | ~v_170;
assign x_10668 = v_3596 | ~v_169;
assign x_10669 = v_3596 | ~v_160;
assign x_10670 = v_3596 | ~v_150;
assign x_10671 = v_3596 | ~v_149;
assign x_10672 = v_3596 | ~v_147;
assign x_10673 = v_3596 | ~v_103;
assign x_10674 = v_3596 | ~v_102;
assign x_10675 = v_3596 | ~v_100;
assign x_10676 = v_3596 | ~v_96;
assign x_10677 = v_3595 | ~v_1769;
assign x_10678 = v_3595 | ~v_1770;
assign x_10679 = v_3595 | ~v_1771;
assign x_10680 = v_3595 | ~v_1772;
assign x_10681 = v_3595 | ~v_1709;
assign x_10682 = v_3595 | ~v_1710;
assign x_10683 = v_3595 | ~v_1711;
assign x_10684 = v_3595 | ~v_1712;
assign x_10685 = v_3595 | ~v_1601;
assign x_10686 = v_3595 | ~v_3475;
assign x_10687 = v_3595 | ~v_3476;
assign x_10688 = v_3595 | ~v_1604;
assign x_10689 = v_3595 | ~v_3477;
assign x_10690 = v_3595 | ~v_3478;
assign x_10691 = v_3595 | ~v_3543;
assign x_10692 = v_3595 | ~v_3544;
assign x_10693 = v_3595 | ~v_3545;
assign x_10694 = v_3595 | ~v_3546;
assign x_10695 = v_3595 | ~v_3579;
assign x_10696 = v_3595 | ~v_3580;
assign x_10697 = v_3595 | ~v_3581;
assign x_10698 = v_3595 | ~v_3582;
assign x_10699 = v_3595 | ~v_3481;
assign x_10700 = v_3595 | ~v_3484;
assign x_10701 = v_3595 | ~v_804;
assign x_10702 = v_3595 | ~v_805;
assign x_10703 = v_3595 | ~v_1066;
assign x_10704 = v_3595 | ~v_1067;
assign x_10705 = v_3595 | ~v_1068;
assign x_10706 = v_3595 | ~v_1069;
assign x_10707 = v_3595 | ~v_1070;
assign x_10708 = v_3595 | ~v_1071;
assign x_10709 = v_3595 | ~v_183;
assign x_10710 = v_3595 | ~v_167;
assign x_10711 = v_3595 | ~v_166;
assign x_10712 = v_3595 | ~v_165;
assign x_10713 = v_3595 | ~v_159;
assign x_10714 = v_3595 | ~v_145;
assign x_10715 = v_3595 | ~v_144;
assign x_10716 = v_3595 | ~v_142;
assign x_10717 = v_3595 | ~v_61;
assign x_10718 = v_3595 | ~v_60;
assign x_10719 = v_3595 | ~v_58;
assign x_10720 = v_3595 | ~v_54;
assign x_10721 = v_3594 | ~v_1760;
assign x_10722 = v_3594 | ~v_1761;
assign x_10723 = v_3594 | ~v_1762;
assign x_10724 = v_3594 | ~v_1763;
assign x_10725 = v_3594 | ~v_1700;
assign x_10726 = v_3594 | ~v_1701;
assign x_10727 = v_3594 | ~v_1702;
assign x_10728 = v_3594 | ~v_1703;
assign x_10729 = v_3594 | ~v_1576;
assign x_10730 = v_3594 | ~v_3460;
assign x_10731 = v_3594 | ~v_3461;
assign x_10732 = v_3594 | ~v_1579;
assign x_10733 = v_3594 | ~v_3462;
assign x_10734 = v_3594 | ~v_3463;
assign x_10735 = v_3594 | ~v_3538;
assign x_10736 = v_3594 | ~v_3539;
assign x_10737 = v_3594 | ~v_3540;
assign x_10738 = v_3594 | ~v_3541;
assign x_10739 = v_3594 | ~v_3574;
assign x_10740 = v_3594 | ~v_3575;
assign x_10741 = v_3594 | ~v_3576;
assign x_10742 = v_3594 | ~v_3577;
assign x_10743 = v_3594 | ~v_3466;
assign x_10744 = v_3594 | ~v_3469;
assign x_10745 = v_3594 | ~v_771;
assign x_10746 = v_3594 | ~v_772;
assign x_10747 = v_3594 | ~v_1051;
assign x_10748 = v_3594 | ~v_1052;
assign x_10749 = v_3594 | ~v_1053;
assign x_10750 = v_3594 | ~v_1054;
assign x_10751 = v_3594 | ~v_1055;
assign x_10752 = v_3594 | ~v_1056;
assign x_10753 = v_3594 | ~v_182;
assign x_10754 = v_3594 | ~v_163;
assign x_10755 = v_3594 | ~v_162;
assign x_10756 = v_3594 | ~v_161;
assign x_10757 = v_3594 | ~v_155;
assign x_10758 = v_3594 | ~v_137;
assign x_10759 = v_3594 | ~v_136;
assign x_10760 = v_3594 | ~v_134;
assign x_10761 = v_3594 | ~v_18;
assign x_10762 = v_3594 | ~v_17;
assign x_10763 = v_3594 | ~v_15;
assign x_10764 = v_3594 | ~v_11;
assign x_10765 = ~v_3592 | ~v_3591 | ~v_3590 | v_3593;
assign x_10766 = v_3592 | ~v_1778;
assign x_10767 = v_3592 | ~v_1779;
assign x_10768 = v_3592 | ~v_1780;
assign x_10769 = v_3592 | ~v_1781;
assign x_10770 = v_3592 | ~v_1690;
assign x_10771 = v_3592 | ~v_1691;
assign x_10772 = v_3592 | ~v_1692;
assign x_10773 = v_3592 | ~v_1693;
assign x_10774 = v_3592 | ~v_1626;
assign x_10775 = v_3592 | ~v_3490;
assign x_10776 = v_3592 | ~v_3491;
assign x_10777 = v_3592 | ~v_1629;
assign x_10778 = v_3592 | ~v_3492;
assign x_10779 = v_3592 | ~v_3493;
assign x_10780 = v_3592 | ~v_3532;
assign x_10781 = v_3592 | ~v_3533;
assign x_10782 = v_3592 | ~v_3534;
assign x_10783 = v_3592 | ~v_3535;
assign x_10784 = v_3592 | ~v_3584;
assign x_10785 = v_3592 | ~v_3585;
assign x_10786 = v_3592 | ~v_3586;
assign x_10787 = v_3592 | ~v_3587;
assign x_10788 = v_3592 | ~v_3496;
assign x_10789 = v_3592 | ~v_3499;
assign x_10790 = v_3592 | ~v_927;
assign x_10791 = v_3592 | ~v_928;
assign x_10792 = v_3592 | ~v_1099;
assign x_10793 = v_3592 | ~v_1100;
assign x_10794 = v_3592 | ~v_1101;
assign x_10795 = v_3592 | ~v_1102;
assign x_10796 = v_3592 | ~v_1085;
assign x_10797 = v_3592 | ~v_1086;
assign x_10798 = v_3592 | ~v_184;
assign x_10799 = v_3592 | ~v_171;
assign x_10800 = v_3592 | ~v_170;
assign x_10801 = v_3592 | ~v_169;
assign x_10802 = v_3592 | ~v_150;
assign x_10803 = v_3592 | ~v_149;
assign x_10804 = v_3592 | ~v_148;
assign x_10805 = v_3592 | ~v_103;
assign x_10806 = v_3592 | ~v_102;
assign x_10807 = v_3592 | ~v_101;
assign x_10808 = v_3592 | ~v_100;
assign x_10809 = v_3592 | ~v_95;
assign x_10810 = v_3591 | ~v_1769;
assign x_10811 = v_3591 | ~v_1770;
assign x_10812 = v_3591 | ~v_1771;
assign x_10813 = v_3591 | ~v_1772;
assign x_10814 = v_3591 | ~v_1681;
assign x_10815 = v_3591 | ~v_1682;
assign x_10816 = v_3591 | ~v_1683;
assign x_10817 = v_3591 | ~v_1684;
assign x_10818 = v_3591 | ~v_1601;
assign x_10819 = v_3591 | ~v_3475;
assign x_10820 = v_3591 | ~v_3476;
assign x_10821 = v_3591 | ~v_1604;
assign x_10822 = v_3591 | ~v_3477;
assign x_10823 = v_3591 | ~v_3478;
assign x_10824 = v_3591 | ~v_3527;
assign x_10825 = v_3591 | ~v_3528;
assign x_10826 = v_3591 | ~v_3529;
assign x_10827 = v_3591 | ~v_3530;
assign x_10828 = v_3591 | ~v_3579;
assign x_10829 = v_3591 | ~v_3580;
assign x_10830 = v_3591 | ~v_3581;
assign x_10831 = v_3591 | ~v_3582;
assign x_10832 = v_3591 | ~v_3481;
assign x_10833 = v_3591 | ~v_3484;
assign x_10834 = v_3591 | ~v_912;
assign x_10835 = v_3591 | ~v_913;
assign x_10836 = v_3591 | ~v_1094;
assign x_10837 = v_3591 | ~v_1095;
assign x_10838 = v_3591 | ~v_1096;
assign x_10839 = v_3591 | ~v_1097;
assign x_10840 = v_3591 | ~v_1070;
assign x_10841 = v_3591 | ~v_1071;
assign x_10842 = v_3591 | ~v_183;
assign x_10843 = v_3591 | ~v_167;
assign x_10844 = v_3591 | ~v_166;
assign x_10845 = v_3591 | ~v_165;
assign x_10846 = v_3591 | ~v_145;
assign x_10847 = v_3591 | ~v_144;
assign x_10848 = v_3591 | ~v_143;
assign x_10849 = v_3591 | ~v_61;
assign x_10850 = v_3591 | ~v_60;
assign x_10851 = v_3591 | ~v_59;
assign x_10852 = v_3591 | ~v_58;
assign x_10853 = v_3591 | ~v_53;
assign x_10854 = v_3590 | ~v_1760;
assign x_10855 = v_3590 | ~v_1761;
assign x_10856 = v_3590 | ~v_1762;
assign x_10857 = v_3590 | ~v_1763;
assign x_10858 = v_3590 | ~v_1672;
assign x_10859 = v_3590 | ~v_1673;
assign x_10860 = v_3590 | ~v_1674;
assign x_10861 = v_3590 | ~v_1675;
assign x_10862 = v_3590 | ~v_1576;
assign x_10863 = v_3590 | ~v_3460;
assign x_10864 = v_3590 | ~v_3461;
assign x_10865 = v_3590 | ~v_1579;
assign x_10866 = v_3590 | ~v_3462;
assign x_10867 = v_3590 | ~v_3463;
assign x_10868 = v_3590 | ~v_3522;
assign x_10869 = v_3590 | ~v_3523;
assign x_10870 = v_3590 | ~v_3524;
assign x_10871 = v_3590 | ~v_3525;
assign x_10872 = v_3590 | ~v_3574;
assign x_10873 = v_3590 | ~v_3575;
assign x_10874 = v_3590 | ~v_3576;
assign x_10875 = v_3590 | ~v_3577;
assign x_10876 = v_3590 | ~v_3466;
assign x_10877 = v_3590 | ~v_3469;
assign x_10878 = v_3590 | ~v_897;
assign x_10879 = v_3590 | ~v_898;
assign x_10880 = v_3590 | ~v_1089;
assign x_10881 = v_3590 | ~v_1090;
assign x_10882 = v_3590 | ~v_1091;
assign x_10883 = v_3590 | ~v_1092;
assign x_10884 = v_3590 | ~v_1055;
assign x_10885 = v_3590 | ~v_1056;
assign x_10886 = v_3590 | ~v_182;
assign x_10887 = v_3590 | ~v_163;
assign x_10888 = v_3590 | ~v_162;
assign x_10889 = v_3590 | ~v_161;
assign x_10890 = v_3590 | ~v_137;
assign x_10891 = v_3590 | ~v_136;
assign x_10892 = v_3590 | ~v_135;
assign x_10893 = v_3590 | ~v_18;
assign x_10894 = v_3590 | ~v_17;
assign x_10895 = v_3590 | ~v_16;
assign x_10896 = v_3590 | ~v_15;
assign x_10897 = v_3590 | ~v_10;
assign x_10898 = ~v_3588 | ~v_3583 | ~v_3578 | v_3589;
assign x_10899 = v_3588 | ~v_1778;
assign x_10900 = v_3588 | ~v_1779;
assign x_10901 = v_3588 | ~v_1780;
assign x_10902 = v_3588 | ~v_1781;
assign x_10903 = v_3588 | ~v_1622;
assign x_10904 = v_3588 | ~v_1623;
assign x_10905 = v_3588 | ~v_1624;
assign x_10906 = v_3588 | ~v_1625;
assign x_10907 = v_3588 | ~v_1626;
assign x_10908 = v_3588 | ~v_3490;
assign x_10909 = v_3588 | ~v_3491;
assign x_10910 = v_3588 | ~v_1629;
assign x_10911 = v_3588 | ~v_3492;
assign x_10912 = v_3588 | ~v_3493;
assign x_10913 = v_3588 | ~v_3494;
assign x_10914 = v_3588 | ~v_3495;
assign x_10915 = v_3588 | ~v_3584;
assign x_10916 = v_3588 | ~v_3585;
assign x_10917 = v_3588 | ~v_3586;
assign x_10918 = v_3588 | ~v_3587;
assign x_10919 = v_3588 | ~v_3496;
assign x_10920 = v_3588 | ~v_3499;
assign x_10921 = v_3588 | ~v_975;
assign x_10922 = v_3588 | ~v_976;
assign x_10923 = v_3588 | ~v_1115;
assign x_10924 = v_3588 | ~v_1116;
assign x_10925 = v_3588 | ~v_1085;
assign x_10926 = v_3588 | ~v_1086;
assign x_10927 = v_3588 | ~v_1117;
assign x_10928 = v_3588 | ~v_1118;
assign x_10929 = v_3588 | ~v_3502;
assign x_10930 = v_3588 | ~v_3503;
assign x_10931 = v_3588 | ~v_184;
assign x_10932 = v_3588 | ~v_171;
assign x_10933 = v_3588 | ~v_170;
assign x_10934 = v_3588 | ~v_169;
assign x_10935 = v_3588 | ~v_151;
assign x_10936 = v_3588 | ~v_150;
assign x_10937 = v_3588 | ~v_149;
assign x_10938 = v_3588 | ~v_148;
assign x_10939 = v_3588 | ~v_147;
assign x_10940 = v_3588 | ~v_103;
assign x_10941 = v_3588 | ~v_101;
assign x_10942 = v_3588 | ~v_100;
assign x_10943 = ~v_128 | ~v_140 | v_3587;
assign x_10944 = ~v_125 | ~v_139 | v_3586;
assign x_10945 = ~v_113 | v_140 | v_3585;
assign x_10946 = ~v_110 | v_139 | v_3584;
assign x_10947 = v_3583 | ~v_1769;
assign x_10948 = v_3583 | ~v_1770;
assign x_10949 = v_3583 | ~v_1771;
assign x_10950 = v_3583 | ~v_1772;
assign x_10951 = v_3583 | ~v_1597;
assign x_10952 = v_3583 | ~v_1598;
assign x_10953 = v_3583 | ~v_1599;
assign x_10954 = v_3583 | ~v_1600;
assign x_10955 = v_3583 | ~v_1601;
assign x_10956 = v_3583 | ~v_3475;
assign x_10957 = v_3583 | ~v_3476;
assign x_10958 = v_3583 | ~v_1604;
assign x_10959 = v_3583 | ~v_3477;
assign x_10960 = v_3583 | ~v_3478;
assign x_10961 = v_3583 | ~v_3479;
assign x_10962 = v_3583 | ~v_3480;
assign x_10963 = v_3583 | ~v_3579;
assign x_10964 = v_3583 | ~v_3580;
assign x_10965 = v_3583 | ~v_3581;
assign x_10966 = v_3583 | ~v_3582;
assign x_10967 = v_3583 | ~v_3481;
assign x_10968 = v_3583 | ~v_3484;
assign x_10969 = v_3583 | ~v_960;
assign x_10970 = v_3583 | ~v_961;
assign x_10971 = v_3583 | ~v_1110;
assign x_10972 = v_3583 | ~v_1111;
assign x_10973 = v_3583 | ~v_1070;
assign x_10974 = v_3583 | ~v_1071;
assign x_10975 = v_3583 | ~v_1112;
assign x_10976 = v_3583 | ~v_1113;
assign x_10977 = v_3583 | ~v_3487;
assign x_10978 = v_3583 | ~v_3488;
assign x_10979 = v_3583 | ~v_183;
assign x_10980 = v_3583 | ~v_167;
assign x_10981 = v_3583 | ~v_166;
assign x_10982 = v_3583 | ~v_165;
assign x_10983 = v_3583 | ~v_146;
assign x_10984 = v_3583 | ~v_145;
assign x_10985 = v_3583 | ~v_144;
assign x_10986 = v_3583 | ~v_143;
assign x_10987 = v_3583 | ~v_142;
assign x_10988 = v_3583 | ~v_61;
assign x_10989 = v_3583 | ~v_59;
assign x_10990 = v_3583 | ~v_58;
assign x_10991 = ~v_86 | ~v_140 | v_3582;
assign x_10992 = ~v_83 | ~v_139 | v_3581;
assign x_10993 = ~v_71 | v_140 | v_3580;
assign x_10994 = ~v_68 | v_139 | v_3579;
assign x_10995 = v_3578 | ~v_1760;
assign x_10996 = v_3578 | ~v_1761;
assign x_10997 = v_3578 | ~v_1762;
assign x_10998 = v_3578 | ~v_1763;
assign x_10999 = v_3578 | ~v_1572;
assign x_11000 = v_3578 | ~v_1573;
assign x_11001 = v_3578 | ~v_1574;
assign x_11002 = v_3578 | ~v_1575;
assign x_11003 = v_3578 | ~v_1576;
assign x_11004 = v_3578 | ~v_3460;
assign x_11005 = v_3578 | ~v_3461;
assign x_11006 = v_3578 | ~v_1579;
assign x_11007 = v_3578 | ~v_3462;
assign x_11008 = v_3578 | ~v_3463;
assign x_11009 = v_3578 | ~v_3464;
assign x_11010 = v_3578 | ~v_3465;
assign x_11011 = v_3578 | ~v_3574;
assign x_11012 = v_3578 | ~v_3575;
assign x_11013 = v_3578 | ~v_3576;
assign x_11014 = v_3578 | ~v_3577;
assign x_11015 = v_3578 | ~v_3466;
assign x_11016 = v_3578 | ~v_3469;
assign x_11017 = v_3578 | ~v_945;
assign x_11018 = v_3578 | ~v_946;
assign x_11019 = v_3578 | ~v_1105;
assign x_11020 = v_3578 | ~v_1106;
assign x_11021 = v_3578 | ~v_1055;
assign x_11022 = v_3578 | ~v_1056;
assign x_11023 = v_3578 | ~v_1107;
assign x_11024 = v_3578 | ~v_1108;
assign x_11025 = v_3578 | ~v_3471;
assign x_11026 = v_3578 | ~v_3472;
assign x_11027 = v_3578 | ~v_182;
assign x_11028 = v_3578 | ~v_163;
assign x_11029 = v_3578 | ~v_162;
assign x_11030 = v_3578 | ~v_161;
assign x_11031 = v_3578 | ~v_138;
assign x_11032 = v_3578 | ~v_137;
assign x_11033 = v_3578 | ~v_136;
assign x_11034 = v_3578 | ~v_135;
assign x_11035 = v_3578 | ~v_134;
assign x_11036 = v_3578 | ~v_18;
assign x_11037 = v_3578 | ~v_16;
assign x_11038 = v_3578 | ~v_15;
assign x_11039 = ~v_44 | ~v_140 | v_3577;
assign x_11040 = ~v_41 | ~v_139 | v_3576;
assign x_11041 = ~v_29 | v_140 | v_3575;
assign x_11042 = ~v_26 | v_139 | v_3574;
assign x_11043 = ~v_3572 | ~v_3571 | ~v_3570 | v_3573;
assign x_11044 = v_3572 | ~v_1690;
assign x_11045 = v_3572 | ~v_1691;
assign x_11046 = v_3572 | ~v_1692;
assign x_11047 = v_3572 | ~v_1693;
assign x_11048 = v_3572 | ~v_1626;
assign x_11049 = v_3572 | ~v_3490;
assign x_11050 = v_3572 | ~v_1627;
assign x_11051 = v_3572 | ~v_3491;
assign x_11052 = v_3572 | ~v_1628;
assign x_11053 = v_3572 | ~v_1629;
assign x_11054 = v_3572 | ~v_3492;
assign x_11055 = v_3572 | ~v_1630;
assign x_11056 = v_3572 | ~v_3493;
assign x_11057 = v_3572 | ~v_1631;
assign x_11058 = v_3572 | ~v_3532;
assign x_11059 = v_3572 | ~v_3533;
assign x_11060 = v_3572 | ~v_3534;
assign x_11061 = v_3572 | ~v_3535;
assign x_11062 = v_3572 | ~v_3496;
assign x_11063 = v_3572 | ~v_3497;
assign x_11064 = v_3572 | ~v_3498;
assign x_11065 = v_3572 | ~v_3499;
assign x_11066 = v_3572 | ~v_3500;
assign x_11067 = v_3572 | ~v_3501;
assign x_11068 = v_3572 | ~v_1037;
assign x_11069 = v_3572 | ~v_1038;
assign x_11070 = v_3572 | ~v_1039;
assign x_11071 = v_3572 | ~v_1040;
assign x_11072 = v_3572 | ~v_927;
assign x_11073 = v_3572 | ~v_928;
assign x_11074 = v_3572 | ~v_839;
assign x_11075 = v_3572 | ~v_840;
assign x_11076 = v_3572 | ~v_184;
assign x_11077 = v_3572 | ~v_169;
assign x_11078 = v_3572 | ~v_151;
assign x_11079 = v_3572 | ~v_150;
assign x_11080 = v_3572 | ~v_149;
assign x_11081 = v_3572 | ~v_148;
assign x_11082 = v_3572 | ~v_147;
assign x_11083 = v_3572 | ~v_103;
assign x_11084 = v_3572 | ~v_101;
assign x_11085 = v_3572 | ~v_100;
assign x_11086 = v_3572 | ~v_98;
assign x_11087 = v_3572 | ~v_94;
assign x_11088 = v_3571 | ~v_1681;
assign x_11089 = v_3571 | ~v_1682;
assign x_11090 = v_3571 | ~v_1683;
assign x_11091 = v_3571 | ~v_1684;
assign x_11092 = v_3571 | ~v_1601;
assign x_11093 = v_3571 | ~v_3475;
assign x_11094 = v_3571 | ~v_1602;
assign x_11095 = v_3571 | ~v_3476;
assign x_11096 = v_3571 | ~v_1603;
assign x_11097 = v_3571 | ~v_1604;
assign x_11098 = v_3571 | ~v_3477;
assign x_11099 = v_3571 | ~v_1605;
assign x_11100 = v_3571 | ~v_3478;
assign x_11101 = v_3571 | ~v_1606;
assign x_11102 = v_3571 | ~v_3527;
assign x_11103 = v_3571 | ~v_3528;
assign x_11104 = v_3571 | ~v_3529;
assign x_11105 = v_3571 | ~v_3530;
assign x_11106 = v_3571 | ~v_3481;
assign x_11107 = v_3571 | ~v_3482;
assign x_11108 = v_3571 | ~v_3483;
assign x_11109 = v_3571 | ~v_3484;
assign x_11110 = v_3571 | ~v_3485;
assign x_11111 = v_3571 | ~v_1032;
assign x_11112 = v_3571 | ~v_1033;
assign x_11113 = v_3571 | ~v_1034;
assign x_11114 = v_3571 | ~v_1035;
assign x_11115 = v_3571 | ~v_912;
assign x_11116 = v_3571 | ~v_913;
assign x_11117 = v_3571 | ~v_806;
assign x_11118 = v_3571 | ~v_807;
assign x_11119 = v_3571 | ~v_3486;
assign x_11120 = v_3571 | ~v_183;
assign x_11121 = v_3571 | ~v_165;
assign x_11122 = v_3571 | ~v_146;
assign x_11123 = v_3571 | ~v_145;
assign x_11124 = v_3571 | ~v_144;
assign x_11125 = v_3571 | ~v_143;
assign x_11126 = v_3571 | ~v_142;
assign x_11127 = v_3571 | ~v_61;
assign x_11128 = v_3571 | ~v_59;
assign x_11129 = v_3571 | ~v_58;
assign x_11130 = v_3571 | ~v_56;
assign x_11131 = v_3571 | ~v_52;
assign x_11132 = v_3570 | ~v_1672;
assign x_11133 = v_3570 | ~v_1673;
assign x_11134 = v_3570 | ~v_1674;
assign x_11135 = v_3570 | ~v_1675;
assign x_11136 = v_3570 | ~v_1576;
assign x_11137 = v_3570 | ~v_3460;
assign x_11138 = v_3570 | ~v_1577;
assign x_11139 = v_3570 | ~v_3461;
assign x_11140 = v_3570 | ~v_1578;
assign x_11141 = v_3570 | ~v_1579;
assign x_11142 = v_3570 | ~v_3462;
assign x_11143 = v_3570 | ~v_1580;
assign x_11144 = v_3570 | ~v_3463;
assign x_11145 = v_3570 | ~v_1581;
assign x_11146 = v_3570 | ~v_3522;
assign x_11147 = v_3570 | ~v_3523;
assign x_11148 = v_3570 | ~v_3524;
assign x_11149 = v_3570 | ~v_3525;
assign x_11150 = v_3570 | ~v_3466;
assign x_11151 = v_3570 | ~v_3467;
assign x_11152 = v_3570 | ~v_3468;
assign x_11153 = v_3570 | ~v_3469;
assign x_11154 = v_3570 | ~v_3470;
assign x_11155 = v_3570 | ~v_1027;
assign x_11156 = v_3570 | ~v_1028;
assign x_11157 = v_3570 | ~v_1029;
assign x_11158 = v_3570 | ~v_1030;
assign x_11159 = v_3570 | ~v_897;
assign x_11160 = v_3570 | ~v_898;
assign x_11161 = v_3570 | ~v_773;
assign x_11162 = v_3570 | ~v_774;
assign x_11163 = v_3570 | ~v_182;
assign x_11164 = v_3570 | ~v_161;
assign x_11165 = v_3570 | ~v_138;
assign x_11166 = v_3570 | ~v_137;
assign x_11167 = v_3570 | ~v_3473;
assign x_11168 = v_3570 | ~v_136;
assign x_11169 = v_3570 | ~v_135;
assign x_11170 = v_3570 | ~v_134;
assign x_11171 = v_3570 | ~v_18;
assign x_11172 = v_3570 | ~v_16;
assign x_11173 = v_3570 | ~v_15;
assign x_11174 = v_3570 | ~v_13;
assign x_11175 = v_3570 | ~v_9;
assign x_11176 = ~v_3568 | ~v_3563 | ~v_3558 | v_3569;
assign x_11177 = v_3568 | ~v_1662;
assign x_11178 = v_3568 | ~v_1663;
assign x_11179 = v_3568 | ~v_1664;
assign x_11180 = v_3568 | ~v_1665;
assign x_11181 = v_3568 | ~v_1626;
assign x_11182 = v_3568 | ~v_3490;
assign x_11183 = v_3568 | ~v_1746;
assign x_11184 = v_3568 | ~v_3491;
assign x_11185 = v_3568 | ~v_1747;
assign x_11186 = v_3568 | ~v_1629;
assign x_11187 = v_3568 | ~v_3492;
assign x_11188 = v_3568 | ~v_1748;
assign x_11189 = v_3568 | ~v_3493;
assign x_11190 = v_3568 | ~v_1749;
assign x_11191 = v_3568 | ~v_3516;
assign x_11192 = v_3568 | ~v_3517;
assign x_11193 = v_3568 | ~v_3518;
assign x_11194 = v_3568 | ~v_3519;
assign x_11195 = v_3568 | ~v_3496;
assign x_11196 = v_3568 | ~v_3564;
assign x_11197 = v_3568 | ~v_3565;
assign x_11198 = v_3568 | ~v_3499;
assign x_11199 = v_3568 | ~v_3566;
assign x_11200 = v_3568 | ~v_3567;
assign x_11201 = v_3568 | ~v_1193;
assign x_11202 = v_3568 | ~v_1241;
assign x_11203 = v_3568 | ~v_1194;
assign x_11204 = v_3568 | ~v_1242;
assign x_11205 = v_3568 | ~v_1023;
assign x_11206 = v_3568 | ~v_1024;
assign x_11207 = v_3568 | ~v_1243;
assign x_11208 = v_3568 | ~v_1244;
assign x_11209 = v_3568 | ~v_184;
assign x_11210 = v_3568 | ~v_171;
assign x_11211 = v_3568 | ~v_170;
assign x_11212 = v_3568 | ~v_169;
assign x_11213 = v_3568 | ~v_148;
assign x_11214 = v_3568 | ~v_147;
assign x_11215 = v_3568 | ~v_103;
assign x_11216 = v_3568 | ~v_102;
assign x_11217 = v_3568 | ~v_101;
assign x_11218 = v_3568 | ~v_100;
assign x_11219 = v_3568 | ~v_99;
assign x_11220 = v_3568 | ~v_97;
assign x_11221 = ~v_19 | ~v_131 | v_3567;
assign x_11222 = ~v_19 | ~v_126 | v_3566;
assign x_11223 = v_19 | ~v_116 | v_3565;
assign x_11224 = v_19 | ~v_111 | v_3564;
assign x_11225 = v_3563 | ~v_1653;
assign x_11226 = v_3563 | ~v_1654;
assign x_11227 = v_3563 | ~v_1655;
assign x_11228 = v_3563 | ~v_1656;
assign x_11229 = v_3563 | ~v_1601;
assign x_11230 = v_3563 | ~v_3475;
assign x_11231 = v_3563 | ~v_1737;
assign x_11232 = v_3563 | ~v_3476;
assign x_11233 = v_3563 | ~v_1738;
assign x_11234 = v_3563 | ~v_1604;
assign x_11235 = v_3563 | ~v_3477;
assign x_11236 = v_3563 | ~v_1739;
assign x_11237 = v_3563 | ~v_3478;
assign x_11238 = v_3563 | ~v_1740;
assign x_11239 = v_3563 | ~v_3511;
assign x_11240 = v_3563 | ~v_3512;
assign x_11241 = v_3563 | ~v_3513;
assign x_11242 = v_3563 | ~v_3514;
assign x_11243 = v_3563 | ~v_3481;
assign x_11244 = v_3563 | ~v_3559;
assign x_11245 = v_3563 | ~v_3560;
assign x_11246 = v_3563 | ~v_3484;
assign x_11247 = v_3563 | ~v_1178;
assign x_11248 = v_3563 | ~v_1236;
assign x_11249 = v_3563 | ~v_1179;
assign x_11250 = v_3563 | ~v_1237;
assign x_11251 = v_3563 | ~v_1008;
assign x_11252 = v_3563 | ~v_1009;
assign x_11253 = v_3563 | ~v_3561;
assign x_11254 = v_3563 | ~v_3562;
assign x_11255 = v_3563 | ~v_1238;
assign x_11256 = v_3563 | ~v_1239;
assign x_11257 = v_3563 | ~v_183;
assign x_11258 = v_3563 | ~v_167;
assign x_11259 = v_3563 | ~v_166;
assign x_11260 = v_3563 | ~v_165;
assign x_11261 = v_3563 | ~v_143;
assign x_11262 = v_3563 | ~v_142;
assign x_11263 = v_3563 | ~v_61;
assign x_11264 = v_3563 | ~v_60;
assign x_11265 = v_3563 | ~v_59;
assign x_11266 = v_3563 | ~v_58;
assign x_11267 = v_3563 | ~v_57;
assign x_11268 = v_3563 | ~v_55;
assign x_11269 = ~v_19 | ~v_84 | v_3562;
assign x_11270 = ~v_19 | ~v_89 | v_3561;
assign x_11271 = v_19 | ~v_74 | v_3560;
assign x_11272 = v_19 | ~v_69 | v_3559;
assign x_11273 = v_3558 | ~v_1644;
assign x_11274 = v_3558 | ~v_1645;
assign x_11275 = v_3558 | ~v_1646;
assign x_11276 = v_3558 | ~v_1647;
assign x_11277 = v_3558 | ~v_1576;
assign x_11278 = v_3558 | ~v_3460;
assign x_11279 = v_3558 | ~v_1728;
assign x_11280 = v_3558 | ~v_3461;
assign x_11281 = v_3558 | ~v_1729;
assign x_11282 = v_3558 | ~v_1579;
assign x_11283 = v_3558 | ~v_3462;
assign x_11284 = v_3558 | ~v_1730;
assign x_11285 = v_3558 | ~v_3463;
assign x_11286 = v_3558 | ~v_1731;
assign x_11287 = v_3558 | ~v_3506;
assign x_11288 = v_3558 | ~v_3507;
assign x_11289 = v_3558 | ~v_3508;
assign x_11290 = v_3558 | ~v_3509;
assign x_11291 = v_3558 | ~v_3466;
assign x_11292 = v_3558 | ~v_3554;
assign x_11293 = v_3558 | ~v_3555;
assign x_11294 = v_3558 | ~v_3469;
assign x_11295 = v_3558 | ~v_3556;
assign x_11296 = v_3558 | ~v_3557;
assign x_11297 = v_3558 | ~v_1163;
assign x_11298 = v_3558 | ~v_1231;
assign x_11299 = v_3558 | ~v_1164;
assign x_11300 = v_3558 | ~v_1232;
assign x_11301 = v_3558 | ~v_1233;
assign x_11302 = v_3558 | ~v_1234;
assign x_11303 = v_3558 | ~v_182;
assign x_11304 = v_3558 | ~v_163;
assign x_11305 = v_3558 | ~v_162;
assign x_11306 = v_3558 | ~v_161;
assign x_11307 = v_3558 | ~v_135;
assign x_11308 = v_3558 | ~v_134;
assign x_11309 = v_3558 | ~v_993;
assign x_11310 = v_3558 | ~v_994;
assign x_11311 = v_3558 | ~v_18;
assign x_11312 = v_3558 | ~v_17;
assign x_11313 = v_3558 | ~v_16;
assign x_11314 = v_3558 | ~v_15;
assign x_11315 = v_3558 | ~v_14;
assign x_11316 = v_3558 | ~v_12;
assign x_11317 = ~v_19 | ~v_47 | v_3557;
assign x_11318 = ~v_19 | ~v_42 | v_3556;
assign x_11319 = ~v_32 | v_19 | v_3555;
assign x_11320 = ~v_27 | v_19 | v_3554;
assign x_11321 = ~v_3552 | ~v_3547 | ~v_3542 | v_3553;
assign x_11322 = v_3552 | ~v_1662;
assign x_11323 = v_3552 | ~v_1663;
assign x_11324 = v_3552 | ~v_1664;
assign x_11325 = v_3552 | ~v_1665;
assign x_11326 = v_3552 | ~v_1718;
assign x_11327 = v_3552 | ~v_1719;
assign x_11328 = v_3552 | ~v_1720;
assign x_11329 = v_3552 | ~v_1721;
assign x_11330 = v_3552 | ~v_1626;
assign x_11331 = v_3552 | ~v_3490;
assign x_11332 = v_3552 | ~v_3491;
assign x_11333 = v_3552 | ~v_1629;
assign x_11334 = v_3552 | ~v_3492;
assign x_11335 = v_3552 | ~v_3493;
assign x_11336 = v_3552 | ~v_3516;
assign x_11337 = v_3552 | ~v_3517;
assign x_11338 = v_3552 | ~v_3518;
assign x_11339 = v_3552 | ~v_3519;
assign x_11340 = v_3552 | ~v_3548;
assign x_11341 = v_3552 | ~v_3549;
assign x_11342 = v_3552 | ~v_3550;
assign x_11343 = v_3552 | ~v_3551;
assign x_11344 = v_3552 | ~v_3496;
assign x_11345 = v_3552 | ~v_3499;
assign x_11346 = v_3552 | ~v_1191;
assign x_11347 = v_3552 | ~v_1192;
assign x_11348 = v_3552 | ~v_1193;
assign x_11349 = v_3552 | ~v_1194;
assign x_11350 = v_3552 | ~v_837;
assign x_11351 = v_3552 | ~v_838;
assign x_11352 = v_3552 | ~v_1195;
assign x_11353 = v_3552 | ~v_1196;
assign x_11354 = v_3552 | ~v_184;
assign x_11355 = v_3552 | ~v_171;
assign x_11356 = v_3552 | ~v_170;
assign x_11357 = v_3552 | ~v_169;
assign x_11358 = v_3552 | ~v_160;
assign x_11359 = v_3552 | ~v_151;
assign x_11360 = v_3552 | ~v_150;
assign x_11361 = v_3552 | ~v_149;
assign x_11362 = v_3552 | ~v_147;
assign x_11363 = v_3552 | ~v_103;
assign x_11364 = v_3552 | ~v_100;
assign x_11365 = v_3552 | ~v_96;
assign x_11366 = ~v_131 | ~v_157 | v_3551;
assign x_11367 = ~v_126 | ~v_156 | v_3550;
assign x_11368 = ~v_116 | v_157 | v_3549;
assign x_11369 = ~v_111 | v_156 | v_3548;
assign x_11370 = v_3547 | ~v_1653;
assign x_11371 = v_3547 | ~v_1654;
assign x_11372 = v_3547 | ~v_1655;
assign x_11373 = v_3547 | ~v_1656;
assign x_11374 = v_3547 | ~v_1709;
assign x_11375 = v_3547 | ~v_1710;
assign x_11376 = v_3547 | ~v_1711;
assign x_11377 = v_3547 | ~v_1712;
assign x_11378 = v_3547 | ~v_1601;
assign x_11379 = v_3547 | ~v_3475;
assign x_11380 = v_3547 | ~v_3476;
assign x_11381 = v_3547 | ~v_1604;
assign x_11382 = v_3547 | ~v_3477;
assign x_11383 = v_3547 | ~v_3478;
assign x_11384 = v_3547 | ~v_3511;
assign x_11385 = v_3547 | ~v_3512;
assign x_11386 = v_3547 | ~v_3513;
assign x_11387 = v_3547 | ~v_3514;
assign x_11388 = v_3547 | ~v_3543;
assign x_11389 = v_3547 | ~v_3544;
assign x_11390 = v_3547 | ~v_3545;
assign x_11391 = v_3547 | ~v_3546;
assign x_11392 = v_3547 | ~v_3481;
assign x_11393 = v_3547 | ~v_3484;
assign x_11394 = v_3547 | ~v_1176;
assign x_11395 = v_3547 | ~v_1177;
assign x_11396 = v_3547 | ~v_1178;
assign x_11397 = v_3547 | ~v_1179;
assign x_11398 = v_3547 | ~v_804;
assign x_11399 = v_3547 | ~v_805;
assign x_11400 = v_3547 | ~v_1180;
assign x_11401 = v_3547 | ~v_1181;
assign x_11402 = v_3547 | ~v_183;
assign x_11403 = v_3547 | ~v_167;
assign x_11404 = v_3547 | ~v_166;
assign x_11405 = v_3547 | ~v_165;
assign x_11406 = v_3547 | ~v_159;
assign x_11407 = v_3547 | ~v_146;
assign x_11408 = v_3547 | ~v_145;
assign x_11409 = v_3547 | ~v_144;
assign x_11410 = v_3547 | ~v_142;
assign x_11411 = v_3547 | ~v_61;
assign x_11412 = v_3547 | ~v_58;
assign x_11413 = v_3547 | ~v_54;
assign x_11414 = ~v_89 | ~v_157 | v_3546;
assign x_11415 = ~v_84 | ~v_156 | v_3545;
assign x_11416 = ~v_74 | v_157 | v_3544;
assign x_11417 = ~v_69 | v_156 | v_3543;
assign x_11418 = v_3542 | ~v_1644;
assign x_11419 = v_3542 | ~v_1645;
assign x_11420 = v_3542 | ~v_1646;
assign x_11421 = v_3542 | ~v_1647;
assign x_11422 = v_3542 | ~v_1700;
assign x_11423 = v_3542 | ~v_1701;
assign x_11424 = v_3542 | ~v_1702;
assign x_11425 = v_3542 | ~v_1703;
assign x_11426 = v_3542 | ~v_1576;
assign x_11427 = v_3542 | ~v_3460;
assign x_11428 = v_3542 | ~v_3461;
assign x_11429 = v_3542 | ~v_1579;
assign x_11430 = v_3542 | ~v_3462;
assign x_11431 = v_3542 | ~v_3463;
assign x_11432 = v_3542 | ~v_3506;
assign x_11433 = v_3542 | ~v_3507;
assign x_11434 = v_3542 | ~v_3508;
assign x_11435 = v_3542 | ~v_3509;
assign x_11436 = v_3542 | ~v_3538;
assign x_11437 = v_3542 | ~v_3539;
assign x_11438 = v_3542 | ~v_3540;
assign x_11439 = v_3542 | ~v_3541;
assign x_11440 = v_3542 | ~v_3466;
assign x_11441 = v_3542 | ~v_3469;
assign x_11442 = v_3542 | ~v_1161;
assign x_11443 = v_3542 | ~v_1162;
assign x_11444 = v_3542 | ~v_1163;
assign x_11445 = v_3542 | ~v_1164;
assign x_11446 = v_3542 | ~v_771;
assign x_11447 = v_3542 | ~v_772;
assign x_11448 = v_3542 | ~v_1165;
assign x_11449 = v_3542 | ~v_1166;
assign x_11450 = v_3542 | ~v_182;
assign x_11451 = v_3542 | ~v_163;
assign x_11452 = v_3542 | ~v_162;
assign x_11453 = v_3542 | ~v_161;
assign x_11454 = v_3542 | ~v_155;
assign x_11455 = v_3542 | ~v_138;
assign x_11456 = v_3542 | ~v_137;
assign x_11457 = v_3542 | ~v_136;
assign x_11458 = v_3542 | ~v_134;
assign x_11459 = v_3542 | ~v_18;
assign x_11460 = v_3542 | ~v_15;
assign x_11461 = v_3542 | ~v_11;
assign x_11462 = ~v_47 | ~v_157 | v_3541;
assign x_11463 = ~v_42 | ~v_156 | v_3540;
assign x_11464 = ~v_32 | v_157 | v_3539;
assign x_11465 = ~v_27 | v_156 | v_3538;
assign x_11466 = ~v_3536 | ~v_3531 | ~v_3526 | v_3537;
assign x_11467 = v_3536 | ~v_1662;
assign x_11468 = v_3536 | ~v_1663;
assign x_11469 = v_3536 | ~v_1664;
assign x_11470 = v_3536 | ~v_1665;
assign x_11471 = v_3536 | ~v_1690;
assign x_11472 = v_3536 | ~v_1691;
assign x_11473 = v_3536 | ~v_1692;
assign x_11474 = v_3536 | ~v_1693;
assign x_11475 = v_3536 | ~v_1626;
assign x_11476 = v_3536 | ~v_3490;
assign x_11477 = v_3536 | ~v_3491;
assign x_11478 = v_3536 | ~v_1629;
assign x_11479 = v_3536 | ~v_3492;
assign x_11480 = v_3536 | ~v_3493;
assign x_11481 = v_3536 | ~v_3516;
assign x_11482 = v_3536 | ~v_3517;
assign x_11483 = v_3536 | ~v_3518;
assign x_11484 = v_3536 | ~v_3519;
assign x_11485 = v_3536 | ~v_3532;
assign x_11486 = v_3536 | ~v_3533;
assign x_11487 = v_3536 | ~v_3534;
assign x_11488 = v_3536 | ~v_3535;
assign x_11489 = v_3536 | ~v_3496;
assign x_11490 = v_3536 | ~v_3499;
assign x_11491 = v_3536 | ~v_1209;
assign x_11492 = v_3536 | ~v_1210;
assign x_11493 = v_3536 | ~v_1193;
assign x_11494 = v_3536 | ~v_1194;
assign x_11495 = v_3536 | ~v_927;
assign x_11496 = v_3536 | ~v_928;
assign x_11497 = v_3536 | ~v_1211;
assign x_11498 = v_3536 | ~v_1212;
assign x_11499 = v_3536 | ~v_184;
assign x_11500 = v_3536 | ~v_172;
assign x_11501 = v_3536 | ~v_171;
assign x_11502 = v_3536 | ~v_170;
assign x_11503 = v_3536 | ~v_169;
assign x_11504 = v_3536 | ~v_150;
assign x_11505 = v_3536 | ~v_149;
assign x_11506 = v_3536 | ~v_148;
assign x_11507 = v_3536 | ~v_147;
assign x_11508 = v_3536 | ~v_102;
assign x_11509 = v_3536 | ~v_101;
assign x_11510 = v_3536 | ~v_100;
assign x_11511 = ~v_131 | ~v_140 | v_3535;
assign x_11512 = ~v_126 | ~v_139 | v_3534;
assign x_11513 = ~v_116 | v_140 | v_3533;
assign x_11514 = ~v_111 | v_139 | v_3532;
assign x_11515 = v_3531 | ~v_1653;
assign x_11516 = v_3531 | ~v_1654;
assign x_11517 = v_3531 | ~v_1655;
assign x_11518 = v_3531 | ~v_1656;
assign x_11519 = v_3531 | ~v_1681;
assign x_11520 = v_3531 | ~v_1682;
assign x_11521 = v_3531 | ~v_1683;
assign x_11522 = v_3531 | ~v_1684;
assign x_11523 = v_3531 | ~v_1601;
assign x_11524 = v_3531 | ~v_3475;
assign x_11525 = v_3531 | ~v_3476;
assign x_11526 = v_3531 | ~v_1604;
assign x_11527 = v_3531 | ~v_3477;
assign x_11528 = v_3531 | ~v_3478;
assign x_11529 = v_3531 | ~v_3511;
assign x_11530 = v_3531 | ~v_3512;
assign x_11531 = v_3531 | ~v_3513;
assign x_11532 = v_3531 | ~v_3514;
assign x_11533 = v_3531 | ~v_3527;
assign x_11534 = v_3531 | ~v_3528;
assign x_11535 = v_3531 | ~v_3529;
assign x_11536 = v_3531 | ~v_3530;
assign x_11537 = v_3531 | ~v_3481;
assign x_11538 = v_3531 | ~v_3484;
assign x_11539 = v_3531 | ~v_1204;
assign x_11540 = v_3531 | ~v_1205;
assign x_11541 = v_3531 | ~v_1178;
assign x_11542 = v_3531 | ~v_1179;
assign x_11543 = v_3531 | ~v_912;
assign x_11544 = v_3531 | ~v_913;
assign x_11545 = v_3531 | ~v_1206;
assign x_11546 = v_3531 | ~v_1207;
assign x_11547 = v_3531 | ~v_183;
assign x_11548 = v_3531 | ~v_168;
assign x_11549 = v_3531 | ~v_167;
assign x_11550 = v_3531 | ~v_166;
assign x_11551 = v_3531 | ~v_165;
assign x_11552 = v_3531 | ~v_145;
assign x_11553 = v_3531 | ~v_144;
assign x_11554 = v_3531 | ~v_143;
assign x_11555 = v_3531 | ~v_142;
assign x_11556 = v_3531 | ~v_60;
assign x_11557 = v_3531 | ~v_59;
assign x_11558 = v_3531 | ~v_58;
assign x_11559 = ~v_89 | ~v_140 | v_3530;
assign x_11560 = ~v_84 | ~v_139 | v_3529;
assign x_11561 = ~v_74 | v_140 | v_3528;
assign x_11562 = ~v_69 | v_139 | v_3527;
assign x_11563 = v_3526 | ~v_1644;
assign x_11564 = v_3526 | ~v_1645;
assign x_11565 = v_3526 | ~v_1646;
assign x_11566 = v_3526 | ~v_1647;
assign x_11567 = v_3526 | ~v_1672;
assign x_11568 = v_3526 | ~v_1673;
assign x_11569 = v_3526 | ~v_1674;
assign x_11570 = v_3526 | ~v_1675;
assign x_11571 = v_3526 | ~v_1576;
assign x_11572 = v_3526 | ~v_3460;
assign x_11573 = v_3526 | ~v_3461;
assign x_11574 = v_3526 | ~v_1579;
assign x_11575 = v_3526 | ~v_3462;
assign x_11576 = v_3526 | ~v_3463;
assign x_11577 = v_3526 | ~v_3506;
assign x_11578 = v_3526 | ~v_3507;
assign x_11579 = v_3526 | ~v_3508;
assign x_11580 = v_3526 | ~v_3509;
assign x_11581 = v_3526 | ~v_3522;
assign x_11582 = v_3526 | ~v_3523;
assign x_11583 = v_3526 | ~v_3524;
assign x_11584 = v_3526 | ~v_3525;
assign x_11585 = v_3526 | ~v_3466;
assign x_11586 = v_3526 | ~v_3469;
assign x_11587 = v_3526 | ~v_1199;
assign x_11588 = v_3526 | ~v_1200;
assign x_11589 = v_3526 | ~v_1163;
assign x_11590 = v_3526 | ~v_1164;
assign x_11591 = v_3526 | ~v_897;
assign x_11592 = v_3526 | ~v_898;
assign x_11593 = v_3526 | ~v_1201;
assign x_11594 = v_3526 | ~v_1202;
assign x_11595 = v_3526 | ~v_182;
assign x_11596 = v_3526 | ~v_164;
assign x_11597 = v_3526 | ~v_163;
assign x_11598 = v_3526 | ~v_162;
assign x_11599 = v_3526 | ~v_161;
assign x_11600 = v_3526 | ~v_137;
assign x_11601 = v_3526 | ~v_136;
assign x_11602 = v_3526 | ~v_135;
assign x_11603 = v_3526 | ~v_134;
assign x_11604 = v_3526 | ~v_17;
assign x_11605 = v_3526 | ~v_16;
assign x_11606 = v_3526 | ~v_15;
assign x_11607 = ~v_47 | ~v_140 | v_3525;
assign x_11608 = ~v_42 | ~v_139 | v_3524;
assign x_11609 = ~v_32 | v_140 | v_3523;
assign x_11610 = ~v_27 | v_139 | v_3522;
assign x_11611 = ~v_3520 | ~v_3515 | ~v_3510 | v_3521;
assign x_11612 = v_3520 | ~v_1662;
assign x_11613 = v_3520 | ~v_1663;
assign x_11614 = v_3520 | ~v_1664;
assign x_11615 = v_3520 | ~v_1665;
assign x_11616 = v_3520 | ~v_1622;
assign x_11617 = v_3520 | ~v_1623;
assign x_11618 = v_3520 | ~v_1624;
assign x_11619 = v_3520 | ~v_1625;
assign x_11620 = v_3520 | ~v_1626;
assign x_11621 = v_3520 | ~v_3490;
assign x_11622 = v_3520 | ~v_3491;
assign x_11623 = v_3520 | ~v_1629;
assign x_11624 = v_3520 | ~v_3492;
assign x_11625 = v_3520 | ~v_3493;
assign x_11626 = v_3520 | ~v_3516;
assign x_11627 = v_3520 | ~v_3517;
assign x_11628 = v_3520 | ~v_3518;
assign x_11629 = v_3520 | ~v_3519;
assign x_11630 = v_3520 | ~v_3494;
assign x_11631 = v_3520 | ~v_3495;
assign x_11632 = v_3520 | ~v_3496;
assign x_11633 = v_3520 | ~v_3499;
assign x_11634 = v_3520 | ~v_1225;
assign x_11635 = v_3520 | ~v_1226;
assign x_11636 = v_3520 | ~v_1227;
assign x_11637 = v_3520 | ~v_1228;
assign x_11638 = v_3520 | ~v_1193;
assign x_11639 = v_3520 | ~v_1194;
assign x_11640 = v_3520 | ~v_975;
assign x_11641 = v_3520 | ~v_976;
assign x_11642 = v_3520 | ~v_3502;
assign x_11643 = v_3520 | ~v_3503;
assign x_11644 = v_3520 | ~v_184;
assign x_11645 = v_3520 | ~v_171;
assign x_11646 = v_3520 | ~v_170;
assign x_11647 = v_3520 | ~v_169;
assign x_11648 = v_3520 | ~v_150;
assign x_11649 = v_3520 | ~v_149;
assign x_11650 = v_3520 | ~v_148;
assign x_11651 = v_3520 | ~v_103;
assign x_11652 = v_3520 | ~v_102;
assign x_11653 = v_3520 | ~v_101;
assign x_11654 = v_3520 | ~v_100;
assign x_11655 = v_3520 | ~v_95;
assign x_11656 = ~v_128 | ~v_153 | v_3519;
assign x_11657 = ~v_125 | ~v_152 | v_3518;
assign x_11658 = ~v_113 | v_153 | v_3517;
assign x_11659 = ~v_110 | v_152 | v_3516;
assign x_11660 = v_3515 | ~v_1653;
assign x_11661 = v_3515 | ~v_1654;
assign x_11662 = v_3515 | ~v_1655;
assign x_11663 = v_3515 | ~v_1656;
assign x_11664 = v_3515 | ~v_1597;
assign x_11665 = v_3515 | ~v_1598;
assign x_11666 = v_3515 | ~v_1599;
assign x_11667 = v_3515 | ~v_1600;
assign x_11668 = v_3515 | ~v_1601;
assign x_11669 = v_3515 | ~v_3475;
assign x_11670 = v_3515 | ~v_3476;
assign x_11671 = v_3515 | ~v_1604;
assign x_11672 = v_3515 | ~v_3477;
assign x_11673 = v_3515 | ~v_3478;
assign x_11674 = v_3515 | ~v_3511;
assign x_11675 = v_3515 | ~v_3512;
assign x_11676 = v_3515 | ~v_3513;
assign x_11677 = v_3515 | ~v_3514;
assign x_11678 = v_3515 | ~v_3479;
assign x_11679 = v_3515 | ~v_3480;
assign x_11680 = v_3515 | ~v_3481;
assign x_11681 = v_3515 | ~v_3484;
assign x_11682 = v_3515 | ~v_1220;
assign x_11683 = v_3515 | ~v_1221;
assign x_11684 = v_3515 | ~v_1222;
assign x_11685 = v_3515 | ~v_1223;
assign x_11686 = v_3515 | ~v_1178;
assign x_11687 = v_3515 | ~v_1179;
assign x_11688 = v_3515 | ~v_960;
assign x_11689 = v_3515 | ~v_961;
assign x_11690 = v_3515 | ~v_3487;
assign x_11691 = v_3515 | ~v_3488;
assign x_11692 = v_3515 | ~v_183;
assign x_11693 = v_3515 | ~v_167;
assign x_11694 = v_3515 | ~v_166;
assign x_11695 = v_3515 | ~v_165;
assign x_11696 = v_3515 | ~v_145;
assign x_11697 = v_3515 | ~v_144;
assign x_11698 = v_3515 | ~v_143;
assign x_11699 = v_3515 | ~v_61;
assign x_11700 = v_3515 | ~v_60;
assign x_11701 = v_3515 | ~v_59;
assign x_11702 = v_3515 | ~v_58;
assign x_11703 = v_3515 | ~v_53;
assign x_11704 = ~v_86 | ~v_153 | v_3514;
assign x_11705 = ~v_83 | ~v_152 | v_3513;
assign x_11706 = ~v_71 | v_153 | v_3512;
assign x_11707 = ~v_68 | v_152 | v_3511;
assign x_11708 = v_3510 | ~v_1644;
assign x_11709 = v_3510 | ~v_1645;
assign x_11710 = v_3510 | ~v_1646;
assign x_11711 = v_3510 | ~v_1647;
assign x_11712 = v_3510 | ~v_1572;
assign x_11713 = v_3510 | ~v_1573;
assign x_11714 = v_3510 | ~v_1574;
assign x_11715 = v_3510 | ~v_1575;
assign x_11716 = v_3510 | ~v_1576;
assign x_11717 = v_3510 | ~v_3460;
assign x_11718 = v_3510 | ~v_3461;
assign x_11719 = v_3510 | ~v_1579;
assign x_11720 = v_3510 | ~v_3462;
assign x_11721 = v_3510 | ~v_3463;
assign x_11722 = v_3510 | ~v_3506;
assign x_11723 = v_3510 | ~v_3507;
assign x_11724 = v_3510 | ~v_3508;
assign x_11725 = v_3510 | ~v_3509;
assign x_11726 = v_3510 | ~v_3464;
assign x_11727 = v_3510 | ~v_3465;
assign x_11728 = v_3510 | ~v_3466;
assign x_11729 = v_3510 | ~v_3469;
assign x_11730 = v_3510 | ~v_1215;
assign x_11731 = v_3510 | ~v_1216;
assign x_11732 = v_3510 | ~v_1217;
assign x_11733 = v_3510 | ~v_1218;
assign x_11734 = v_3510 | ~v_1163;
assign x_11735 = v_3510 | ~v_1164;
assign x_11736 = v_3510 | ~v_945;
assign x_11737 = v_3510 | ~v_946;
assign x_11738 = v_3510 | ~v_3471;
assign x_11739 = v_3510 | ~v_3472;
assign x_11740 = v_3510 | ~v_182;
assign x_11741 = v_3510 | ~v_163;
assign x_11742 = v_3510 | ~v_162;
assign x_11743 = v_3510 | ~v_161;
assign x_11744 = v_3510 | ~v_137;
assign x_11745 = v_3510 | ~v_136;
assign x_11746 = v_3510 | ~v_135;
assign x_11747 = v_3510 | ~v_18;
assign x_11748 = v_3510 | ~v_17;
assign x_11749 = v_3510 | ~v_16;
assign x_11750 = v_3510 | ~v_15;
assign x_11751 = v_3510 | ~v_10;
assign x_11752 = ~v_44 | ~v_153 | v_3509;
assign x_11753 = ~v_41 | ~v_152 | v_3508;
assign x_11754 = ~v_29 | v_153 | v_3507;
assign x_11755 = ~v_26 | v_152 | v_3506;
assign x_11756 = ~v_3504 | ~v_3489 | ~v_3474 | v_3505;
assign x_11757 = v_3504 | ~v_1622;
assign x_11758 = v_3504 | ~v_1623;
assign x_11759 = v_3504 | ~v_1624;
assign x_11760 = v_3504 | ~v_1625;
assign x_11761 = v_3504 | ~v_1626;
assign x_11762 = v_3504 | ~v_3490;
assign x_11763 = v_3504 | ~v_1627;
assign x_11764 = v_3504 | ~v_3491;
assign x_11765 = v_3504 | ~v_1628;
assign x_11766 = v_3504 | ~v_1629;
assign x_11767 = v_3504 | ~v_3492;
assign x_11768 = v_3504 | ~v_1630;
assign x_11769 = v_3504 | ~v_3493;
assign x_11770 = v_3504 | ~v_1631;
assign x_11771 = v_3504 | ~v_3494;
assign x_11772 = v_3504 | ~v_3495;
assign x_11773 = v_3504 | ~v_3496;
assign x_11774 = v_3504 | ~v_3497;
assign x_11775 = v_3504 | ~v_3498;
assign x_11776 = v_3504 | ~v_3499;
assign x_11777 = v_3504 | ~v_3500;
assign x_11778 = v_3504 | ~v_3501;
assign x_11779 = v_3504 | ~v_1147;
assign x_11780 = v_3504 | ~v_1148;
assign x_11781 = v_3504 | ~v_975;
assign x_11782 = v_3504 | ~v_976;
assign x_11783 = v_3504 | ~v_839;
assign x_11784 = v_3504 | ~v_840;
assign x_11785 = v_3504 | ~v_1149;
assign x_11786 = v_3504 | ~v_1150;
assign x_11787 = v_3504 | ~v_3502;
assign x_11788 = v_3504 | ~v_3503;
assign x_11789 = v_3504 | ~v_184;
assign x_11790 = v_3504 | ~v_169;
assign x_11791 = v_3504 | ~v_150;
assign x_11792 = v_3504 | ~v_149;
assign x_11793 = v_3504 | ~v_148;
assign x_11794 = v_3504 | ~v_147;
assign x_11795 = v_3504 | ~v_103;
assign x_11796 = v_3504 | ~v_102;
assign x_11797 = v_3504 | ~v_101;
assign x_11798 = v_3504 | ~v_100;
assign x_11799 = v_3504 | ~v_98;
assign x_11800 = v_3504 | ~v_94;
assign x_11801 = ~v_131 | ~v_153 | v_3503;
assign x_11802 = ~v_116 | v_153 | v_3502;
assign x_11803 = ~v_19 | ~v_128 | v_3501;
assign x_11804 = ~v_19 | ~v_125 | v_3500;
assign x_11805 = ~v_19 | ~v_124 | v_3499;
assign x_11806 = v_19 | ~v_113 | v_3498;
assign x_11807 = v_19 | ~v_110 | v_3497;
assign x_11808 = v_19 | ~v_109 | v_3496;
assign x_11809 = ~v_126 | ~v_152 | v_3495;
assign x_11810 = ~v_111 | v_152 | v_3494;
assign x_11811 = ~v_123 | ~v_156 | v_3493;
assign x_11812 = ~v_120 | ~v_157 | v_3492;
assign x_11813 = ~v_108 | v_156 | v_3491;
assign x_11814 = ~v_105 | v_157 | v_3490;
assign x_11815 = v_3489 | ~v_1597;
assign x_11816 = v_3489 | ~v_1598;
assign x_11817 = v_3489 | ~v_1599;
assign x_11818 = v_3489 | ~v_1600;
assign x_11819 = v_3489 | ~v_1601;
assign x_11820 = v_3489 | ~v_3475;
assign x_11821 = v_3489 | ~v_1602;
assign x_11822 = v_3489 | ~v_3476;
assign x_11823 = v_3489 | ~v_1603;
assign x_11824 = v_3489 | ~v_1604;
assign x_11825 = v_3489 | ~v_3477;
assign x_11826 = v_3489 | ~v_1605;
assign x_11827 = v_3489 | ~v_3478;
assign x_11828 = v_3489 | ~v_1606;
assign x_11829 = v_3489 | ~v_3479;
assign x_11830 = v_3489 | ~v_3480;
assign x_11831 = v_3489 | ~v_3481;
assign x_11832 = v_3489 | ~v_3482;
assign x_11833 = v_3489 | ~v_3483;
assign x_11834 = v_3489 | ~v_3484;
assign x_11835 = v_3489 | ~v_3485;
assign x_11836 = v_3489 | ~v_1142;
assign x_11837 = v_3489 | ~v_1143;
assign x_11838 = v_3489 | ~v_960;
assign x_11839 = v_3489 | ~v_961;
assign x_11840 = v_3489 | ~v_806;
assign x_11841 = v_3489 | ~v_807;
assign x_11842 = v_3489 | ~v_3486;
assign x_11843 = v_3489 | ~v_1144;
assign x_11844 = v_3489 | ~v_1145;
assign x_11845 = v_3489 | ~v_3487;
assign x_11846 = v_3489 | ~v_3488;
assign x_11847 = v_3489 | ~v_183;
assign x_11848 = v_3489 | ~v_165;
assign x_11849 = v_3489 | ~v_145;
assign x_11850 = v_3489 | ~v_144;
assign x_11851 = v_3489 | ~v_143;
assign x_11852 = v_3489 | ~v_142;
assign x_11853 = v_3489 | ~v_61;
assign x_11854 = v_3489 | ~v_60;
assign x_11855 = v_3489 | ~v_59;
assign x_11856 = v_3489 | ~v_58;
assign x_11857 = v_3489 | ~v_56;
assign x_11858 = v_3489 | ~v_52;
assign x_11859 = ~v_89 | ~v_153 | v_3488;
assign x_11860 = ~v_74 | v_153 | v_3487;
assign x_11861 = ~v_19 | ~v_83 | v_3486;
assign x_11862 = ~v_19 | ~v_86 | v_3485;
assign x_11863 = ~v_19 | ~v_82 | v_3484;
assign x_11864 = v_19 | ~v_71 | v_3483;
assign x_11865 = v_19 | ~v_68 | v_3482;
assign x_11866 = v_19 | ~v_67 | v_3481;
assign x_11867 = ~v_84 | ~v_152 | v_3480;
assign x_11868 = ~v_69 | v_152 | v_3479;
assign x_11869 = ~v_81 | ~v_156 | v_3478;
assign x_11870 = ~v_78 | ~v_157 | v_3477;
assign x_11871 = ~v_66 | v_156 | v_3476;
assign x_11872 = ~v_63 | v_157 | v_3475;
assign x_11873 = v_3474 | ~v_1572;
assign x_11874 = v_3474 | ~v_1573;
assign x_11875 = v_3474 | ~v_1574;
assign x_11876 = v_3474 | ~v_1575;
assign x_11877 = v_3474 | ~v_1576;
assign x_11878 = v_3474 | ~v_3460;
assign x_11879 = v_3474 | ~v_1577;
assign x_11880 = v_3474 | ~v_3461;
assign x_11881 = v_3474 | ~v_1578;
assign x_11882 = v_3474 | ~v_1579;
assign x_11883 = v_3474 | ~v_3462;
assign x_11884 = v_3474 | ~v_1580;
assign x_11885 = v_3474 | ~v_3463;
assign x_11886 = v_3474 | ~v_1581;
assign x_11887 = v_3474 | ~v_3464;
assign x_11888 = v_3474 | ~v_3465;
assign x_11889 = v_3474 | ~v_3466;
assign x_11890 = v_3474 | ~v_3467;
assign x_11891 = v_3474 | ~v_3468;
assign x_11892 = v_3474 | ~v_3469;
assign x_11893 = v_3474 | ~v_3470;
assign x_11894 = v_3474 | ~v_1137;
assign x_11895 = v_3474 | ~v_1138;
assign x_11896 = v_3474 | ~v_945;
assign x_11897 = v_3474 | ~v_946;
assign x_11898 = v_3474 | ~v_773;
assign x_11899 = v_3474 | ~v_774;
assign x_11900 = v_3474 | ~v_1139;
assign x_11901 = v_3474 | ~v_1140;
assign x_11902 = v_3474 | ~v_3471;
assign x_11903 = v_3474 | ~v_3472;
assign x_11904 = v_3474 | ~v_182;
assign x_11905 = v_3474 | ~v_161;
assign x_11906 = v_3474 | ~v_137;
assign x_11907 = v_3474 | ~v_3473;
assign x_11908 = v_3474 | ~v_136;
assign x_11909 = v_3474 | ~v_135;
assign x_11910 = v_3474 | ~v_134;
assign x_11911 = v_3474 | ~v_18;
assign x_11912 = v_3474 | ~v_17;
assign x_11913 = v_3474 | ~v_16;
assign x_11914 = v_3474 | ~v_15;
assign x_11915 = v_3474 | ~v_13;
assign x_11916 = v_3474 | ~v_9;
assign x_11917 = ~v_19 | ~v_41 | v_3473;
assign x_11918 = ~v_47 | ~v_153 | v_3472;
assign x_11919 = ~v_32 | v_153 | v_3471;
assign x_11920 = ~v_19 | ~v_44 | v_3470;
assign x_11921 = ~v_19 | ~v_40 | v_3469;
assign x_11922 = ~v_29 | v_19 | v_3468;
assign x_11923 = ~v_26 | v_19 | v_3467;
assign x_11924 = ~v_25 | v_19 | v_3466;
assign x_11925 = ~v_42 | ~v_152 | v_3465;
assign x_11926 = ~v_27 | v_152 | v_3464;
assign x_11927 = ~v_39 | ~v_156 | v_3463;
assign x_11928 = ~v_36 | ~v_157 | v_3462;
assign x_11929 = ~v_24 | v_156 | v_3461;
assign x_11930 = ~v_21 | v_157 | v_3460;
assign x_11931 = v_3459 | ~v_2406;
assign x_11932 = v_3459 | ~v_735;
assign x_11933 = v_3458 | ~v_1566;
assign x_11934 = v_3458 | ~v_730;
assign x_11935 = ~v_725 | ~v_724 | ~v_723 | ~v_722 | ~v_3456 | ~v_3452 | ~v_3448 | ~v_3444 | ~v_3440 | ~v_3424 | ~v_3420 | ~v_3416 | ~v_3412 | ~v_3408 | ~v_3392 | ~v_3388 | ~v_3372 | ~v_3356 | ~v_3340 | ~v_3324 | ~v_3278 | v_3457;
assign x_11936 = v_3456 | ~v_3453;
assign x_11937 = v_3456 | ~v_3454;
assign x_11938 = v_3456 | ~v_3455;
assign x_11939 = v_98 | v_103 | v_101 | v_97 | v_100 | v_95 | v_94 | v_99 | v_102 | ~v_719 | ~v_718 | v_169 | v_148 | v_184 | ~v_483 | ~v_717 | ~v_299 | ~v_482 | ~v_716 | ~v_298 | ~v_3386 | ~v_3320 | ~v_3385 | ~v_3319 | ~v_3318 | ~v_3384 | ~v_3317 | ~v_3383 | ~v_3316 | ~v_3315 | ~v_1460 | ~v_1342 | ~v_3312 | ~v_1459 | ~v_1341 | ~v_3311 | ~v_1340 | ~v_1458 | ~v_1339 | ~v_3310 | ~v_1457 | ~v_1338 | ~v_3309 | ~v_1337 | v_3455;
assign x_11940 = v_53 | v_56 | v_55 | v_61 | v_52 | v_60 | v_59 | v_58 | v_57 | ~v_714 | ~v_713 | v_143 | v_165 | v_183 | ~v_3381 | ~v_3305 | ~v_266 | ~v_3380 | ~v_468 | ~v_712 | ~v_467 | ~v_711 | ~v_265 | ~v_3304 | ~v_3303 | ~v_3379 | ~v_3302 | ~v_3378 | ~v_3301 | ~v_3300 | ~v_1451 | ~v_1317 | ~v_3297 | ~v_1450 | ~v_1316 | ~v_3296 | ~v_1315 | ~v_1449 | ~v_1314 | ~v_3295 | ~v_1448 | ~v_1313 | ~v_3294 | ~v_1312 | v_3454;
assign x_11941 = v_13 | v_9 | v_18 | v_17 | v_16 | v_15 | v_14 | v_12 | v_10 | ~v_453 | ~v_709 | ~v_452 | ~v_708 | v_135 | ~v_707 | ~v_706 | ~v_3292 | v_161 | v_182 | ~v_233 | ~v_232 | ~v_3376 | ~v_3289 | ~v_3375 | ~v_3288 | ~v_3374 | ~v_3287 | ~v_3373 | ~v_3286 | ~v_3285 | ~v_1442 | ~v_1292 | ~v_3282 | ~v_1441 | ~v_1291 | ~v_3281 | ~v_1290 | ~v_1440 | ~v_1289 | ~v_3280 | ~v_1439 | ~v_1288 | ~v_3279 | ~v_1287 | v_3453;
assign x_11942 = v_3452 | ~v_3449;
assign x_11943 = v_3452 | ~v_3450;
assign x_11944 = v_3452 | ~v_3451;
assign x_11945 = v_103 | v_101 | v_97 | v_99 | v_93 | v_102 | v_171 | v_170 | v_148 | v_147 | v_184 | v_181 | ~v_483 | ~v_482 | ~v_481 | ~v_480 | ~v_345 | ~v_479 | ~v_478 | ~v_344 | ~v_3386 | ~v_3385 | ~v_3318 | ~v_3384 | ~v_3383 | ~v_3315 | ~v_3438 | ~v_3437 | ~v_3436 | ~v_3435 | ~v_1460 | ~v_3312 | ~v_1459 | ~v_3311 | ~v_1340 | ~v_1458 | ~v_3310 | ~v_1457 | ~v_3309 | ~v_1337 | ~v_1536 | ~v_1535 | ~v_1534 | ~v_1533 | v_3451;
assign x_11946 = v_55 | v_61 | v_51 | v_60 | v_59 | v_57 | v_180 | v_143 | v_142 | v_167 | v_166 | v_183 | ~v_3381 | ~v_3380 | ~v_468 | ~v_467 | ~v_466 | ~v_465 | ~v_330 | ~v_464 | ~v_463 | ~v_329 | ~v_3303 | ~v_3379 | ~v_3378 | ~v_3300 | ~v_3433 | ~v_3432 | ~v_3431 | ~v_3430 | ~v_1451 | ~v_3297 | ~v_1450 | ~v_3296 | ~v_1315 | ~v_1449 | ~v_3295 | ~v_1448 | ~v_3294 | ~v_1312 | ~v_1527 | ~v_1526 | ~v_1525 | ~v_1524 | v_3450;
assign x_11947 = v_18 | v_17 | v_16 | v_8 | v_14 | v_12 | ~v_453 | ~v_452 | v_135 | v_134 | v_179 | v_163 | v_162 | v_182 | ~v_451 | ~v_450 | ~v_315 | ~v_449 | ~v_448 | ~v_314 | ~v_3376 | ~v_3375 | ~v_3288 | ~v_3374 | ~v_3373 | ~v_3285 | ~v_3428 | ~v_3427 | ~v_3426 | ~v_3425 | ~v_1442 | ~v_3282 | ~v_1441 | ~v_3281 | ~v_1290 | ~v_1440 | ~v_3280 | ~v_1439 | ~v_3279 | ~v_1287 | ~v_1518 | ~v_1517 | ~v_1516 | ~v_1515 | v_3449;
assign x_11948 = v_3448 | ~v_3445;
assign x_11949 = v_3448 | ~v_3446;
assign x_11950 = v_3448 | ~v_3447;
assign x_11951 = v_103 | v_96 | v_95 | v_93 | v_102 | v_171 | v_170 | v_160 | v_150 | v_149 | v_184 | v_181 | ~v_297 | ~v_296 | ~v_345 | ~v_344 | ~v_343 | ~v_342 | ~v_341 | ~v_340 | ~v_3318 | ~v_3315 | ~v_3370 | ~v_3369 | ~v_3368 | ~v_3367 | ~v_3438 | ~v_3437 | ~v_3436 | ~v_3435 | ~v_3312 | ~v_3311 | ~v_1340 | ~v_3310 | ~v_3309 | ~v_1337 | ~v_1536 | ~v_1535 | ~v_1534 | ~v_1533 | ~v_1432 | ~v_1431 | ~v_1430 | ~v_1429 | v_3447;
assign x_11952 = v_54 | v_53 | v_61 | v_51 | v_60 | v_144 | v_180 | v_159 | v_145 | v_167 | v_166 | v_183 | ~v_264 | ~v_263 | ~v_330 | ~v_329 | ~v_328 | ~v_327 | ~v_326 | ~v_325 | ~v_3303 | ~v_3300 | ~v_3365 | ~v_3364 | ~v_3363 | ~v_3362 | ~v_3433 | ~v_3432 | ~v_3431 | ~v_3430 | ~v_3297 | ~v_3296 | ~v_1315 | ~v_3295 | ~v_3294 | ~v_1312 | ~v_1527 | ~v_1526 | ~v_1525 | ~v_1524 | ~v_1423 | ~v_1422 | ~v_1421 | ~v_1420 | v_3446;
assign x_11953 = v_18 | v_17 | v_8 | v_11 | v_10 | v_136 | v_137 | v_179 | v_163 | v_162 | v_155 | v_182 | ~v_231 | ~v_230 | ~v_315 | ~v_314 | ~v_313 | ~v_312 | ~v_311 | ~v_310 | ~v_3288 | ~v_3285 | ~v_3360 | ~v_3359 | ~v_3358 | ~v_3357 | ~v_3428 | ~v_3427 | ~v_3426 | ~v_3425 | ~v_3282 | ~v_3281 | ~v_1290 | ~v_3280 | ~v_3279 | ~v_1287 | ~v_1518 | ~v_1517 | ~v_1516 | ~v_1515 | ~v_1414 | ~v_1413 | ~v_1412 | ~v_1411 | v_3445;
assign x_11954 = v_3444 | ~v_3441;
assign x_11955 = v_3444 | ~v_3442;
assign x_11956 = v_3444 | ~v_3443;
assign x_11957 = v_103 | v_101 | v_93 | v_102 | v_171 | v_170 | v_150 | v_149 | v_148 | v_147 | v_184 | v_181 | ~v_391 | ~v_390 | ~v_387 | ~v_386 | ~v_345 | ~v_344 | ~v_385 | ~v_384 | ~v_3318 | ~v_3315 | ~v_3354 | ~v_3353 | ~v_3352 | ~v_3351 | ~v_3438 | ~v_3437 | ~v_3436 | ~v_3435 | ~v_3312 | ~v_3311 | ~v_1340 | ~v_3310 | ~v_3309 | ~v_1337 | ~v_1536 | ~v_1535 | ~v_1534 | ~v_1533 | ~v_1404 | ~v_1403 | ~v_1402 | ~v_1401 | v_3443;
assign x_11958 = v_61 | v_51 | v_60 | v_59 | v_144 | v_180 | v_145 | v_143 | v_142 | v_167 | v_166 | v_183 | ~v_376 | ~v_375 | ~v_372 | ~v_371 | ~v_330 | ~v_329 | ~v_370 | ~v_369 | ~v_3303 | ~v_3300 | ~v_3349 | ~v_3348 | ~v_3347 | ~v_3346 | ~v_3433 | ~v_3432 | ~v_3431 | ~v_3430 | ~v_3297 | ~v_3296 | ~v_1315 | ~v_3295 | ~v_3294 | ~v_1312 | ~v_1527 | ~v_1526 | ~v_1525 | ~v_1524 | ~v_1395 | ~v_1394 | ~v_1393 | ~v_1392 | v_3442;
assign x_11959 = v_18 | v_17 | v_16 | v_8 | v_136 | v_135 | v_134 | v_137 | v_179 | v_163 | v_162 | v_182 | ~v_361 | ~v_360 | ~v_357 | ~v_356 | ~v_315 | ~v_314 | ~v_355 | ~v_354 | ~v_3288 | ~v_3285 | ~v_3344 | ~v_3343 | ~v_3342 | ~v_3341 | ~v_3428 | ~v_3427 | ~v_3426 | ~v_3425 | ~v_3282 | ~v_3281 | ~v_1290 | ~v_3280 | ~v_3279 | ~v_1287 | ~v_1518 | ~v_1517 | ~v_1516 | ~v_1515 | ~v_1386 | ~v_1385 | ~v_1384 | ~v_1383 | v_3441;
assign x_11960 = v_3440 | ~v_3429;
assign x_11961 = v_3440 | ~v_3434;
assign x_11962 = v_3440 | ~v_3439;
assign x_11963 = v_101 | v_93 | v_102 | v_172 | v_171 | v_170 | v_150 | v_149 | v_148 | v_147 | v_184 | v_181 | ~v_3322 | ~v_3321 | ~v_437 | ~v_436 | ~v_435 | ~v_434 | ~v_345 | ~v_344 | ~v_433 | ~v_432 | ~v_3318 | ~v_3315 | ~v_3314 | ~v_3313 | ~v_3438 | ~v_3437 | ~v_3436 | ~v_3435 | ~v_3312 | ~v_3311 | ~v_1340 | ~v_3310 | ~v_3309 | ~v_1337 | ~v_1536 | ~v_1535 | ~v_1534 | ~v_1533 | ~v_1336 | ~v_1335 | ~v_1334 | ~v_1333 | v_3439;
assign x_11964 = v_3438 | v_157;
assign x_11965 = v_3438 | v_128;
assign x_11966 = v_3437 | v_156;
assign x_11967 = v_3437 | v_125;
assign x_11968 = v_3436 | ~v_157;
assign x_11969 = v_3436 | v_113;
assign x_11970 = v_3435 | ~v_156;
assign x_11971 = v_3435 | v_110;
assign x_11972 = v_51 | v_60 | v_59 | v_144 | v_180 | v_145 | v_143 | v_142 | v_168 | v_167 | v_166 | v_183 | ~v_3307 | ~v_3306 | ~v_422 | ~v_421 | ~v_420 | ~v_419 | ~v_330 | ~v_329 | ~v_418 | ~v_417 | ~v_3303 | ~v_3300 | ~v_3299 | ~v_3298 | ~v_3433 | ~v_3432 | ~v_3431 | ~v_3430 | ~v_3297 | ~v_3296 | ~v_1315 | ~v_3295 | ~v_3294 | ~v_1312 | ~v_1527 | ~v_1526 | ~v_1525 | ~v_1524 | ~v_1311 | ~v_1310 | ~v_1309 | ~v_1308 | v_3434;
assign x_11973 = v_3433 | v_157;
assign x_11974 = v_3433 | v_86;
assign x_11975 = v_3432 | v_156;
assign x_11976 = v_3432 | v_83;
assign x_11977 = v_3431 | ~v_157;
assign x_11978 = v_3431 | v_71;
assign x_11979 = v_3430 | ~v_156;
assign x_11980 = v_3430 | v_68;
assign x_11981 = v_17 | v_16 | v_8 | v_136 | v_135 | v_134 | v_137 | v_179 | v_164 | v_163 | v_162 | v_182 | ~v_3291 | ~v_3290 | ~v_407 | ~v_406 | ~v_405 | ~v_404 | ~v_315 | ~v_314 | ~v_403 | ~v_402 | ~v_3288 | ~v_3285 | ~v_3284 | ~v_3283 | ~v_3428 | ~v_3427 | ~v_3426 | ~v_3425 | ~v_3282 | ~v_3281 | ~v_1290 | ~v_3280 | ~v_3279 | ~v_1287 | ~v_1518 | ~v_1517 | ~v_1516 | ~v_1515 | ~v_1286 | ~v_1285 | ~v_1284 | ~v_1283 | v_3429;
assign x_11982 = v_3428 | v_157;
assign x_11983 = v_3428 | v_44;
assign x_11984 = v_3427 | v_156;
assign x_11985 = v_3427 | v_41;
assign x_11986 = v_3426 | ~v_157;
assign x_11987 = v_3426 | v_29;
assign x_11988 = v_3425 | ~v_156;
assign x_11989 = v_3425 | v_26;
assign x_11990 = v_3424 | ~v_3421;
assign x_11991 = v_3424 | ~v_3422;
assign x_11992 = v_3424 | ~v_3423;
assign x_11993 = v_98 | v_103 | v_96 | v_100 | v_94 | v_102 | v_169 | v_160 | v_150 | v_149 | v_147 | v_184 | ~v_299 | ~v_298 | ~v_297 | ~v_296 | ~v_295 | ~v_294 | ~v_293 | ~v_292 | ~v_3320 | ~v_3319 | ~v_3318 | ~v_3317 | ~v_3316 | ~v_3315 | ~v_3370 | ~v_3369 | ~v_3368 | ~v_3367 | ~v_1342 | ~v_3312 | ~v_1341 | ~v_3311 | ~v_1340 | ~v_1339 | ~v_3310 | ~v_1338 | ~v_3309 | ~v_1337 | ~v_1432 | ~v_1431 | ~v_1430 | ~v_1429 | v_3423;
assign x_11994 = v_54 | v_56 | v_61 | v_52 | v_60 | v_58 | v_144 | v_159 | v_145 | v_142 | v_165 | v_183 | ~v_3305 | ~v_266 | ~v_265 | ~v_264 | ~v_263 | ~v_262 | ~v_261 | ~v_260 | ~v_259 | ~v_3304 | ~v_3303 | ~v_3302 | ~v_3301 | ~v_3300 | ~v_3365 | ~v_3364 | ~v_3363 | ~v_3362 | ~v_1317 | ~v_3297 | ~v_1316 | ~v_3296 | ~v_1315 | ~v_1314 | ~v_3295 | ~v_1313 | ~v_3294 | ~v_1312 | ~v_1423 | ~v_1422 | ~v_1421 | ~v_1420 | v_3422;
assign x_11995 = v_13 | v_9 | v_18 | v_17 | v_15 | v_11 | v_136 | v_134 | ~v_3292 | v_137 | v_161 | v_155 | v_182 | ~v_233 | ~v_232 | ~v_231 | ~v_230 | ~v_229 | ~v_228 | ~v_227 | ~v_226 | ~v_3289 | ~v_3288 | ~v_3287 | ~v_3286 | ~v_3285 | ~v_3360 | ~v_3359 | ~v_3358 | ~v_3357 | ~v_1292 | ~v_3282 | ~v_1291 | ~v_3281 | ~v_1290 | ~v_1289 | ~v_3280 | ~v_1288 | ~v_3279 | ~v_1287 | ~v_1414 | ~v_1413 | ~v_1412 | ~v_1411 | v_3421;
assign x_11996 = v_3420 | ~v_3417;
assign x_11997 = v_3420 | ~v_3418;
assign x_11998 = v_3420 | ~v_3419;
assign x_11999 = v_101 | v_97 | v_100 | v_99 | v_102 | v_172 | v_171 | v_170 | v_169 | v_148 | v_147 | v_184 | ~v_483 | ~v_482 | ~v_593 | ~v_592 | ~v_545 | ~v_591 | ~v_590 | ~v_544 | ~v_3386 | ~v_3385 | ~v_3318 | ~v_3384 | ~v_3383 | ~v_3315 | ~v_3406 | ~v_3405 | ~v_3404 | ~v_3403 | ~v_1460 | ~v_3312 | ~v_1459 | ~v_3311 | ~v_1340 | ~v_1458 | ~v_3310 | ~v_1457 | ~v_3309 | ~v_1337 | ~v_1492 | ~v_1491 | ~v_1490 | ~v_1489 | v_3419;
assign x_12000 = v_55 | v_60 | v_59 | v_58 | v_57 | v_143 | v_142 | v_168 | v_167 | v_166 | v_165 | v_183 | ~v_3381 | ~v_3380 | ~v_468 | ~v_467 | ~v_588 | ~v_587 | ~v_530 | ~v_586 | ~v_585 | ~v_529 | ~v_3303 | ~v_3379 | ~v_3378 | ~v_3300 | ~v_3401 | ~v_3400 | ~v_3399 | ~v_3398 | ~v_1451 | ~v_3297 | ~v_1450 | ~v_3296 | ~v_1315 | ~v_1449 | ~v_3295 | ~v_1448 | ~v_3294 | ~v_1312 | ~v_1483 | ~v_1482 | ~v_1481 | ~v_1480 | v_3418;
assign x_12001 = v_17 | v_16 | v_15 | v_14 | v_12 | ~v_453 | ~v_452 | v_135 | v_134 | v_164 | v_163 | v_162 | v_161 | v_182 | ~v_583 | ~v_582 | ~v_515 | ~v_581 | ~v_580 | ~v_514 | ~v_3376 | ~v_3375 | ~v_3288 | ~v_3374 | ~v_3373 | ~v_3285 | ~v_3396 | ~v_3395 | ~v_3394 | ~v_3393 | ~v_1442 | ~v_3282 | ~v_1441 | ~v_3281 | ~v_1290 | ~v_1440 | ~v_3280 | ~v_1439 | ~v_3279 | ~v_1287 | ~v_1474 | ~v_1473 | ~v_1472 | ~v_1471 | v_3417;
assign x_12002 = v_3416 | ~v_3413;
assign x_12003 = v_3416 | ~v_3414;
assign x_12004 = v_3416 | ~v_3415;
assign x_12005 = v_103 | v_96 | v_100 | v_102 | v_171 | v_170 | v_169 | v_160 | v_150 | v_149 | v_147 | v_184 | ~v_545 | ~v_544 | ~v_543 | ~v_542 | ~v_541 | ~v_540 | ~v_297 | ~v_296 | ~v_3318 | ~v_3315 | ~v_3406 | ~v_3405 | ~v_3404 | ~v_3403 | ~v_3370 | ~v_3369 | ~v_3368 | ~v_3367 | ~v_3312 | ~v_3311 | ~v_1340 | ~v_3310 | ~v_3309 | ~v_1337 | ~v_1432 | ~v_1431 | ~v_1430 | ~v_1429 | ~v_1492 | ~v_1491 | ~v_1490 | ~v_1489 | v_3415;
assign x_12006 = v_54 | v_61 | v_60 | v_58 | v_144 | v_159 | v_145 | v_142 | v_167 | v_166 | v_165 | v_183 | ~v_530 | ~v_529 | ~v_528 | ~v_527 | ~v_526 | ~v_525 | ~v_264 | ~v_263 | ~v_3303 | ~v_3300 | ~v_3401 | ~v_3400 | ~v_3399 | ~v_3398 | ~v_3365 | ~v_3364 | ~v_3363 | ~v_3362 | ~v_3297 | ~v_3296 | ~v_1315 | ~v_3295 | ~v_3294 | ~v_1312 | ~v_1423 | ~v_1422 | ~v_1421 | ~v_1420 | ~v_1483 | ~v_1482 | ~v_1481 | ~v_1480 | v_3414;
assign x_12007 = v_18 | v_17 | v_15 | v_11 | v_136 | v_134 | v_137 | v_163 | v_162 | v_161 | v_155 | v_182 | ~v_515 | ~v_514 | ~v_513 | ~v_512 | ~v_511 | ~v_510 | ~v_231 | ~v_230 | ~v_3288 | ~v_3285 | ~v_3396 | ~v_3395 | ~v_3394 | ~v_3393 | ~v_3360 | ~v_3359 | ~v_3358 | ~v_3357 | ~v_3282 | ~v_3281 | ~v_1290 | ~v_3280 | ~v_3279 | ~v_1287 | ~v_1414 | ~v_1413 | ~v_1412 | ~v_1411 | ~v_1474 | ~v_1473 | ~v_1472 | ~v_1471 | v_3413;
assign x_12008 = v_3412 | ~v_3409;
assign x_12009 = v_3412 | ~v_3410;
assign x_12010 = v_3412 | ~v_3411;
assign x_12011 = v_103 | v_101 | v_100 | v_95 | v_102 | v_171 | v_170 | v_169 | v_150 | v_149 | v_148 | v_184 | ~v_545 | ~v_544 | ~v_561 | ~v_560 | ~v_559 | ~v_558 | ~v_387 | ~v_386 | ~v_3318 | ~v_3315 | ~v_3406 | ~v_3405 | ~v_3404 | ~v_3403 | ~v_3354 | ~v_3353 | ~v_3352 | ~v_3351 | ~v_3312 | ~v_3311 | ~v_1340 | ~v_3310 | ~v_3309 | ~v_1337 | ~v_1404 | ~v_1403 | ~v_1402 | ~v_1401 | ~v_1492 | ~v_1491 | ~v_1490 | ~v_1489 | v_3411;
assign x_12012 = v_53 | v_61 | v_60 | v_59 | v_58 | v_144 | v_145 | v_143 | v_167 | v_166 | v_165 | v_183 | ~v_530 | ~v_529 | ~v_556 | ~v_555 | ~v_554 | ~v_553 | ~v_372 | ~v_371 | ~v_3303 | ~v_3300 | ~v_3401 | ~v_3400 | ~v_3399 | ~v_3398 | ~v_3349 | ~v_3348 | ~v_3347 | ~v_3346 | ~v_3297 | ~v_3296 | ~v_1315 | ~v_3295 | ~v_3294 | ~v_1312 | ~v_1395 | ~v_1394 | ~v_1393 | ~v_1392 | ~v_1483 | ~v_1482 | ~v_1481 | ~v_1480 | v_3410;
assign x_12013 = v_18 | v_17 | v_16 | v_15 | v_10 | v_136 | v_135 | v_137 | v_163 | v_162 | v_161 | v_182 | ~v_515 | ~v_514 | ~v_551 | ~v_550 | ~v_549 | ~v_548 | ~v_357 | ~v_356 | ~v_3288 | ~v_3285 | ~v_3396 | ~v_3395 | ~v_3394 | ~v_3393 | ~v_3344 | ~v_3343 | ~v_3342 | ~v_3341 | ~v_3282 | ~v_3281 | ~v_1290 | ~v_3280 | ~v_3279 | ~v_1287 | ~v_1386 | ~v_1385 | ~v_1384 | ~v_1383 | ~v_1474 | ~v_1473 | ~v_1472 | ~v_1471 | v_3409;
assign x_12014 = v_3408 | ~v_3397;
assign x_12015 = v_3408 | ~v_3402;
assign x_12016 = v_3408 | ~v_3407;
assign x_12017 = v_103 | v_101 | v_100 | v_151 | v_171 | v_170 | v_169 | v_150 | v_149 | v_148 | v_147 | v_184 | ~v_3322 | ~v_3321 | ~v_577 | ~v_576 | ~v_545 | ~v_544 | ~v_575 | ~v_574 | ~v_435 | ~v_434 | ~v_3318 | ~v_3315 | ~v_3406 | ~v_3405 | ~v_3404 | ~v_3403 | ~v_3314 | ~v_3313 | ~v_3312 | ~v_3311 | ~v_1340 | ~v_3310 | ~v_3309 | ~v_1337 | ~v_1336 | ~v_1335 | ~v_1334 | ~v_1333 | ~v_1492 | ~v_1491 | ~v_1490 | ~v_1489 | v_3407;
assign x_12018 = v_3406 | v_140;
assign x_12019 = v_3406 | v_128;
assign x_12020 = v_3405 | v_139;
assign x_12021 = v_3405 | v_125;
assign x_12022 = v_3404 | ~v_140;
assign x_12023 = v_3404 | v_113;
assign x_12024 = v_3403 | ~v_139;
assign x_12025 = v_3403 | v_110;
assign x_12026 = v_61 | v_59 | v_58 | v_144 | v_145 | v_143 | v_142 | v_167 | v_166 | v_165 | v_146 | v_183 | ~v_3307 | ~v_3306 | ~v_572 | ~v_571 | ~v_530 | ~v_529 | ~v_570 | ~v_569 | ~v_420 | ~v_419 | ~v_3303 | ~v_3300 | ~v_3401 | ~v_3400 | ~v_3399 | ~v_3398 | ~v_3299 | ~v_3298 | ~v_3297 | ~v_3296 | ~v_1315 | ~v_3295 | ~v_3294 | ~v_1312 | ~v_1311 | ~v_1310 | ~v_1309 | ~v_1308 | ~v_1483 | ~v_1482 | ~v_1481 | ~v_1480 | v_3402;
assign x_12027 = v_3401 | v_140;
assign x_12028 = v_3401 | v_86;
assign x_12029 = v_3400 | v_139;
assign x_12030 = v_3400 | v_83;
assign x_12031 = v_3399 | ~v_140;
assign x_12032 = v_3399 | v_71;
assign x_12033 = v_3398 | ~v_139;
assign x_12034 = v_3398 | v_68;
assign x_12035 = v_18 | v_16 | v_15 | v_136 | v_135 | v_134 | v_137 | v_138 | v_163 | v_162 | v_161 | v_182 | ~v_3291 | ~v_3290 | ~v_567 | ~v_566 | ~v_515 | ~v_514 | ~v_565 | ~v_564 | ~v_405 | ~v_404 | ~v_3288 | ~v_3285 | ~v_3396 | ~v_3395 | ~v_3394 | ~v_3393 | ~v_3284 | ~v_3283 | ~v_3282 | ~v_3281 | ~v_1290 | ~v_3280 | ~v_3279 | ~v_1287 | ~v_1286 | ~v_1285 | ~v_1284 | ~v_1283 | ~v_1474 | ~v_1473 | ~v_1472 | ~v_1471 | v_3397;
assign x_12036 = v_3396 | v_140;
assign x_12037 = v_3396 | v_44;
assign x_12038 = v_3395 | v_139;
assign x_12039 = v_3395 | v_41;
assign x_12040 = v_3394 | ~v_140;
assign x_12041 = v_3394 | v_29;
assign x_12042 = v_3393 | ~v_139;
assign x_12043 = v_3393 | v_26;
assign x_12044 = v_3392 | ~v_3389;
assign x_12045 = v_3392 | ~v_3390;
assign x_12046 = v_3392 | ~v_3391;
assign x_12047 = v_98 | v_103 | v_101 | v_100 | v_94 | v_151 | v_169 | v_150 | v_149 | v_148 | v_147 | v_184 | ~v_299 | ~v_298 | ~v_387 | ~v_386 | ~v_499 | ~v_498 | ~v_497 | ~v_496 | ~v_3320 | ~v_3319 | ~v_3318 | ~v_3317 | ~v_3316 | ~v_3315 | ~v_3354 | ~v_3353 | ~v_3352 | ~v_3351 | ~v_1342 | ~v_3312 | ~v_1341 | ~v_3311 | ~v_1340 | ~v_1339 | ~v_3310 | ~v_1338 | ~v_3309 | ~v_1337 | ~v_1404 | ~v_1403 | ~v_1402 | ~v_1401 | v_3391;
assign x_12048 = v_56 | v_61 | v_52 | v_59 | v_58 | v_144 | v_145 | v_143 | v_142 | v_165 | v_146 | v_183 | ~v_3305 | ~v_266 | ~v_265 | ~v_372 | ~v_371 | ~v_494 | ~v_493 | ~v_492 | ~v_491 | ~v_3304 | ~v_3303 | ~v_3302 | ~v_3301 | ~v_3300 | ~v_3349 | ~v_3348 | ~v_3347 | ~v_3346 | ~v_1317 | ~v_3297 | ~v_1316 | ~v_3296 | ~v_1315 | ~v_1314 | ~v_3295 | ~v_1313 | ~v_3294 | ~v_1312 | ~v_1395 | ~v_1394 | ~v_1393 | ~v_1392 | v_3390;
assign x_12049 = v_13 | v_9 | v_18 | v_16 | v_15 | v_136 | v_135 | v_134 | ~v_3292 | v_137 | v_138 | v_161 | v_182 | ~v_233 | ~v_232 | ~v_357 | ~v_356 | ~v_489 | ~v_488 | ~v_487 | ~v_486 | ~v_3289 | ~v_3288 | ~v_3287 | ~v_3286 | ~v_3285 | ~v_3344 | ~v_3343 | ~v_3342 | ~v_3341 | ~v_1292 | ~v_3282 | ~v_1291 | ~v_3281 | ~v_1290 | ~v_1289 | ~v_3280 | ~v_1288 | ~v_3279 | ~v_1287 | ~v_1386 | ~v_1385 | ~v_1384 | ~v_1383 | v_3389;
assign x_12050 = v_3388 | ~v_3377;
assign x_12051 = v_3388 | ~v_3382;
assign x_12052 = v_3388 | ~v_3387;
assign x_12053 = v_103 | v_101 | v_97 | v_100 | v_99 | v_102 | v_171 | v_170 | v_169 | v_148 | v_147 | v_184 | ~v_703 | ~v_702 | ~v_483 | ~v_482 | ~v_701 | ~v_653 | ~v_700 | ~v_652 | ~v_3386 | ~v_3385 | ~v_3318 | ~v_3384 | ~v_3383 | ~v_3315 | ~v_3338 | ~v_3337 | ~v_3336 | ~v_3335 | ~v_1460 | ~v_3312 | ~v_1459 | ~v_3311 | ~v_1340 | ~v_1458 | ~v_3310 | ~v_1457 | ~v_3309 | ~v_1337 | ~v_1376 | ~v_1375 | ~v_1374 | ~v_1373 | v_3387;
assign x_12054 = v_3386 | v_131;
assign x_12055 = v_3386 | v_19;
assign x_12056 = v_3385 | v_126;
assign x_12057 = v_3385 | v_19;
assign x_12058 = v_3384 | v_116;
assign x_12059 = v_3384 | ~v_19;
assign x_12060 = v_3383 | v_111;
assign x_12061 = v_3383 | ~v_19;
assign x_12062 = v_55 | v_61 | v_60 | v_59 | v_58 | v_57 | v_143 | v_142 | v_167 | v_166 | v_165 | v_183 | ~v_698 | ~v_697 | ~v_3381 | ~v_3380 | ~v_468 | ~v_467 | ~v_696 | ~v_638 | ~v_695 | ~v_637 | ~v_3303 | ~v_3379 | ~v_3378 | ~v_3300 | ~v_3333 | ~v_3332 | ~v_3331 | ~v_3330 | ~v_1451 | ~v_3297 | ~v_1450 | ~v_3296 | ~v_1315 | ~v_1449 | ~v_3295 | ~v_1448 | ~v_3294 | ~v_1312 | ~v_1367 | ~v_1366 | ~v_1365 | ~v_1364 | v_3382;
assign x_12063 = v_3381 | v_84;
assign x_12064 = v_3381 | v_19;
assign x_12065 = v_3380 | v_89;
assign x_12066 = v_3380 | v_19;
assign x_12067 = v_3379 | v_74;
assign x_12068 = v_3379 | ~v_19;
assign x_12069 = v_3378 | v_69;
assign x_12070 = v_3378 | ~v_19;
assign x_12071 = v_18 | v_17 | v_16 | v_15 | v_14 | v_12 | ~v_453 | ~v_452 | v_135 | v_134 | v_163 | v_162 | v_161 | v_182 | ~v_693 | ~v_692 | ~v_691 | ~v_623 | ~v_690 | ~v_622 | ~v_3376 | ~v_3375 | ~v_3288 | ~v_3374 | ~v_3373 | ~v_3285 | ~v_3328 | ~v_3327 | ~v_3326 | ~v_3325 | ~v_1442 | ~v_3282 | ~v_1441 | ~v_3281 | ~v_1290 | ~v_1440 | ~v_3280 | ~v_1439 | ~v_3279 | ~v_1287 | ~v_1358 | ~v_1357 | ~v_1356 | ~v_1355 | v_3377;
assign x_12072 = v_3376 | v_47;
assign x_12073 = v_3376 | v_19;
assign x_12074 = v_3375 | v_42;
assign x_12075 = v_3375 | v_19;
assign x_12076 = v_3374 | v_32;
assign x_12077 = v_3374 | ~v_19;
assign x_12078 = v_3373 | v_27;
assign x_12079 = v_3373 | ~v_19;
assign x_12080 = v_3372 | ~v_3361;
assign x_12081 = v_3372 | ~v_3366;
assign x_12082 = v_3372 | ~v_3371;
assign x_12083 = v_103 | v_96 | v_100 | v_151 | v_171 | v_170 | v_169 | v_160 | v_150 | v_149 | v_147 | v_184 | ~v_655 | ~v_654 | ~v_297 | ~v_296 | ~v_653 | ~v_652 | ~v_651 | ~v_650 | ~v_3318 | ~v_3315 | ~v_3370 | ~v_3369 | ~v_3368 | ~v_3367 | ~v_3338 | ~v_3337 | ~v_3336 | ~v_3335 | ~v_3312 | ~v_3311 | ~v_1340 | ~v_3310 | ~v_3309 | ~v_1337 | ~v_1432 | ~v_1431 | ~v_1430 | ~v_1429 | ~v_1376 | ~v_1375 | ~v_1374 | ~v_1373 | v_3371;
assign x_12084 = v_3370 | v_157;
assign x_12085 = v_3370 | v_131;
assign x_12086 = v_3369 | v_156;
assign x_12087 = v_3369 | v_126;
assign x_12088 = v_3368 | ~v_157;
assign x_12089 = v_3368 | v_116;
assign x_12090 = v_3367 | ~v_156;
assign x_12091 = v_3367 | v_111;
assign x_12092 = v_54 | v_61 | v_58 | v_144 | v_159 | v_145 | v_142 | v_167 | v_166 | v_165 | v_146 | v_183 | ~v_640 | ~v_639 | ~v_264 | ~v_263 | ~v_638 | ~v_637 | ~v_636 | ~v_635 | ~v_3303 | ~v_3300 | ~v_3365 | ~v_3364 | ~v_3363 | ~v_3362 | ~v_3333 | ~v_3332 | ~v_3331 | ~v_3330 | ~v_3297 | ~v_3296 | ~v_1315 | ~v_3295 | ~v_3294 | ~v_1312 | ~v_1423 | ~v_1422 | ~v_1421 | ~v_1420 | ~v_1367 | ~v_1366 | ~v_1365 | ~v_1364 | v_3366;
assign x_12093 = v_3365 | v_157;
assign x_12094 = v_3365 | v_89;
assign x_12095 = v_3364 | v_156;
assign x_12096 = v_3364 | v_84;
assign x_12097 = v_3363 | ~v_157;
assign x_12098 = v_3363 | v_74;
assign x_12099 = v_3362 | ~v_156;
assign x_12100 = v_3362 | v_69;
assign x_12101 = v_18 | v_15 | v_11 | v_136 | v_134 | v_137 | v_138 | v_163 | v_162 | v_161 | v_155 | v_182 | ~v_625 | ~v_624 | ~v_231 | ~v_230 | ~v_623 | ~v_622 | ~v_621 | ~v_620 | ~v_3288 | ~v_3285 | ~v_3360 | ~v_3359 | ~v_3358 | ~v_3357 | ~v_3328 | ~v_3327 | ~v_3326 | ~v_3325 | ~v_3282 | ~v_3281 | ~v_1290 | ~v_3280 | ~v_3279 | ~v_1287 | ~v_1414 | ~v_1413 | ~v_1412 | ~v_1411 | ~v_1358 | ~v_1357 | ~v_1356 | ~v_1355 | v_3361;
assign x_12102 = v_3360 | v_157;
assign x_12103 = v_3360 | v_47;
assign x_12104 = v_3359 | v_156;
assign x_12105 = v_3359 | v_42;
assign x_12106 = v_3358 | ~v_157;
assign x_12107 = v_3358 | v_32;
assign x_12108 = v_3357 | ~v_156;
assign x_12109 = v_3357 | v_27;
assign x_12110 = v_3356 | ~v_3345;
assign x_12111 = v_3356 | ~v_3350;
assign x_12112 = v_3356 | ~v_3355;
assign x_12113 = v_101 | v_100 | v_102 | v_172 | v_171 | v_170 | v_169 | v_150 | v_149 | v_148 | v_147 | v_184 | ~v_671 | ~v_670 | ~v_387 | ~v_386 | ~v_653 | ~v_652 | ~v_669 | ~v_668 | ~v_3318 | ~v_3315 | ~v_3354 | ~v_3353 | ~v_3352 | ~v_3351 | ~v_3338 | ~v_3337 | ~v_3336 | ~v_3335 | ~v_3312 | ~v_3311 | ~v_1340 | ~v_3310 | ~v_3309 | ~v_1337 | ~v_1404 | ~v_1403 | ~v_1402 | ~v_1401 | ~v_1376 | ~v_1375 | ~v_1374 | ~v_1373 | v_3355;
assign x_12114 = v_3354 | v_140;
assign x_12115 = v_3354 | v_131;
assign x_12116 = v_3353 | v_139;
assign x_12117 = v_3353 | v_126;
assign x_12118 = v_3352 | ~v_140;
assign x_12119 = v_3352 | v_116;
assign x_12120 = v_3351 | ~v_139;
assign x_12121 = v_3351 | v_111;
assign x_12122 = v_60 | v_59 | v_58 | v_144 | v_145 | v_143 | v_142 | v_168 | v_167 | v_166 | v_165 | v_183 | ~v_666 | ~v_665 | ~v_372 | ~v_371 | ~v_638 | ~v_637 | ~v_664 | ~v_663 | ~v_3303 | ~v_3300 | ~v_3349 | ~v_3348 | ~v_3347 | ~v_3346 | ~v_3333 | ~v_3332 | ~v_3331 | ~v_3330 | ~v_3297 | ~v_3296 | ~v_1315 | ~v_3295 | ~v_3294 | ~v_1312 | ~v_1395 | ~v_1394 | ~v_1393 | ~v_1392 | ~v_1367 | ~v_1366 | ~v_1365 | ~v_1364 | v_3350;
assign x_12123 = v_3349 | v_140;
assign x_12124 = v_3349 | v_89;
assign x_12125 = v_3348 | v_139;
assign x_12126 = v_3348 | v_84;
assign x_12127 = v_3347 | ~v_140;
assign x_12128 = v_3347 | v_74;
assign x_12129 = v_3346 | ~v_139;
assign x_12130 = v_3346 | v_69;
assign x_12131 = v_17 | v_16 | v_15 | v_136 | v_135 | v_134 | v_137 | v_164 | v_163 | v_162 | v_161 | v_182 | ~v_661 | ~v_660 | ~v_357 | ~v_356 | ~v_623 | ~v_622 | ~v_659 | ~v_658 | ~v_3288 | ~v_3285 | ~v_3344 | ~v_3343 | ~v_3342 | ~v_3341 | ~v_3328 | ~v_3327 | ~v_3326 | ~v_3325 | ~v_3282 | ~v_3281 | ~v_1290 | ~v_3280 | ~v_3279 | ~v_1287 | ~v_1386 | ~v_1385 | ~v_1384 | ~v_1383 | ~v_1358 | ~v_1357 | ~v_1356 | ~v_1355 | v_3345;
assign x_12132 = v_3344 | v_140;
assign x_12133 = v_3344 | v_47;
assign x_12134 = v_3343 | v_139;
assign x_12135 = v_3343 | v_42;
assign x_12136 = v_3342 | ~v_140;
assign x_12137 = v_3342 | v_32;
assign x_12138 = v_3341 | ~v_139;
assign x_12139 = v_3341 | v_27;
assign x_12140 = v_3340 | ~v_3329;
assign x_12141 = v_3340 | ~v_3334;
assign x_12142 = v_3340 | ~v_3339;
assign x_12143 = v_103 | v_101 | v_100 | v_95 | v_102 | v_171 | v_170 | v_169 | v_150 | v_149 | v_148 | v_184 | ~v_3322 | ~v_3321 | ~v_435 | ~v_434 | ~v_653 | ~v_652 | ~v_687 | ~v_686 | ~v_685 | ~v_684 | ~v_3318 | ~v_3315 | ~v_3314 | ~v_3313 | ~v_3338 | ~v_3337 | ~v_3336 | ~v_3335 | ~v_3312 | ~v_3311 | ~v_1340 | ~v_3310 | ~v_3309 | ~v_1337 | ~v_1336 | ~v_1335 | ~v_1334 | ~v_1333 | ~v_1376 | ~v_1375 | ~v_1374 | ~v_1373 | v_3339;
assign x_12144 = v_3338 | v_153;
assign x_12145 = v_3338 | v_128;
assign x_12146 = v_3337 | v_152;
assign x_12147 = v_3337 | v_125;
assign x_12148 = v_3336 | ~v_153;
assign x_12149 = v_3336 | v_113;
assign x_12150 = v_3335 | ~v_152;
assign x_12151 = v_3335 | v_110;
assign x_12152 = v_53 | v_61 | v_60 | v_59 | v_58 | v_144 | v_145 | v_143 | v_167 | v_166 | v_165 | v_183 | ~v_3307 | ~v_3306 | ~v_420 | ~v_419 | ~v_638 | ~v_637 | ~v_682 | ~v_681 | ~v_680 | ~v_679 | ~v_3303 | ~v_3300 | ~v_3299 | ~v_3298 | ~v_3333 | ~v_3332 | ~v_3331 | ~v_3330 | ~v_3297 | ~v_3296 | ~v_1315 | ~v_3295 | ~v_3294 | ~v_1312 | ~v_1311 | ~v_1310 | ~v_1309 | ~v_1308 | ~v_1367 | ~v_1366 | ~v_1365 | ~v_1364 | v_3334;
assign x_12153 = v_3333 | v_153;
assign x_12154 = v_3333 | v_86;
assign x_12155 = v_3332 | v_152;
assign x_12156 = v_3332 | v_83;
assign x_12157 = v_3331 | ~v_153;
assign x_12158 = v_3331 | v_71;
assign x_12159 = v_3330 | ~v_152;
assign x_12160 = v_3330 | v_68;
assign x_12161 = v_18 | v_17 | v_16 | v_15 | v_10 | v_136 | v_135 | v_137 | v_163 | v_162 | v_161 | v_182 | ~v_3291 | ~v_3290 | ~v_405 | ~v_404 | ~v_623 | ~v_622 | ~v_677 | ~v_676 | ~v_675 | ~v_674 | ~v_3288 | ~v_3285 | ~v_3284 | ~v_3283 | ~v_3328 | ~v_3327 | ~v_3326 | ~v_3325 | ~v_3282 | ~v_3281 | ~v_1290 | ~v_3280 | ~v_3279 | ~v_1287 | ~v_1286 | ~v_1285 | ~v_1284 | ~v_1283 | ~v_1358 | ~v_1357 | ~v_1356 | ~v_1355 | v_3329;
assign x_12162 = v_3328 | v_153;
assign x_12163 = v_3328 | v_44;
assign x_12164 = v_3327 | v_152;
assign x_12165 = v_3327 | v_41;
assign x_12166 = v_3326 | ~v_153;
assign x_12167 = v_3326 | v_29;
assign x_12168 = v_3325 | ~v_152;
assign x_12169 = v_3325 | v_26;
assign x_12170 = v_3324 | ~v_3293;
assign x_12171 = v_3324 | ~v_3308;
assign x_12172 = v_3324 | ~v_3323;
assign x_12173 = v_98 | v_103 | v_101 | v_100 | v_94 | v_102 | v_169 | v_150 | v_149 | v_148 | v_147 | v_184 | ~v_609 | ~v_608 | ~v_3322 | ~v_3321 | ~v_299 | ~v_298 | ~v_435 | ~v_434 | ~v_607 | ~v_606 | ~v_3320 | ~v_3319 | ~v_3318 | ~v_3317 | ~v_3316 | ~v_3315 | ~v_3314 | ~v_3313 | ~v_1342 | ~v_3312 | ~v_1341 | ~v_3311 | ~v_1340 | ~v_1339 | ~v_3310 | ~v_1338 | ~v_3309 | ~v_1337 | ~v_1336 | ~v_1335 | ~v_1334 | ~v_1333 | v_3323;
assign x_12174 = v_3322 | v_153;
assign x_12175 = v_3322 | v_131;
assign x_12176 = v_3321 | ~v_153;
assign x_12177 = v_3321 | v_116;
assign x_12178 = v_3320 | v_128;
assign x_12179 = v_3320 | v_19;
assign x_12180 = v_3319 | v_125;
assign x_12181 = v_3319 | v_19;
assign x_12182 = v_3318 | v_124;
assign x_12183 = v_3318 | v_19;
assign x_12184 = v_3317 | v_113;
assign x_12185 = v_3317 | ~v_19;
assign x_12186 = v_3316 | v_110;
assign x_12187 = v_3316 | ~v_19;
assign x_12188 = v_3315 | v_109;
assign x_12189 = v_3315 | ~v_19;
assign x_12190 = v_3314 | v_152;
assign x_12191 = v_3314 | v_126;
assign x_12192 = v_3313 | ~v_152;
assign x_12193 = v_3313 | v_111;
assign x_12194 = v_3312 | v_156;
assign x_12195 = v_3312 | v_123;
assign x_12196 = v_3311 | v_157;
assign x_12197 = v_3311 | v_120;
assign x_12198 = v_3310 | ~v_156;
assign x_12199 = v_3310 | v_108;
assign x_12200 = v_3309 | ~v_157;
assign x_12201 = v_3309 | v_105;
assign x_12202 = v_56 | v_61 | v_52 | v_60 | v_59 | v_58 | v_144 | v_145 | v_143 | v_142 | v_165 | v_183 | ~v_604 | ~v_603 | ~v_3307 | ~v_3306 | ~v_3305 | ~v_266 | ~v_265 | ~v_420 | ~v_419 | ~v_602 | ~v_601 | ~v_3304 | ~v_3303 | ~v_3302 | ~v_3301 | ~v_3300 | ~v_3299 | ~v_3298 | ~v_1317 | ~v_3297 | ~v_1316 | ~v_3296 | ~v_1315 | ~v_1314 | ~v_3295 | ~v_1313 | ~v_3294 | ~v_1312 | ~v_1311 | ~v_1310 | ~v_1309 | ~v_1308 | v_3308;
assign x_12203 = v_3307 | v_153;
assign x_12204 = v_3307 | v_89;
assign x_12205 = v_3306 | ~v_153;
assign x_12206 = v_3306 | v_74;
assign x_12207 = v_3305 | v_83;
assign x_12208 = v_3305 | v_19;
assign x_12209 = v_3304 | v_86;
assign x_12210 = v_3304 | v_19;
assign x_12211 = v_3303 | v_82;
assign x_12212 = v_3303 | v_19;
assign x_12213 = v_3302 | v_71;
assign x_12214 = v_3302 | ~v_19;
assign x_12215 = v_3301 | v_68;
assign x_12216 = v_3301 | ~v_19;
assign x_12217 = v_3300 | v_67;
assign x_12218 = v_3300 | ~v_19;
assign x_12219 = v_3299 | v_152;
assign x_12220 = v_3299 | v_84;
assign x_12221 = v_3298 | ~v_152;
assign x_12222 = v_3298 | v_69;
assign x_12223 = v_3297 | v_156;
assign x_12224 = v_3297 | v_81;
assign x_12225 = v_3296 | v_157;
assign x_12226 = v_3296 | v_78;
assign x_12227 = v_3295 | ~v_156;
assign x_12228 = v_3295 | v_66;
assign x_12229 = v_3294 | ~v_157;
assign x_12230 = v_3294 | v_63;
assign x_12231 = v_13 | v_9 | v_18 | v_17 | v_16 | v_15 | v_136 | v_135 | v_134 | ~v_3292 | v_137 | v_161 | v_182 | ~v_599 | ~v_598 | ~v_3291 | ~v_3290 | ~v_233 | ~v_232 | ~v_405 | ~v_404 | ~v_597 | ~v_596 | ~v_3289 | ~v_3288 | ~v_3287 | ~v_3286 | ~v_3285 | ~v_3284 | ~v_3283 | ~v_1292 | ~v_3282 | ~v_1291 | ~v_3281 | ~v_1290 | ~v_1289 | ~v_3280 | ~v_1288 | ~v_3279 | ~v_1287 | ~v_1286 | ~v_1285 | ~v_1284 | ~v_1283 | v_3293;
assign x_12232 = v_3292 | v_41;
assign x_12233 = v_3292 | v_19;
assign x_12234 = v_3291 | v_153;
assign x_12235 = v_3291 | v_47;
assign x_12236 = v_3290 | ~v_153;
assign x_12237 = v_3290 | v_32;
assign x_12238 = v_3289 | v_44;
assign x_12239 = v_3289 | v_19;
assign x_12240 = v_3288 | v_40;
assign x_12241 = v_3288 | v_19;
assign x_12242 = v_3287 | v_29;
assign x_12243 = v_3287 | ~v_19;
assign x_12244 = v_3286 | v_26;
assign x_12245 = v_3286 | ~v_19;
assign x_12246 = v_3285 | v_25;
assign x_12247 = v_3285 | ~v_19;
assign x_12248 = v_3284 | v_152;
assign x_12249 = v_3284 | v_42;
assign x_12250 = v_3283 | ~v_152;
assign x_12251 = v_3283 | v_27;
assign x_12252 = v_3282 | v_156;
assign x_12253 = v_3282 | v_39;
assign x_12254 = v_3281 | v_157;
assign x_12255 = v_3281 | v_36;
assign x_12256 = v_3280 | ~v_156;
assign x_12257 = v_3280 | v_24;
assign x_12258 = v_3279 | ~v_157;
assign x_12259 = v_3279 | v_21;
assign x_12260 = v_3278 | ~v_3276;
assign x_12261 = v_3278 | ~v_3277;
assign x_12262 = v_3278 | ~v_194;
assign x_12263 = v_3278 | ~v_196;
assign x_12264 = v_3278 | ~v_157;
assign x_12265 = v_3278 | ~v_156;
assign x_12266 = ~v_195 | ~v_2221 | v_3277;
assign x_12267 = ~v_188 | ~v_1276 | v_3276;
assign x_12268 = v_3275 | ~v_3092;
assign x_12269 = v_3275 | ~v_3274;
assign x_12270 = v_157 | v_156 | ~v_3273 | ~v_738 | ~v_736 | ~v_3094 | ~v_3093 | v_3274;
assign x_12271 = v_3273 | ~v_3140;
assign x_12272 = v_3273 | ~v_3156;
assign x_12273 = v_3273 | ~v_3172;
assign x_12274 = v_3273 | ~v_3188;
assign x_12275 = v_3273 | ~v_3204;
assign x_12276 = v_3273 | ~v_3208;
assign x_12277 = v_3273 | ~v_3224;
assign x_12278 = v_3273 | ~v_3228;
assign x_12279 = v_3273 | ~v_3232;
assign x_12280 = v_3273 | ~v_3236;
assign x_12281 = v_3273 | ~v_3240;
assign x_12282 = v_3273 | ~v_3256;
assign x_12283 = v_3273 | ~v_3260;
assign x_12284 = v_3273 | ~v_3264;
assign x_12285 = v_3273 | ~v_3268;
assign x_12286 = v_3273 | ~v_3272;
assign x_12287 = v_3273 | ~v_1263;
assign x_12288 = v_3273 | ~v_1264;
assign x_12289 = v_3273 | ~v_1265;
assign x_12290 = v_3273 | ~v_1266;
assign x_12291 = ~v_3271 | ~v_3270 | ~v_3269 | v_3272;
assign x_12292 = v_3271 | ~v_3125;
assign x_12293 = v_3271 | ~v_3126;
assign x_12294 = v_3271 | ~v_817;
assign x_12295 = v_3271 | ~v_818;
assign x_12296 = v_3271 | ~v_1011;
assign x_12297 = v_3271 | ~v_819;
assign x_12298 = v_3271 | ~v_1012;
assign x_12299 = v_3271 | ~v_3127;
assign x_12300 = v_3271 | ~v_3128;
assign x_12301 = v_3271 | ~v_820;
assign x_12302 = v_3271 | ~v_821;
assign x_12303 = v_3271 | ~v_1013;
assign x_12304 = v_3271 | ~v_822;
assign x_12305 = v_3271 | ~v_1014;
assign x_12306 = v_3271 | ~v_3133;
assign x_12307 = v_3271 | ~v_3134;
assign x_12308 = v_3271 | ~v_3199;
assign x_12309 = v_3271 | ~v_3135;
assign x_12310 = v_3271 | ~v_839;
assign x_12311 = v_3271 | ~v_3200;
assign x_12312 = v_3271 | ~v_1257;
assign x_12313 = v_3271 | ~v_1023;
assign x_12314 = v_3271 | ~v_3136;
assign x_12315 = v_3271 | ~v_3137;
assign x_12316 = v_3271 | ~v_3201;
assign x_12317 = v_3271 | ~v_3138;
assign x_12318 = v_3271 | ~v_840;
assign x_12319 = v_3271 | ~v_3202;
assign x_12320 = v_3271 | ~v_1258;
assign x_12321 = v_3271 | ~v_1024;
assign x_12322 = v_3271 | ~v_184;
assign x_12323 = v_3271 | ~v_170;
assign x_12324 = v_3271 | ~v_149;
assign x_12325 = v_3271 | ~v_1259;
assign x_12326 = v_3271 | ~v_1260;
assign x_12327 = v_3271 | ~v_103;
assign x_12328 = v_3271 | ~v_102;
assign x_12329 = v_3271 | ~v_101;
assign x_12330 = v_3271 | ~v_100;
assign x_12331 = v_3271 | ~v_99;
assign x_12332 = v_3271 | ~v_98;
assign x_12333 = v_3271 | ~v_96;
assign x_12334 = v_3271 | ~v_95;
assign x_12335 = v_3271 | ~v_93;
assign x_12336 = v_3270 | ~v_3110;
assign x_12337 = v_3270 | ~v_3111;
assign x_12338 = v_3270 | ~v_784;
assign x_12339 = v_3270 | ~v_785;
assign x_12340 = v_3270 | ~v_996;
assign x_12341 = v_3270 | ~v_786;
assign x_12342 = v_3270 | ~v_997;
assign x_12343 = v_3270 | ~v_3112;
assign x_12344 = v_3270 | ~v_3113;
assign x_12345 = v_3270 | ~v_787;
assign x_12346 = v_3270 | ~v_788;
assign x_12347 = v_3270 | ~v_998;
assign x_12348 = v_3270 | ~v_789;
assign x_12349 = v_3270 | ~v_999;
assign x_12350 = v_3270 | ~v_3118;
assign x_12351 = v_3270 | ~v_3119;
assign x_12352 = v_3270 | ~v_3194;
assign x_12353 = v_3270 | ~v_3120;
assign x_12354 = v_3270 | ~v_806;
assign x_12355 = v_3270 | ~v_3195;
assign x_12356 = v_3270 | ~v_1252;
assign x_12357 = v_3270 | ~v_1008;
assign x_12358 = v_3270 | ~v_3121;
assign x_12359 = v_3270 | ~v_3122;
assign x_12360 = v_3270 | ~v_1253;
assign x_12361 = v_3270 | ~v_1009;
assign x_12362 = v_3270 | ~v_3123;
assign x_12363 = v_3270 | ~v_807;
assign x_12364 = v_3270 | ~v_3196;
assign x_12365 = v_3270 | ~v_183;
assign x_12366 = v_3270 | ~v_166;
assign x_12367 = v_3270 | ~v_144;
assign x_12368 = v_3270 | ~v_3197;
assign x_12369 = v_3270 | ~v_1254;
assign x_12370 = v_3270 | ~v_1255;
assign x_12371 = v_3270 | ~v_61;
assign x_12372 = v_3270 | ~v_60;
assign x_12373 = v_3270 | ~v_59;
assign x_12374 = v_3270 | ~v_58;
assign x_12375 = v_3270 | ~v_57;
assign x_12376 = v_3270 | ~v_56;
assign x_12377 = v_3270 | ~v_54;
assign x_12378 = v_3270 | ~v_53;
assign x_12379 = v_3270 | ~v_51;
assign x_12380 = v_3269 | ~v_3095;
assign x_12381 = v_3269 | ~v_3096;
assign x_12382 = v_3269 | ~v_751;
assign x_12383 = v_3269 | ~v_752;
assign x_12384 = v_3269 | ~v_981;
assign x_12385 = v_3269 | ~v_753;
assign x_12386 = v_3269 | ~v_982;
assign x_12387 = v_3269 | ~v_3097;
assign x_12388 = v_3269 | ~v_3098;
assign x_12389 = v_3269 | ~v_754;
assign x_12390 = v_3269 | ~v_755;
assign x_12391 = v_3269 | ~v_983;
assign x_12392 = v_3269 | ~v_756;
assign x_12393 = v_3269 | ~v_984;
assign x_12394 = v_3269 | ~v_3103;
assign x_12395 = v_3269 | ~v_3189;
assign x_12396 = v_3269 | ~v_3104;
assign x_12397 = v_3269 | ~v_773;
assign x_12398 = v_3269 | ~v_3190;
assign x_12399 = v_3269 | ~v_3105;
assign x_12400 = v_3269 | ~v_3191;
assign x_12401 = v_3269 | ~v_3106;
assign x_12402 = v_3269 | ~v_774;
assign x_12403 = v_3269 | ~v_3192;
assign x_12404 = v_3269 | ~v_182;
assign x_12405 = v_3269 | ~v_162;
assign x_12406 = v_3269 | ~v_1247;
assign x_12407 = v_3269 | ~v_1248;
assign x_12408 = v_3269 | ~v_136;
assign x_12409 = v_3269 | ~v_3107;
assign x_12410 = v_3269 | ~v_1249;
assign x_12411 = v_3269 | ~v_993;
assign x_12412 = v_3269 | ~v_3108;
assign x_12413 = v_3269 | ~v_1250;
assign x_12414 = v_3269 | ~v_994;
assign x_12415 = v_3269 | ~v_18;
assign x_12416 = v_3269 | ~v_17;
assign x_12417 = v_3269 | ~v_16;
assign x_12418 = v_3269 | ~v_15;
assign x_12419 = v_3269 | ~v_14;
assign x_12420 = v_3269 | ~v_13;
assign x_12421 = v_3269 | ~v_11;
assign x_12422 = v_3269 | ~v_10;
assign x_12423 = v_3269 | ~v_8;
assign x_12424 = ~v_3267 | ~v_3266 | ~v_3265 | v_3268;
assign x_12425 = v_3267 | ~v_873;
assign x_12426 = v_3267 | ~v_874;
assign x_12427 = v_3267 | ~v_875;
assign x_12428 = v_3267 | ~v_876;
assign x_12429 = v_3267 | ~v_3125;
assign x_12430 = v_3267 | ~v_3126;
assign x_12431 = v_3267 | ~v_817;
assign x_12432 = v_3267 | ~v_1011;
assign x_12433 = v_3267 | ~v_1012;
assign x_12434 = v_3267 | ~v_3127;
assign x_12435 = v_3267 | ~v_3128;
assign x_12436 = v_3267 | ~v_820;
assign x_12437 = v_3267 | ~v_1013;
assign x_12438 = v_3267 | ~v_1014;
assign x_12439 = v_3267 | ~v_3251;
assign x_12440 = v_3267 | ~v_3252;
assign x_12441 = v_3267 | ~v_885;
assign x_12442 = v_3267 | ~v_1019;
assign x_12443 = v_3267 | ~v_1020;
assign x_12444 = v_3267 | ~v_3253;
assign x_12445 = v_3267 | ~v_3254;
assign x_12446 = v_3267 | ~v_886;
assign x_12447 = v_3267 | ~v_1021;
assign x_12448 = v_3267 | ~v_1022;
assign x_12449 = v_3267 | ~v_3133;
assign x_12450 = v_3267 | ~v_3199;
assign x_12451 = v_3267 | ~v_3200;
assign x_12452 = v_3267 | ~v_1023;
assign x_12453 = v_3267 | ~v_3136;
assign x_12454 = v_3267 | ~v_3201;
assign x_12455 = v_3267 | ~v_3202;
assign x_12456 = v_3267 | ~v_1024;
assign x_12457 = v_3267 | ~v_184;
assign x_12458 = v_3267 | ~v_181;
assign x_12459 = v_3267 | ~v_171;
assign x_12460 = v_3267 | ~v_169;
assign x_12461 = v_3267 | ~v_149;
assign x_12462 = v_3267 | ~v_147;
assign x_12463 = v_3267 | ~v_103;
assign x_12464 = v_3267 | ~v_102;
assign x_12465 = v_3267 | ~v_101;
assign x_12466 = v_3267 | ~v_99;
assign x_12467 = v_3267 | ~v_96;
assign x_12468 = v_3267 | ~v_94;
assign x_12469 = v_3266 | ~v_858;
assign x_12470 = v_3266 | ~v_859;
assign x_12471 = v_3266 | ~v_860;
assign x_12472 = v_3266 | ~v_861;
assign x_12473 = v_3266 | ~v_3110;
assign x_12474 = v_3266 | ~v_3111;
assign x_12475 = v_3266 | ~v_784;
assign x_12476 = v_3266 | ~v_996;
assign x_12477 = v_3266 | ~v_997;
assign x_12478 = v_3266 | ~v_3112;
assign x_12479 = v_3266 | ~v_3113;
assign x_12480 = v_3266 | ~v_787;
assign x_12481 = v_3266 | ~v_998;
assign x_12482 = v_3266 | ~v_999;
assign x_12483 = v_3266 | ~v_3246;
assign x_12484 = v_3266 | ~v_3247;
assign x_12485 = v_3266 | ~v_870;
assign x_12486 = v_3266 | ~v_1004;
assign x_12487 = v_3266 | ~v_1005;
assign x_12488 = v_3266 | ~v_3248;
assign x_12489 = v_3266 | ~v_3249;
assign x_12490 = v_3266 | ~v_871;
assign x_12491 = v_3266 | ~v_1006;
assign x_12492 = v_3266 | ~v_1007;
assign x_12493 = v_3266 | ~v_3118;
assign x_12494 = v_3266 | ~v_3194;
assign x_12495 = v_3266 | ~v_3195;
assign x_12496 = v_3266 | ~v_1008;
assign x_12497 = v_3266 | ~v_3121;
assign x_12498 = v_3266 | ~v_1009;
assign x_12499 = v_3266 | ~v_3196;
assign x_12500 = v_3266 | ~v_183;
assign x_12501 = v_3266 | ~v_180;
assign x_12502 = v_3266 | ~v_167;
assign x_12503 = v_3266 | ~v_165;
assign x_12504 = v_3266 | ~v_144;
assign x_12505 = v_3266 | ~v_142;
assign x_12506 = v_3266 | ~v_3197;
assign x_12507 = v_3266 | ~v_61;
assign x_12508 = v_3266 | ~v_60;
assign x_12509 = v_3266 | ~v_59;
assign x_12510 = v_3266 | ~v_57;
assign x_12511 = v_3266 | ~v_54;
assign x_12512 = v_3266 | ~v_52;
assign x_12513 = v_3265 | ~v_843;
assign x_12514 = v_3265 | ~v_844;
assign x_12515 = v_3265 | ~v_845;
assign x_12516 = v_3265 | ~v_846;
assign x_12517 = v_3265 | ~v_3095;
assign x_12518 = v_3265 | ~v_3096;
assign x_12519 = v_3265 | ~v_751;
assign x_12520 = v_3265 | ~v_981;
assign x_12521 = v_3265 | ~v_982;
assign x_12522 = v_3265 | ~v_3097;
assign x_12523 = v_3265 | ~v_3098;
assign x_12524 = v_3265 | ~v_754;
assign x_12525 = v_3265 | ~v_983;
assign x_12526 = v_3265 | ~v_984;
assign x_12527 = v_3265 | ~v_3241;
assign x_12528 = v_3265 | ~v_3242;
assign x_12529 = v_3265 | ~v_855;
assign x_12530 = v_3265 | ~v_989;
assign x_12531 = v_3265 | ~v_990;
assign x_12532 = v_3265 | ~v_3243;
assign x_12533 = v_3265 | ~v_3244;
assign x_12534 = v_3265 | ~v_856;
assign x_12535 = v_3265 | ~v_991;
assign x_12536 = v_3265 | ~v_992;
assign x_12537 = v_3265 | ~v_3189;
assign x_12538 = v_3265 | ~v_3190;
assign x_12539 = v_3265 | ~v_3191;
assign x_12540 = v_3265 | ~v_3192;
assign x_12541 = v_3265 | ~v_182;
assign x_12542 = v_3265 | ~v_179;
assign x_12543 = v_3265 | ~v_163;
assign x_12544 = v_3265 | ~v_161;
assign x_12545 = v_3265 | ~v_136;
assign x_12546 = v_3265 | ~v_134;
assign x_12547 = v_3265 | ~v_3107;
assign x_12548 = v_3265 | ~v_993;
assign x_12549 = v_3265 | ~v_3108;
assign x_12550 = v_3265 | ~v_994;
assign x_12551 = v_3265 | ~v_18;
assign x_12552 = v_3265 | ~v_17;
assign x_12553 = v_3265 | ~v_16;
assign x_12554 = v_3265 | ~v_14;
assign x_12555 = v_3265 | ~v_11;
assign x_12556 = v_3265 | ~v_9;
assign x_12557 = ~v_3263 | ~v_3262 | ~v_3261 | v_3264;
assign x_12558 = v_3263 | ~v_813;
assign x_12559 = v_3263 | ~v_814;
assign x_12560 = v_3263 | ~v_815;
assign x_12561 = v_3263 | ~v_816;
assign x_12562 = v_3263 | ~v_873;
assign x_12563 = v_3263 | ~v_874;
assign x_12564 = v_3263 | ~v_875;
assign x_12565 = v_3263 | ~v_876;
assign x_12566 = v_3263 | ~v_3125;
assign x_12567 = v_3263 | ~v_3126;
assign x_12568 = v_3263 | ~v_817;
assign x_12569 = v_3263 | ~v_3127;
assign x_12570 = v_3263 | ~v_3128;
assign x_12571 = v_3263 | ~v_820;
assign x_12572 = v_3263 | ~v_881;
assign x_12573 = v_3263 | ~v_882;
assign x_12574 = v_3263 | ~v_883;
assign x_12575 = v_3263 | ~v_884;
assign x_12576 = v_3263 | ~v_3251;
assign x_12577 = v_3263 | ~v_3252;
assign x_12578 = v_3263 | ~v_885;
assign x_12579 = v_3263 | ~v_3253;
assign x_12580 = v_3263 | ~v_3254;
assign x_12581 = v_3263 | ~v_886;
assign x_12582 = v_3263 | ~v_3183;
assign x_12583 = v_3263 | ~v_3184;
assign x_12584 = v_3263 | ~v_837;
assign x_12585 = v_3263 | ~v_3185;
assign x_12586 = v_3263 | ~v_3186;
assign x_12587 = v_3263 | ~v_838;
assign x_12588 = v_3263 | ~v_3133;
assign x_12589 = v_3263 | ~v_3136;
assign x_12590 = v_3263 | ~v_184;
assign x_12591 = v_3263 | ~v_181;
assign x_12592 = v_3263 | ~v_171;
assign x_12593 = v_3263 | ~v_169;
assign x_12594 = v_3263 | ~v_160;
assign x_12595 = v_3263 | ~v_150;
assign x_12596 = v_3263 | ~v_148;
assign x_12597 = v_3263 | ~v_103;
assign x_12598 = v_3263 | ~v_102;
assign x_12599 = v_3263 | ~v_97;
assign x_12600 = v_3263 | ~v_95;
assign x_12601 = v_3263 | ~v_94;
assign x_12602 = v_3262 | ~v_780;
assign x_12603 = v_3262 | ~v_781;
assign x_12604 = v_3262 | ~v_782;
assign x_12605 = v_3262 | ~v_783;
assign x_12606 = v_3262 | ~v_858;
assign x_12607 = v_3262 | ~v_859;
assign x_12608 = v_3262 | ~v_860;
assign x_12609 = v_3262 | ~v_861;
assign x_12610 = v_3262 | ~v_3110;
assign x_12611 = v_3262 | ~v_3111;
assign x_12612 = v_3262 | ~v_784;
assign x_12613 = v_3262 | ~v_3112;
assign x_12614 = v_3262 | ~v_3113;
assign x_12615 = v_3262 | ~v_787;
assign x_12616 = v_3262 | ~v_866;
assign x_12617 = v_3262 | ~v_867;
assign x_12618 = v_3262 | ~v_868;
assign x_12619 = v_3262 | ~v_869;
assign x_12620 = v_3262 | ~v_3246;
assign x_12621 = v_3262 | ~v_3247;
assign x_12622 = v_3262 | ~v_870;
assign x_12623 = v_3262 | ~v_3248;
assign x_12624 = v_3262 | ~v_3249;
assign x_12625 = v_3262 | ~v_871;
assign x_12626 = v_3262 | ~v_3178;
assign x_12627 = v_3262 | ~v_3179;
assign x_12628 = v_3262 | ~v_804;
assign x_12629 = v_3262 | ~v_3180;
assign x_12630 = v_3262 | ~v_3181;
assign x_12631 = v_3262 | ~v_805;
assign x_12632 = v_3262 | ~v_3118;
assign x_12633 = v_3262 | ~v_3121;
assign x_12634 = v_3262 | ~v_183;
assign x_12635 = v_3262 | ~v_180;
assign x_12636 = v_3262 | ~v_167;
assign x_12637 = v_3262 | ~v_165;
assign x_12638 = v_3262 | ~v_159;
assign x_12639 = v_3262 | ~v_145;
assign x_12640 = v_3262 | ~v_143;
assign x_12641 = v_3262 | ~v_61;
assign x_12642 = v_3262 | ~v_60;
assign x_12643 = v_3262 | ~v_55;
assign x_12644 = v_3262 | ~v_53;
assign x_12645 = v_3262 | ~v_52;
assign x_12646 = v_3261 | ~v_747;
assign x_12647 = v_3261 | ~v_748;
assign x_12648 = v_3261 | ~v_749;
assign x_12649 = v_3261 | ~v_750;
assign x_12650 = v_3261 | ~v_843;
assign x_12651 = v_3261 | ~v_844;
assign x_12652 = v_3261 | ~v_845;
assign x_12653 = v_3261 | ~v_846;
assign x_12654 = v_3261 | ~v_3095;
assign x_12655 = v_3261 | ~v_3096;
assign x_12656 = v_3261 | ~v_751;
assign x_12657 = v_3261 | ~v_3097;
assign x_12658 = v_3261 | ~v_3098;
assign x_12659 = v_3261 | ~v_754;
assign x_12660 = v_3261 | ~v_851;
assign x_12661 = v_3261 | ~v_852;
assign x_12662 = v_3261 | ~v_853;
assign x_12663 = v_3261 | ~v_854;
assign x_12664 = v_3261 | ~v_3241;
assign x_12665 = v_3261 | ~v_3242;
assign x_12666 = v_3261 | ~v_855;
assign x_12667 = v_3261 | ~v_3243;
assign x_12668 = v_3261 | ~v_3244;
assign x_12669 = v_3261 | ~v_856;
assign x_12670 = v_3261 | ~v_3173;
assign x_12671 = v_3261 | ~v_3174;
assign x_12672 = v_3261 | ~v_771;
assign x_12673 = v_3261 | ~v_3175;
assign x_12674 = v_3261 | ~v_3176;
assign x_12675 = v_3261 | ~v_772;
assign x_12676 = v_3261 | ~v_182;
assign x_12677 = v_3261 | ~v_179;
assign x_12678 = v_3261 | ~v_163;
assign x_12679 = v_3261 | ~v_161;
assign x_12680 = v_3261 | ~v_155;
assign x_12681 = v_3261 | ~v_137;
assign x_12682 = v_3261 | ~v_135;
assign x_12683 = v_3261 | ~v_3107;
assign x_12684 = v_3261 | ~v_3108;
assign x_12685 = v_3261 | ~v_18;
assign x_12686 = v_3261 | ~v_17;
assign x_12687 = v_3261 | ~v_12;
assign x_12688 = v_3261 | ~v_10;
assign x_12689 = v_3261 | ~v_9;
assign x_12690 = ~v_3259 | ~v_3258 | ~v_3257 | v_3260;
assign x_12691 = v_3259 | ~v_919;
assign x_12692 = v_3259 | ~v_920;
assign x_12693 = v_3259 | ~v_873;
assign x_12694 = v_3259 | ~v_874;
assign x_12695 = v_3259 | ~v_875;
assign x_12696 = v_3259 | ~v_876;
assign x_12697 = v_3259 | ~v_3125;
assign x_12698 = v_3259 | ~v_3126;
assign x_12699 = v_3259 | ~v_817;
assign x_12700 = v_3259 | ~v_3127;
assign x_12701 = v_3259 | ~v_3128;
assign x_12702 = v_3259 | ~v_820;
assign x_12703 = v_3259 | ~v_925;
assign x_12704 = v_3259 | ~v_926;
assign x_12705 = v_3259 | ~v_3251;
assign x_12706 = v_3259 | ~v_3252;
assign x_12707 = v_3259 | ~v_885;
assign x_12708 = v_3259 | ~v_3253;
assign x_12709 = v_3259 | ~v_3254;
assign x_12710 = v_3259 | ~v_886;
assign x_12711 = v_3259 | ~v_3167;
assign x_12712 = v_3259 | ~v_3168;
assign x_12713 = v_3259 | ~v_927;
assign x_12714 = v_3259 | ~v_3169;
assign x_12715 = v_3259 | ~v_3170;
assign x_12716 = v_3259 | ~v_928;
assign x_12717 = v_3259 | ~v_3133;
assign x_12718 = v_3259 | ~v_3136;
assign x_12719 = v_3259 | ~v_929;
assign x_12720 = v_3259 | ~v_930;
assign x_12721 = v_3259 | ~v_931;
assign x_12722 = v_3259 | ~v_932;
assign x_12723 = v_3259 | ~v_184;
assign x_12724 = v_3259 | ~v_181;
assign x_12725 = v_3259 | ~v_171;
assign x_12726 = v_3259 | ~v_169;
assign x_12727 = v_3259 | ~v_150;
assign x_12728 = v_3259 | ~v_149;
assign x_12729 = v_3259 | ~v_148;
assign x_12730 = v_3259 | ~v_147;
assign x_12731 = v_3259 | ~v_103;
assign x_12732 = v_3259 | ~v_102;
assign x_12733 = v_3259 | ~v_101;
assign x_12734 = v_3259 | ~v_94;
assign x_12735 = v_3258 | ~v_904;
assign x_12736 = v_3258 | ~v_905;
assign x_12737 = v_3258 | ~v_858;
assign x_12738 = v_3258 | ~v_859;
assign x_12739 = v_3258 | ~v_860;
assign x_12740 = v_3258 | ~v_861;
assign x_12741 = v_3258 | ~v_3110;
assign x_12742 = v_3258 | ~v_3111;
assign x_12743 = v_3258 | ~v_784;
assign x_12744 = v_3258 | ~v_3112;
assign x_12745 = v_3258 | ~v_3113;
assign x_12746 = v_3258 | ~v_787;
assign x_12747 = v_3258 | ~v_910;
assign x_12748 = v_3258 | ~v_911;
assign x_12749 = v_3258 | ~v_3246;
assign x_12750 = v_3258 | ~v_3247;
assign x_12751 = v_3258 | ~v_870;
assign x_12752 = v_3258 | ~v_3248;
assign x_12753 = v_3258 | ~v_3249;
assign x_12754 = v_3258 | ~v_871;
assign x_12755 = v_3258 | ~v_3162;
assign x_12756 = v_3258 | ~v_3163;
assign x_12757 = v_3258 | ~v_912;
assign x_12758 = v_3258 | ~v_3164;
assign x_12759 = v_3258 | ~v_3165;
assign x_12760 = v_3258 | ~v_913;
assign x_12761 = v_3258 | ~v_3118;
assign x_12762 = v_3258 | ~v_3121;
assign x_12763 = v_3258 | ~v_914;
assign x_12764 = v_3258 | ~v_915;
assign x_12765 = v_3258 | ~v_916;
assign x_12766 = v_3258 | ~v_917;
assign x_12767 = v_3258 | ~v_183;
assign x_12768 = v_3258 | ~v_180;
assign x_12769 = v_3258 | ~v_167;
assign x_12770 = v_3258 | ~v_165;
assign x_12771 = v_3258 | ~v_145;
assign x_12772 = v_3258 | ~v_144;
assign x_12773 = v_3258 | ~v_143;
assign x_12774 = v_3258 | ~v_142;
assign x_12775 = v_3258 | ~v_61;
assign x_12776 = v_3258 | ~v_60;
assign x_12777 = v_3258 | ~v_59;
assign x_12778 = v_3258 | ~v_52;
assign x_12779 = v_3257 | ~v_889;
assign x_12780 = v_3257 | ~v_890;
assign x_12781 = v_3257 | ~v_843;
assign x_12782 = v_3257 | ~v_844;
assign x_12783 = v_3257 | ~v_845;
assign x_12784 = v_3257 | ~v_846;
assign x_12785 = v_3257 | ~v_3095;
assign x_12786 = v_3257 | ~v_3096;
assign x_12787 = v_3257 | ~v_751;
assign x_12788 = v_3257 | ~v_3097;
assign x_12789 = v_3257 | ~v_3098;
assign x_12790 = v_3257 | ~v_754;
assign x_12791 = v_3257 | ~v_895;
assign x_12792 = v_3257 | ~v_896;
assign x_12793 = v_3257 | ~v_3241;
assign x_12794 = v_3257 | ~v_3242;
assign x_12795 = v_3257 | ~v_855;
assign x_12796 = v_3257 | ~v_3243;
assign x_12797 = v_3257 | ~v_3244;
assign x_12798 = v_3257 | ~v_856;
assign x_12799 = v_3257 | ~v_3157;
assign x_12800 = v_3257 | ~v_3158;
assign x_12801 = v_3257 | ~v_897;
assign x_12802 = v_3257 | ~v_3159;
assign x_12803 = v_3257 | ~v_3160;
assign x_12804 = v_3257 | ~v_898;
assign x_12805 = v_3257 | ~v_899;
assign x_12806 = v_3257 | ~v_900;
assign x_12807 = v_3257 | ~v_901;
assign x_12808 = v_3257 | ~v_902;
assign x_12809 = v_3257 | ~v_182;
assign x_12810 = v_3257 | ~v_179;
assign x_12811 = v_3257 | ~v_163;
assign x_12812 = v_3257 | ~v_161;
assign x_12813 = v_3257 | ~v_137;
assign x_12814 = v_3257 | ~v_136;
assign x_12815 = v_3257 | ~v_135;
assign x_12816 = v_3257 | ~v_134;
assign x_12817 = v_3257 | ~v_3107;
assign x_12818 = v_3257 | ~v_3108;
assign x_12819 = v_3257 | ~v_18;
assign x_12820 = v_3257 | ~v_17;
assign x_12821 = v_3257 | ~v_16;
assign x_12822 = v_3257 | ~v_9;
assign x_12823 = ~v_3255 | ~v_3250 | ~v_3245 | v_3256;
assign x_12824 = v_3255 | ~v_965;
assign x_12825 = v_3255 | ~v_966;
assign x_12826 = v_3255 | ~v_967;
assign x_12827 = v_3255 | ~v_968;
assign x_12828 = v_3255 | ~v_873;
assign x_12829 = v_3255 | ~v_874;
assign x_12830 = v_3255 | ~v_875;
assign x_12831 = v_3255 | ~v_876;
assign x_12832 = v_3255 | ~v_3125;
assign x_12833 = v_3255 | ~v_3126;
assign x_12834 = v_3255 | ~v_817;
assign x_12835 = v_3255 | ~v_3127;
assign x_12836 = v_3255 | ~v_3128;
assign x_12837 = v_3255 | ~v_820;
assign x_12838 = v_3255 | ~v_973;
assign x_12839 = v_3255 | ~v_974;
assign x_12840 = v_3255 | ~v_3251;
assign x_12841 = v_3255 | ~v_3252;
assign x_12842 = v_3255 | ~v_885;
assign x_12843 = v_3255 | ~v_3253;
assign x_12844 = v_3255 | ~v_3254;
assign x_12845 = v_3255 | ~v_886;
assign x_12846 = v_3255 | ~v_3129;
assign x_12847 = v_3255 | ~v_3130;
assign x_12848 = v_3255 | ~v_975;
assign x_12849 = v_3255 | ~v_3131;
assign x_12850 = v_3255 | ~v_3132;
assign x_12851 = v_3255 | ~v_976;
assign x_12852 = v_3255 | ~v_3133;
assign x_12853 = v_3255 | ~v_3136;
assign x_12854 = v_3255 | ~v_977;
assign x_12855 = v_3255 | ~v_978;
assign x_12856 = v_3255 | ~v_184;
assign x_12857 = v_3255 | ~v_181;
assign x_12858 = v_3255 | ~v_172;
assign x_12859 = v_3255 | ~v_171;
assign x_12860 = v_3255 | ~v_169;
assign x_12861 = v_3255 | ~v_150;
assign x_12862 = v_3255 | ~v_149;
assign x_12863 = v_3255 | ~v_148;
assign x_12864 = v_3255 | ~v_147;
assign x_12865 = v_3255 | ~v_102;
assign x_12866 = v_3255 | ~v_101;
assign x_12867 = v_3255 | ~v_94;
assign x_12868 = ~v_127 | ~v_157 | v_3254;
assign x_12869 = ~v_121 | ~v_156 | v_3253;
assign x_12870 = ~v_112 | v_157 | v_3252;
assign x_12871 = ~v_106 | v_156 | v_3251;
assign x_12872 = v_3250 | ~v_950;
assign x_12873 = v_3250 | ~v_951;
assign x_12874 = v_3250 | ~v_952;
assign x_12875 = v_3250 | ~v_953;
assign x_12876 = v_3250 | ~v_858;
assign x_12877 = v_3250 | ~v_859;
assign x_12878 = v_3250 | ~v_860;
assign x_12879 = v_3250 | ~v_861;
assign x_12880 = v_3250 | ~v_3110;
assign x_12881 = v_3250 | ~v_3111;
assign x_12882 = v_3250 | ~v_784;
assign x_12883 = v_3250 | ~v_3112;
assign x_12884 = v_3250 | ~v_3113;
assign x_12885 = v_3250 | ~v_787;
assign x_12886 = v_3250 | ~v_958;
assign x_12887 = v_3250 | ~v_959;
assign x_12888 = v_3250 | ~v_3246;
assign x_12889 = v_3250 | ~v_3247;
assign x_12890 = v_3250 | ~v_870;
assign x_12891 = v_3250 | ~v_3248;
assign x_12892 = v_3250 | ~v_3249;
assign x_12893 = v_3250 | ~v_871;
assign x_12894 = v_3250 | ~v_3114;
assign x_12895 = v_3250 | ~v_3115;
assign x_12896 = v_3250 | ~v_960;
assign x_12897 = v_3250 | ~v_3116;
assign x_12898 = v_3250 | ~v_3117;
assign x_12899 = v_3250 | ~v_961;
assign x_12900 = v_3250 | ~v_3118;
assign x_12901 = v_3250 | ~v_3121;
assign x_12902 = v_3250 | ~v_962;
assign x_12903 = v_3250 | ~v_963;
assign x_12904 = v_3250 | ~v_183;
assign x_12905 = v_3250 | ~v_180;
assign x_12906 = v_3250 | ~v_168;
assign x_12907 = v_3250 | ~v_167;
assign x_12908 = v_3250 | ~v_165;
assign x_12909 = v_3250 | ~v_145;
assign x_12910 = v_3250 | ~v_144;
assign x_12911 = v_3250 | ~v_143;
assign x_12912 = v_3250 | ~v_142;
assign x_12913 = v_3250 | ~v_60;
assign x_12914 = v_3250 | ~v_59;
assign x_12915 = v_3250 | ~v_52;
assign x_12916 = ~v_85 | ~v_157 | v_3249;
assign x_12917 = ~v_79 | ~v_156 | v_3248;
assign x_12918 = ~v_70 | v_157 | v_3247;
assign x_12919 = ~v_64 | v_156 | v_3246;
assign x_12920 = v_3245 | ~v_935;
assign x_12921 = v_3245 | ~v_936;
assign x_12922 = v_3245 | ~v_937;
assign x_12923 = v_3245 | ~v_938;
assign x_12924 = v_3245 | ~v_843;
assign x_12925 = v_3245 | ~v_844;
assign x_12926 = v_3245 | ~v_845;
assign x_12927 = v_3245 | ~v_846;
assign x_12928 = v_3245 | ~v_3095;
assign x_12929 = v_3245 | ~v_3096;
assign x_12930 = v_3245 | ~v_751;
assign x_12931 = v_3245 | ~v_3097;
assign x_12932 = v_3245 | ~v_3098;
assign x_12933 = v_3245 | ~v_754;
assign x_12934 = v_3245 | ~v_943;
assign x_12935 = v_3245 | ~v_944;
assign x_12936 = v_3245 | ~v_3241;
assign x_12937 = v_3245 | ~v_3242;
assign x_12938 = v_3245 | ~v_855;
assign x_12939 = v_3245 | ~v_3243;
assign x_12940 = v_3245 | ~v_3244;
assign x_12941 = v_3245 | ~v_856;
assign x_12942 = v_3245 | ~v_3099;
assign x_12943 = v_3245 | ~v_3100;
assign x_12944 = v_3245 | ~v_945;
assign x_12945 = v_3245 | ~v_3101;
assign x_12946 = v_3245 | ~v_3102;
assign x_12947 = v_3245 | ~v_946;
assign x_12948 = v_3245 | ~v_947;
assign x_12949 = v_3245 | ~v_948;
assign x_12950 = v_3245 | ~v_182;
assign x_12951 = v_3245 | ~v_179;
assign x_12952 = v_3245 | ~v_164;
assign x_12953 = v_3245 | ~v_163;
assign x_12954 = v_3245 | ~v_161;
assign x_12955 = v_3245 | ~v_137;
assign x_12956 = v_3245 | ~v_136;
assign x_12957 = v_3245 | ~v_135;
assign x_12958 = v_3245 | ~v_134;
assign x_12959 = v_3245 | ~v_3107;
assign x_12960 = v_3245 | ~v_3108;
assign x_12961 = v_3245 | ~v_17;
assign x_12962 = v_3245 | ~v_16;
assign x_12963 = v_3245 | ~v_9;
assign x_12964 = ~v_43 | ~v_157 | v_3244;
assign x_12965 = ~v_37 | ~v_156 | v_3243;
assign x_12966 = ~v_28 | v_157 | v_3242;
assign x_12967 = ~v_22 | v_156 | v_3241;
assign x_12968 = ~v_3239 | ~v_3238 | ~v_3237 | v_3240;
assign x_12969 = v_3239 | ~v_813;
assign x_12970 = v_3239 | ~v_814;
assign x_12971 = v_3239 | ~v_815;
assign x_12972 = v_3239 | ~v_816;
assign x_12973 = v_3239 | ~v_3125;
assign x_12974 = v_3239 | ~v_3126;
assign x_12975 = v_3239 | ~v_817;
assign x_12976 = v_3239 | ~v_818;
assign x_12977 = v_3239 | ~v_819;
assign x_12978 = v_3239 | ~v_3127;
assign x_12979 = v_3239 | ~v_3128;
assign x_12980 = v_3239 | ~v_820;
assign x_12981 = v_3239 | ~v_821;
assign x_12982 = v_3239 | ~v_822;
assign x_12983 = v_3239 | ~v_833;
assign x_12984 = v_3239 | ~v_834;
assign x_12985 = v_3239 | ~v_835;
assign x_12986 = v_3239 | ~v_836;
assign x_12987 = v_3239 | ~v_3183;
assign x_12988 = v_3239 | ~v_3184;
assign x_12989 = v_3239 | ~v_837;
assign x_12990 = v_3239 | ~v_3185;
assign x_12991 = v_3239 | ~v_3186;
assign x_12992 = v_3239 | ~v_838;
assign x_12993 = v_3239 | ~v_3133;
assign x_12994 = v_3239 | ~v_3134;
assign x_12995 = v_3239 | ~v_3135;
assign x_12996 = v_3239 | ~v_839;
assign x_12997 = v_3239 | ~v_3136;
assign x_12998 = v_3239 | ~v_3137;
assign x_12999 = v_3239 | ~v_3138;
assign x_13000 = v_3239 | ~v_840;
assign x_13001 = v_3239 | ~v_184;
assign x_13002 = v_3239 | ~v_170;
assign x_13003 = v_3239 | ~v_160;
assign x_13004 = v_3239 | ~v_150;
assign x_13005 = v_3239 | ~v_148;
assign x_13006 = v_3239 | ~v_147;
assign x_13007 = v_3239 | ~v_103;
assign x_13008 = v_3239 | ~v_102;
assign x_13009 = v_3239 | ~v_100;
assign x_13010 = v_3239 | ~v_98;
assign x_13011 = v_3239 | ~v_97;
assign x_13012 = v_3239 | ~v_93;
assign x_13013 = v_3238 | ~v_780;
assign x_13014 = v_3238 | ~v_781;
assign x_13015 = v_3238 | ~v_782;
assign x_13016 = v_3238 | ~v_783;
assign x_13017 = v_3238 | ~v_3110;
assign x_13018 = v_3238 | ~v_3111;
assign x_13019 = v_3238 | ~v_784;
assign x_13020 = v_3238 | ~v_785;
assign x_13021 = v_3238 | ~v_786;
assign x_13022 = v_3238 | ~v_3112;
assign x_13023 = v_3238 | ~v_3113;
assign x_13024 = v_3238 | ~v_787;
assign x_13025 = v_3238 | ~v_788;
assign x_13026 = v_3238 | ~v_789;
assign x_13027 = v_3238 | ~v_800;
assign x_13028 = v_3238 | ~v_801;
assign x_13029 = v_3238 | ~v_802;
assign x_13030 = v_3238 | ~v_803;
assign x_13031 = v_3238 | ~v_3178;
assign x_13032 = v_3238 | ~v_3179;
assign x_13033 = v_3238 | ~v_804;
assign x_13034 = v_3238 | ~v_3180;
assign x_13035 = v_3238 | ~v_3181;
assign x_13036 = v_3238 | ~v_805;
assign x_13037 = v_3238 | ~v_3118;
assign x_13038 = v_3238 | ~v_3119;
assign x_13039 = v_3238 | ~v_3120;
assign x_13040 = v_3238 | ~v_806;
assign x_13041 = v_3238 | ~v_3121;
assign x_13042 = v_3238 | ~v_3122;
assign x_13043 = v_3238 | ~v_3123;
assign x_13044 = v_3238 | ~v_807;
assign x_13045 = v_3238 | ~v_183;
assign x_13046 = v_3238 | ~v_166;
assign x_13047 = v_3238 | ~v_159;
assign x_13048 = v_3238 | ~v_145;
assign x_13049 = v_3238 | ~v_143;
assign x_13050 = v_3238 | ~v_142;
assign x_13051 = v_3238 | ~v_61;
assign x_13052 = v_3238 | ~v_60;
assign x_13053 = v_3238 | ~v_58;
assign x_13054 = v_3238 | ~v_56;
assign x_13055 = v_3238 | ~v_55;
assign x_13056 = v_3238 | ~v_51;
assign x_13057 = v_3237 | ~v_747;
assign x_13058 = v_3237 | ~v_748;
assign x_13059 = v_3237 | ~v_749;
assign x_13060 = v_3237 | ~v_750;
assign x_13061 = v_3237 | ~v_3095;
assign x_13062 = v_3237 | ~v_3096;
assign x_13063 = v_3237 | ~v_751;
assign x_13064 = v_3237 | ~v_752;
assign x_13065 = v_3237 | ~v_753;
assign x_13066 = v_3237 | ~v_3097;
assign x_13067 = v_3237 | ~v_3098;
assign x_13068 = v_3237 | ~v_754;
assign x_13069 = v_3237 | ~v_755;
assign x_13070 = v_3237 | ~v_756;
assign x_13071 = v_3237 | ~v_767;
assign x_13072 = v_3237 | ~v_768;
assign x_13073 = v_3237 | ~v_769;
assign x_13074 = v_3237 | ~v_770;
assign x_13075 = v_3237 | ~v_3173;
assign x_13076 = v_3237 | ~v_3174;
assign x_13077 = v_3237 | ~v_771;
assign x_13078 = v_3237 | ~v_3175;
assign x_13079 = v_3237 | ~v_3176;
assign x_13080 = v_3237 | ~v_772;
assign x_13081 = v_3237 | ~v_3103;
assign x_13082 = v_3237 | ~v_3104;
assign x_13083 = v_3237 | ~v_773;
assign x_13084 = v_3237 | ~v_3105;
assign x_13085 = v_3237 | ~v_3106;
assign x_13086 = v_3237 | ~v_774;
assign x_13087 = v_3237 | ~v_182;
assign x_13088 = v_3237 | ~v_162;
assign x_13089 = v_3237 | ~v_155;
assign x_13090 = v_3237 | ~v_137;
assign x_13091 = v_3237 | ~v_135;
assign x_13092 = v_3237 | ~v_134;
assign x_13093 = v_3237 | ~v_3107;
assign x_13094 = v_3237 | ~v_3108;
assign x_13095 = v_3237 | ~v_18;
assign x_13096 = v_3237 | ~v_17;
assign x_13097 = v_3237 | ~v_15;
assign x_13098 = v_3237 | ~v_13;
assign x_13099 = v_3237 | ~v_12;
assign x_13100 = v_3237 | ~v_8;
assign x_13101 = ~v_3235 | ~v_3234 | ~v_3233 | v_3236;
assign x_13102 = v_3235 | ~v_1073;
assign x_13103 = v_3235 | ~v_1074;
assign x_13104 = v_3235 | ~v_1075;
assign x_13105 = v_3235 | ~v_1076;
assign x_13106 = v_3235 | ~v_3125;
assign x_13107 = v_3235 | ~v_3126;
assign x_13108 = v_3235 | ~v_817;
assign x_13109 = v_3235 | ~v_1011;
assign x_13110 = v_3235 | ~v_1012;
assign x_13111 = v_3235 | ~v_3127;
assign x_13112 = v_3235 | ~v_3128;
assign x_13113 = v_3235 | ~v_820;
assign x_13114 = v_3235 | ~v_1013;
assign x_13115 = v_3235 | ~v_1014;
assign x_13116 = v_3235 | ~v_3219;
assign x_13117 = v_3235 | ~v_3220;
assign x_13118 = v_3235 | ~v_1085;
assign x_13119 = v_3235 | ~v_1131;
assign x_13120 = v_3235 | ~v_1132;
assign x_13121 = v_3235 | ~v_3221;
assign x_13122 = v_3235 | ~v_3222;
assign x_13123 = v_3235 | ~v_1086;
assign x_13124 = v_3235 | ~v_1133;
assign x_13125 = v_3235 | ~v_1134;
assign x_13126 = v_3235 | ~v_3133;
assign x_13127 = v_3235 | ~v_3199;
assign x_13128 = v_3235 | ~v_3200;
assign x_13129 = v_3235 | ~v_1023;
assign x_13130 = v_3235 | ~v_3136;
assign x_13131 = v_3235 | ~v_3201;
assign x_13132 = v_3235 | ~v_3202;
assign x_13133 = v_3235 | ~v_1024;
assign x_13134 = v_3235 | ~v_184;
assign x_13135 = v_3235 | ~v_172;
assign x_13136 = v_3235 | ~v_171;
assign x_13137 = v_3235 | ~v_170;
assign x_13138 = v_3235 | ~v_169;
assign x_13139 = v_3235 | ~v_149;
assign x_13140 = v_3235 | ~v_147;
assign x_13141 = v_3235 | ~v_102;
assign x_13142 = v_3235 | ~v_101;
assign x_13143 = v_3235 | ~v_100;
assign x_13144 = v_3235 | ~v_99;
assign x_13145 = v_3235 | ~v_96;
assign x_13146 = v_3234 | ~v_1058;
assign x_13147 = v_3234 | ~v_1059;
assign x_13148 = v_3234 | ~v_1060;
assign x_13149 = v_3234 | ~v_1061;
assign x_13150 = v_3234 | ~v_3110;
assign x_13151 = v_3234 | ~v_3111;
assign x_13152 = v_3234 | ~v_784;
assign x_13153 = v_3234 | ~v_996;
assign x_13154 = v_3234 | ~v_997;
assign x_13155 = v_3234 | ~v_3112;
assign x_13156 = v_3234 | ~v_3113;
assign x_13157 = v_3234 | ~v_787;
assign x_13158 = v_3234 | ~v_998;
assign x_13159 = v_3234 | ~v_999;
assign x_13160 = v_3234 | ~v_3214;
assign x_13161 = v_3234 | ~v_3215;
assign x_13162 = v_3234 | ~v_1070;
assign x_13163 = v_3234 | ~v_1126;
assign x_13164 = v_3234 | ~v_1127;
assign x_13165 = v_3234 | ~v_3216;
assign x_13166 = v_3234 | ~v_3217;
assign x_13167 = v_3234 | ~v_1071;
assign x_13168 = v_3234 | ~v_1128;
assign x_13169 = v_3234 | ~v_1129;
assign x_13170 = v_3234 | ~v_3118;
assign x_13171 = v_3234 | ~v_3194;
assign x_13172 = v_3234 | ~v_3195;
assign x_13173 = v_3234 | ~v_1008;
assign x_13174 = v_3234 | ~v_3121;
assign x_13175 = v_3234 | ~v_1009;
assign x_13176 = v_3234 | ~v_3196;
assign x_13177 = v_3234 | ~v_183;
assign x_13178 = v_3234 | ~v_168;
assign x_13179 = v_3234 | ~v_167;
assign x_13180 = v_3234 | ~v_166;
assign x_13181 = v_3234 | ~v_165;
assign x_13182 = v_3234 | ~v_144;
assign x_13183 = v_3234 | ~v_142;
assign x_13184 = v_3234 | ~v_3197;
assign x_13185 = v_3234 | ~v_60;
assign x_13186 = v_3234 | ~v_59;
assign x_13187 = v_3234 | ~v_58;
assign x_13188 = v_3234 | ~v_57;
assign x_13189 = v_3234 | ~v_54;
assign x_13190 = v_3233 | ~v_1043;
assign x_13191 = v_3233 | ~v_1044;
assign x_13192 = v_3233 | ~v_1045;
assign x_13193 = v_3233 | ~v_1046;
assign x_13194 = v_3233 | ~v_3095;
assign x_13195 = v_3233 | ~v_3096;
assign x_13196 = v_3233 | ~v_751;
assign x_13197 = v_3233 | ~v_981;
assign x_13198 = v_3233 | ~v_982;
assign x_13199 = v_3233 | ~v_3097;
assign x_13200 = v_3233 | ~v_3098;
assign x_13201 = v_3233 | ~v_754;
assign x_13202 = v_3233 | ~v_983;
assign x_13203 = v_3233 | ~v_984;
assign x_13204 = v_3233 | ~v_3209;
assign x_13205 = v_3233 | ~v_3210;
assign x_13206 = v_3233 | ~v_1055;
assign x_13207 = v_3233 | ~v_1121;
assign x_13208 = v_3233 | ~v_1122;
assign x_13209 = v_3233 | ~v_3211;
assign x_13210 = v_3233 | ~v_3212;
assign x_13211 = v_3233 | ~v_1056;
assign x_13212 = v_3233 | ~v_1123;
assign x_13213 = v_3233 | ~v_1124;
assign x_13214 = v_3233 | ~v_3189;
assign x_13215 = v_3233 | ~v_3190;
assign x_13216 = v_3233 | ~v_3191;
assign x_13217 = v_3233 | ~v_3192;
assign x_13218 = v_3233 | ~v_182;
assign x_13219 = v_3233 | ~v_164;
assign x_13220 = v_3233 | ~v_163;
assign x_13221 = v_3233 | ~v_162;
assign x_13222 = v_3233 | ~v_161;
assign x_13223 = v_3233 | ~v_136;
assign x_13224 = v_3233 | ~v_134;
assign x_13225 = v_3233 | ~v_3107;
assign x_13226 = v_3233 | ~v_993;
assign x_13227 = v_3233 | ~v_3108;
assign x_13228 = v_3233 | ~v_994;
assign x_13229 = v_3233 | ~v_17;
assign x_13230 = v_3233 | ~v_16;
assign x_13231 = v_3233 | ~v_15;
assign x_13232 = v_3233 | ~v_14;
assign x_13233 = v_3233 | ~v_11;
assign x_13234 = ~v_3231 | ~v_3230 | ~v_3229 | v_3232;
assign x_13235 = v_3231 | ~v_1073;
assign x_13236 = v_3231 | ~v_1074;
assign x_13237 = v_3231 | ~v_1075;
assign x_13238 = v_3231 | ~v_1076;
assign x_13239 = v_3231 | ~v_813;
assign x_13240 = v_3231 | ~v_814;
assign x_13241 = v_3231 | ~v_815;
assign x_13242 = v_3231 | ~v_816;
assign x_13243 = v_3231 | ~v_3125;
assign x_13244 = v_3231 | ~v_3126;
assign x_13245 = v_3231 | ~v_817;
assign x_13246 = v_3231 | ~v_3127;
assign x_13247 = v_3231 | ~v_3128;
assign x_13248 = v_3231 | ~v_820;
assign x_13249 = v_3231 | ~v_3183;
assign x_13250 = v_3231 | ~v_3184;
assign x_13251 = v_3231 | ~v_837;
assign x_13252 = v_3231 | ~v_3185;
assign x_13253 = v_3231 | ~v_3186;
assign x_13254 = v_3231 | ~v_838;
assign x_13255 = v_3231 | ~v_1081;
assign x_13256 = v_3231 | ~v_1082;
assign x_13257 = v_3231 | ~v_1083;
assign x_13258 = v_3231 | ~v_1084;
assign x_13259 = v_3231 | ~v_3219;
assign x_13260 = v_3231 | ~v_3220;
assign x_13261 = v_3231 | ~v_1085;
assign x_13262 = v_3231 | ~v_3221;
assign x_13263 = v_3231 | ~v_3222;
assign x_13264 = v_3231 | ~v_1086;
assign x_13265 = v_3231 | ~v_3133;
assign x_13266 = v_3231 | ~v_3136;
assign x_13267 = v_3231 | ~v_184;
assign x_13268 = v_3231 | ~v_171;
assign x_13269 = v_3231 | ~v_170;
assign x_13270 = v_3231 | ~v_169;
assign x_13271 = v_3231 | ~v_160;
assign x_13272 = v_3231 | ~v_150;
assign x_13273 = v_3231 | ~v_148;
assign x_13274 = v_3231 | ~v_147;
assign x_13275 = v_3231 | ~v_103;
assign x_13276 = v_3231 | ~v_102;
assign x_13277 = v_3231 | ~v_100;
assign x_13278 = v_3231 | ~v_97;
assign x_13279 = v_3230 | ~v_1058;
assign x_13280 = v_3230 | ~v_1059;
assign x_13281 = v_3230 | ~v_1060;
assign x_13282 = v_3230 | ~v_1061;
assign x_13283 = v_3230 | ~v_780;
assign x_13284 = v_3230 | ~v_781;
assign x_13285 = v_3230 | ~v_782;
assign x_13286 = v_3230 | ~v_783;
assign x_13287 = v_3230 | ~v_3110;
assign x_13288 = v_3230 | ~v_3111;
assign x_13289 = v_3230 | ~v_784;
assign x_13290 = v_3230 | ~v_3112;
assign x_13291 = v_3230 | ~v_3113;
assign x_13292 = v_3230 | ~v_787;
assign x_13293 = v_3230 | ~v_3178;
assign x_13294 = v_3230 | ~v_3179;
assign x_13295 = v_3230 | ~v_804;
assign x_13296 = v_3230 | ~v_3180;
assign x_13297 = v_3230 | ~v_3181;
assign x_13298 = v_3230 | ~v_805;
assign x_13299 = v_3230 | ~v_1066;
assign x_13300 = v_3230 | ~v_1067;
assign x_13301 = v_3230 | ~v_1068;
assign x_13302 = v_3230 | ~v_1069;
assign x_13303 = v_3230 | ~v_3214;
assign x_13304 = v_3230 | ~v_3215;
assign x_13305 = v_3230 | ~v_1070;
assign x_13306 = v_3230 | ~v_3216;
assign x_13307 = v_3230 | ~v_3217;
assign x_13308 = v_3230 | ~v_1071;
assign x_13309 = v_3230 | ~v_3118;
assign x_13310 = v_3230 | ~v_3121;
assign x_13311 = v_3230 | ~v_183;
assign x_13312 = v_3230 | ~v_167;
assign x_13313 = v_3230 | ~v_166;
assign x_13314 = v_3230 | ~v_165;
assign x_13315 = v_3230 | ~v_159;
assign x_13316 = v_3230 | ~v_145;
assign x_13317 = v_3230 | ~v_143;
assign x_13318 = v_3230 | ~v_142;
assign x_13319 = v_3230 | ~v_61;
assign x_13320 = v_3230 | ~v_60;
assign x_13321 = v_3230 | ~v_58;
assign x_13322 = v_3230 | ~v_55;
assign x_13323 = v_3229 | ~v_1043;
assign x_13324 = v_3229 | ~v_1044;
assign x_13325 = v_3229 | ~v_1045;
assign x_13326 = v_3229 | ~v_1046;
assign x_13327 = v_3229 | ~v_747;
assign x_13328 = v_3229 | ~v_748;
assign x_13329 = v_3229 | ~v_749;
assign x_13330 = v_3229 | ~v_750;
assign x_13331 = v_3229 | ~v_3095;
assign x_13332 = v_3229 | ~v_3096;
assign x_13333 = v_3229 | ~v_751;
assign x_13334 = v_3229 | ~v_3097;
assign x_13335 = v_3229 | ~v_3098;
assign x_13336 = v_3229 | ~v_754;
assign x_13337 = v_3229 | ~v_3173;
assign x_13338 = v_3229 | ~v_3174;
assign x_13339 = v_3229 | ~v_771;
assign x_13340 = v_3229 | ~v_3175;
assign x_13341 = v_3229 | ~v_3176;
assign x_13342 = v_3229 | ~v_772;
assign x_13343 = v_3229 | ~v_1051;
assign x_13344 = v_3229 | ~v_1052;
assign x_13345 = v_3229 | ~v_1053;
assign x_13346 = v_3229 | ~v_1054;
assign x_13347 = v_3229 | ~v_3209;
assign x_13348 = v_3229 | ~v_3210;
assign x_13349 = v_3229 | ~v_1055;
assign x_13350 = v_3229 | ~v_3211;
assign x_13351 = v_3229 | ~v_3212;
assign x_13352 = v_3229 | ~v_1056;
assign x_13353 = v_3229 | ~v_182;
assign x_13354 = v_3229 | ~v_163;
assign x_13355 = v_3229 | ~v_162;
assign x_13356 = v_3229 | ~v_161;
assign x_13357 = v_3229 | ~v_155;
assign x_13358 = v_3229 | ~v_137;
assign x_13359 = v_3229 | ~v_135;
assign x_13360 = v_3229 | ~v_134;
assign x_13361 = v_3229 | ~v_3107;
assign x_13362 = v_3229 | ~v_3108;
assign x_13363 = v_3229 | ~v_18;
assign x_13364 = v_3229 | ~v_17;
assign x_13365 = v_3229 | ~v_15;
assign x_13366 = v_3229 | ~v_12;
assign x_13367 = ~v_3227 | ~v_3226 | ~v_3225 | v_3228;
assign x_13368 = v_3227 | ~v_1073;
assign x_13369 = v_3227 | ~v_1074;
assign x_13370 = v_3227 | ~v_1075;
assign x_13371 = v_3227 | ~v_1076;
assign x_13372 = v_3227 | ~v_919;
assign x_13373 = v_3227 | ~v_920;
assign x_13374 = v_3227 | ~v_3125;
assign x_13375 = v_3227 | ~v_3126;
assign x_13376 = v_3227 | ~v_817;
assign x_13377 = v_3227 | ~v_3127;
assign x_13378 = v_3227 | ~v_3128;
assign x_13379 = v_3227 | ~v_820;
assign x_13380 = v_3227 | ~v_3167;
assign x_13381 = v_3227 | ~v_3168;
assign x_13382 = v_3227 | ~v_927;
assign x_13383 = v_3227 | ~v_3169;
assign x_13384 = v_3227 | ~v_3170;
assign x_13385 = v_3227 | ~v_928;
assign x_13386 = v_3227 | ~v_1099;
assign x_13387 = v_3227 | ~v_1100;
assign x_13388 = v_3227 | ~v_1101;
assign x_13389 = v_3227 | ~v_1102;
assign x_13390 = v_3227 | ~v_3219;
assign x_13391 = v_3227 | ~v_3220;
assign x_13392 = v_3227 | ~v_1085;
assign x_13393 = v_3227 | ~v_3221;
assign x_13394 = v_3227 | ~v_3222;
assign x_13395 = v_3227 | ~v_1086;
assign x_13396 = v_3227 | ~v_3133;
assign x_13397 = v_3227 | ~v_3136;
assign x_13398 = v_3227 | ~v_931;
assign x_13399 = v_3227 | ~v_932;
assign x_13400 = v_3227 | ~v_184;
assign x_13401 = v_3227 | ~v_171;
assign x_13402 = v_3227 | ~v_170;
assign x_13403 = v_3227 | ~v_169;
assign x_13404 = v_3227 | ~v_150;
assign x_13405 = v_3227 | ~v_149;
assign x_13406 = v_3227 | ~v_148;
assign x_13407 = v_3227 | ~v_103;
assign x_13408 = v_3227 | ~v_102;
assign x_13409 = v_3227 | ~v_101;
assign x_13410 = v_3227 | ~v_100;
assign x_13411 = v_3227 | ~v_95;
assign x_13412 = v_3226 | ~v_1058;
assign x_13413 = v_3226 | ~v_1059;
assign x_13414 = v_3226 | ~v_1060;
assign x_13415 = v_3226 | ~v_1061;
assign x_13416 = v_3226 | ~v_904;
assign x_13417 = v_3226 | ~v_905;
assign x_13418 = v_3226 | ~v_3110;
assign x_13419 = v_3226 | ~v_3111;
assign x_13420 = v_3226 | ~v_784;
assign x_13421 = v_3226 | ~v_3112;
assign x_13422 = v_3226 | ~v_3113;
assign x_13423 = v_3226 | ~v_787;
assign x_13424 = v_3226 | ~v_3162;
assign x_13425 = v_3226 | ~v_3163;
assign x_13426 = v_3226 | ~v_912;
assign x_13427 = v_3226 | ~v_3164;
assign x_13428 = v_3226 | ~v_3165;
assign x_13429 = v_3226 | ~v_913;
assign x_13430 = v_3226 | ~v_1094;
assign x_13431 = v_3226 | ~v_1095;
assign x_13432 = v_3226 | ~v_1096;
assign x_13433 = v_3226 | ~v_1097;
assign x_13434 = v_3226 | ~v_3214;
assign x_13435 = v_3226 | ~v_3215;
assign x_13436 = v_3226 | ~v_1070;
assign x_13437 = v_3226 | ~v_3216;
assign x_13438 = v_3226 | ~v_3217;
assign x_13439 = v_3226 | ~v_1071;
assign x_13440 = v_3226 | ~v_3118;
assign x_13441 = v_3226 | ~v_3121;
assign x_13442 = v_3226 | ~v_916;
assign x_13443 = v_3226 | ~v_917;
assign x_13444 = v_3226 | ~v_183;
assign x_13445 = v_3226 | ~v_167;
assign x_13446 = v_3226 | ~v_166;
assign x_13447 = v_3226 | ~v_165;
assign x_13448 = v_3226 | ~v_145;
assign x_13449 = v_3226 | ~v_144;
assign x_13450 = v_3226 | ~v_143;
assign x_13451 = v_3226 | ~v_61;
assign x_13452 = v_3226 | ~v_60;
assign x_13453 = v_3226 | ~v_59;
assign x_13454 = v_3226 | ~v_58;
assign x_13455 = v_3226 | ~v_53;
assign x_13456 = v_3225 | ~v_1043;
assign x_13457 = v_3225 | ~v_1044;
assign x_13458 = v_3225 | ~v_1045;
assign x_13459 = v_3225 | ~v_1046;
assign x_13460 = v_3225 | ~v_889;
assign x_13461 = v_3225 | ~v_890;
assign x_13462 = v_3225 | ~v_3095;
assign x_13463 = v_3225 | ~v_3096;
assign x_13464 = v_3225 | ~v_751;
assign x_13465 = v_3225 | ~v_3097;
assign x_13466 = v_3225 | ~v_3098;
assign x_13467 = v_3225 | ~v_754;
assign x_13468 = v_3225 | ~v_3157;
assign x_13469 = v_3225 | ~v_3158;
assign x_13470 = v_3225 | ~v_897;
assign x_13471 = v_3225 | ~v_3159;
assign x_13472 = v_3225 | ~v_3160;
assign x_13473 = v_3225 | ~v_898;
assign x_13474 = v_3225 | ~v_1089;
assign x_13475 = v_3225 | ~v_1090;
assign x_13476 = v_3225 | ~v_1091;
assign x_13477 = v_3225 | ~v_1092;
assign x_13478 = v_3225 | ~v_3209;
assign x_13479 = v_3225 | ~v_3210;
assign x_13480 = v_3225 | ~v_1055;
assign x_13481 = v_3225 | ~v_3211;
assign x_13482 = v_3225 | ~v_3212;
assign x_13483 = v_3225 | ~v_1056;
assign x_13484 = v_3225 | ~v_901;
assign x_13485 = v_3225 | ~v_902;
assign x_13486 = v_3225 | ~v_182;
assign x_13487 = v_3225 | ~v_163;
assign x_13488 = v_3225 | ~v_162;
assign x_13489 = v_3225 | ~v_161;
assign x_13490 = v_3225 | ~v_137;
assign x_13491 = v_3225 | ~v_136;
assign x_13492 = v_3225 | ~v_135;
assign x_13493 = v_3225 | ~v_3107;
assign x_13494 = v_3225 | ~v_3108;
assign x_13495 = v_3225 | ~v_18;
assign x_13496 = v_3225 | ~v_17;
assign x_13497 = v_3225 | ~v_16;
assign x_13498 = v_3225 | ~v_15;
assign x_13499 = v_3225 | ~v_10;
assign x_13500 = ~v_3223 | ~v_3218 | ~v_3213 | v_3224;
assign x_13501 = v_3223 | ~v_1073;
assign x_13502 = v_3223 | ~v_1074;
assign x_13503 = v_3223 | ~v_1075;
assign x_13504 = v_3223 | ~v_1076;
assign x_13505 = v_3223 | ~v_965;
assign x_13506 = v_3223 | ~v_966;
assign x_13507 = v_3223 | ~v_967;
assign x_13508 = v_3223 | ~v_968;
assign x_13509 = v_3223 | ~v_3125;
assign x_13510 = v_3223 | ~v_3126;
assign x_13511 = v_3223 | ~v_817;
assign x_13512 = v_3223 | ~v_3127;
assign x_13513 = v_3223 | ~v_3128;
assign x_13514 = v_3223 | ~v_820;
assign x_13515 = v_3223 | ~v_3129;
assign x_13516 = v_3223 | ~v_3130;
assign x_13517 = v_3223 | ~v_975;
assign x_13518 = v_3223 | ~v_3131;
assign x_13519 = v_3223 | ~v_3132;
assign x_13520 = v_3223 | ~v_976;
assign x_13521 = v_3223 | ~v_1115;
assign x_13522 = v_3223 | ~v_1116;
assign x_13523 = v_3223 | ~v_3219;
assign x_13524 = v_3223 | ~v_3220;
assign x_13525 = v_3223 | ~v_1085;
assign x_13526 = v_3223 | ~v_3221;
assign x_13527 = v_3223 | ~v_3222;
assign x_13528 = v_3223 | ~v_1086;
assign x_13529 = v_3223 | ~v_3133;
assign x_13530 = v_3223 | ~v_3136;
assign x_13531 = v_3223 | ~v_1117;
assign x_13532 = v_3223 | ~v_1118;
assign x_13533 = v_3223 | ~v_184;
assign x_13534 = v_3223 | ~v_171;
assign x_13535 = v_3223 | ~v_170;
assign x_13536 = v_3223 | ~v_169;
assign x_13537 = v_3223 | ~v_151;
assign x_13538 = v_3223 | ~v_150;
assign x_13539 = v_3223 | ~v_149;
assign x_13540 = v_3223 | ~v_148;
assign x_13541 = v_3223 | ~v_147;
assign x_13542 = v_3223 | ~v_103;
assign x_13543 = v_3223 | ~v_101;
assign x_13544 = v_3223 | ~v_100;
assign x_13545 = ~v_127 | ~v_140 | v_3222;
assign x_13546 = ~v_121 | ~v_139 | v_3221;
assign x_13547 = ~v_112 | v_140 | v_3220;
assign x_13548 = ~v_106 | v_139 | v_3219;
assign x_13549 = v_3218 | ~v_1058;
assign x_13550 = v_3218 | ~v_1059;
assign x_13551 = v_3218 | ~v_1060;
assign x_13552 = v_3218 | ~v_1061;
assign x_13553 = v_3218 | ~v_950;
assign x_13554 = v_3218 | ~v_951;
assign x_13555 = v_3218 | ~v_952;
assign x_13556 = v_3218 | ~v_953;
assign x_13557 = v_3218 | ~v_3110;
assign x_13558 = v_3218 | ~v_3111;
assign x_13559 = v_3218 | ~v_784;
assign x_13560 = v_3218 | ~v_3112;
assign x_13561 = v_3218 | ~v_3113;
assign x_13562 = v_3218 | ~v_787;
assign x_13563 = v_3218 | ~v_3114;
assign x_13564 = v_3218 | ~v_3115;
assign x_13565 = v_3218 | ~v_960;
assign x_13566 = v_3218 | ~v_3116;
assign x_13567 = v_3218 | ~v_3117;
assign x_13568 = v_3218 | ~v_961;
assign x_13569 = v_3218 | ~v_1110;
assign x_13570 = v_3218 | ~v_1111;
assign x_13571 = v_3218 | ~v_3214;
assign x_13572 = v_3218 | ~v_3215;
assign x_13573 = v_3218 | ~v_1070;
assign x_13574 = v_3218 | ~v_3216;
assign x_13575 = v_3218 | ~v_3217;
assign x_13576 = v_3218 | ~v_1071;
assign x_13577 = v_3218 | ~v_3118;
assign x_13578 = v_3218 | ~v_3121;
assign x_13579 = v_3218 | ~v_1112;
assign x_13580 = v_3218 | ~v_1113;
assign x_13581 = v_3218 | ~v_183;
assign x_13582 = v_3218 | ~v_167;
assign x_13583 = v_3218 | ~v_166;
assign x_13584 = v_3218 | ~v_165;
assign x_13585 = v_3218 | ~v_146;
assign x_13586 = v_3218 | ~v_145;
assign x_13587 = v_3218 | ~v_144;
assign x_13588 = v_3218 | ~v_143;
assign x_13589 = v_3218 | ~v_142;
assign x_13590 = v_3218 | ~v_61;
assign x_13591 = v_3218 | ~v_59;
assign x_13592 = v_3218 | ~v_58;
assign x_13593 = ~v_85 | ~v_140 | v_3217;
assign x_13594 = ~v_79 | ~v_139 | v_3216;
assign x_13595 = ~v_70 | v_140 | v_3215;
assign x_13596 = ~v_64 | v_139 | v_3214;
assign x_13597 = v_3213 | ~v_1043;
assign x_13598 = v_3213 | ~v_1044;
assign x_13599 = v_3213 | ~v_1045;
assign x_13600 = v_3213 | ~v_1046;
assign x_13601 = v_3213 | ~v_935;
assign x_13602 = v_3213 | ~v_936;
assign x_13603 = v_3213 | ~v_937;
assign x_13604 = v_3213 | ~v_938;
assign x_13605 = v_3213 | ~v_3095;
assign x_13606 = v_3213 | ~v_3096;
assign x_13607 = v_3213 | ~v_751;
assign x_13608 = v_3213 | ~v_3097;
assign x_13609 = v_3213 | ~v_3098;
assign x_13610 = v_3213 | ~v_754;
assign x_13611 = v_3213 | ~v_3099;
assign x_13612 = v_3213 | ~v_3100;
assign x_13613 = v_3213 | ~v_945;
assign x_13614 = v_3213 | ~v_3101;
assign x_13615 = v_3213 | ~v_3102;
assign x_13616 = v_3213 | ~v_946;
assign x_13617 = v_3213 | ~v_1105;
assign x_13618 = v_3213 | ~v_1106;
assign x_13619 = v_3213 | ~v_3209;
assign x_13620 = v_3213 | ~v_3210;
assign x_13621 = v_3213 | ~v_1055;
assign x_13622 = v_3213 | ~v_3211;
assign x_13623 = v_3213 | ~v_3212;
assign x_13624 = v_3213 | ~v_1056;
assign x_13625 = v_3213 | ~v_1107;
assign x_13626 = v_3213 | ~v_1108;
assign x_13627 = v_3213 | ~v_182;
assign x_13628 = v_3213 | ~v_163;
assign x_13629 = v_3213 | ~v_162;
assign x_13630 = v_3213 | ~v_161;
assign x_13631 = v_3213 | ~v_138;
assign x_13632 = v_3213 | ~v_137;
assign x_13633 = v_3213 | ~v_136;
assign x_13634 = v_3213 | ~v_135;
assign x_13635 = v_3213 | ~v_134;
assign x_13636 = v_3213 | ~v_3107;
assign x_13637 = v_3213 | ~v_3108;
assign x_13638 = v_3213 | ~v_18;
assign x_13639 = v_3213 | ~v_16;
assign x_13640 = v_3213 | ~v_15;
assign x_13641 = ~v_43 | ~v_140 | v_3212;
assign x_13642 = ~v_37 | ~v_139 | v_3211;
assign x_13643 = ~v_28 | v_140 | v_3210;
assign x_13644 = ~v_22 | v_139 | v_3209;
assign x_13645 = ~v_3207 | ~v_3206 | ~v_3205 | v_3208;
assign x_13646 = v_3207 | ~v_919;
assign x_13647 = v_3207 | ~v_920;
assign x_13648 = v_3207 | ~v_3125;
assign x_13649 = v_3207 | ~v_3126;
assign x_13650 = v_3207 | ~v_817;
assign x_13651 = v_3207 | ~v_818;
assign x_13652 = v_3207 | ~v_819;
assign x_13653 = v_3207 | ~v_3127;
assign x_13654 = v_3207 | ~v_3128;
assign x_13655 = v_3207 | ~v_820;
assign x_13656 = v_3207 | ~v_821;
assign x_13657 = v_3207 | ~v_822;
assign x_13658 = v_3207 | ~v_1037;
assign x_13659 = v_3207 | ~v_1038;
assign x_13660 = v_3207 | ~v_1039;
assign x_13661 = v_3207 | ~v_1040;
assign x_13662 = v_3207 | ~v_3167;
assign x_13663 = v_3207 | ~v_3168;
assign x_13664 = v_3207 | ~v_927;
assign x_13665 = v_3207 | ~v_3169;
assign x_13666 = v_3207 | ~v_3170;
assign x_13667 = v_3207 | ~v_928;
assign x_13668 = v_3207 | ~v_3133;
assign x_13669 = v_3207 | ~v_3134;
assign x_13670 = v_3207 | ~v_3135;
assign x_13671 = v_3207 | ~v_839;
assign x_13672 = v_3207 | ~v_3136;
assign x_13673 = v_3207 | ~v_3137;
assign x_13674 = v_3207 | ~v_3138;
assign x_13675 = v_3207 | ~v_840;
assign x_13676 = v_3207 | ~v_931;
assign x_13677 = v_3207 | ~v_932;
assign x_13678 = v_3207 | ~v_184;
assign x_13679 = v_3207 | ~v_170;
assign x_13680 = v_3207 | ~v_151;
assign x_13681 = v_3207 | ~v_150;
assign x_13682 = v_3207 | ~v_149;
assign x_13683 = v_3207 | ~v_148;
assign x_13684 = v_3207 | ~v_147;
assign x_13685 = v_3207 | ~v_103;
assign x_13686 = v_3207 | ~v_101;
assign x_13687 = v_3207 | ~v_100;
assign x_13688 = v_3207 | ~v_98;
assign x_13689 = v_3207 | ~v_93;
assign x_13690 = v_3206 | ~v_904;
assign x_13691 = v_3206 | ~v_905;
assign x_13692 = v_3206 | ~v_3110;
assign x_13693 = v_3206 | ~v_3111;
assign x_13694 = v_3206 | ~v_784;
assign x_13695 = v_3206 | ~v_785;
assign x_13696 = v_3206 | ~v_786;
assign x_13697 = v_3206 | ~v_3112;
assign x_13698 = v_3206 | ~v_3113;
assign x_13699 = v_3206 | ~v_787;
assign x_13700 = v_3206 | ~v_788;
assign x_13701 = v_3206 | ~v_789;
assign x_13702 = v_3206 | ~v_1032;
assign x_13703 = v_3206 | ~v_1033;
assign x_13704 = v_3206 | ~v_1034;
assign x_13705 = v_3206 | ~v_1035;
assign x_13706 = v_3206 | ~v_3162;
assign x_13707 = v_3206 | ~v_3163;
assign x_13708 = v_3206 | ~v_912;
assign x_13709 = v_3206 | ~v_3164;
assign x_13710 = v_3206 | ~v_3165;
assign x_13711 = v_3206 | ~v_913;
assign x_13712 = v_3206 | ~v_3118;
assign x_13713 = v_3206 | ~v_3119;
assign x_13714 = v_3206 | ~v_3120;
assign x_13715 = v_3206 | ~v_806;
assign x_13716 = v_3206 | ~v_3121;
assign x_13717 = v_3206 | ~v_3122;
assign x_13718 = v_3206 | ~v_3123;
assign x_13719 = v_3206 | ~v_807;
assign x_13720 = v_3206 | ~v_916;
assign x_13721 = v_3206 | ~v_917;
assign x_13722 = v_3206 | ~v_183;
assign x_13723 = v_3206 | ~v_166;
assign x_13724 = v_3206 | ~v_146;
assign x_13725 = v_3206 | ~v_145;
assign x_13726 = v_3206 | ~v_144;
assign x_13727 = v_3206 | ~v_143;
assign x_13728 = v_3206 | ~v_142;
assign x_13729 = v_3206 | ~v_61;
assign x_13730 = v_3206 | ~v_59;
assign x_13731 = v_3206 | ~v_58;
assign x_13732 = v_3206 | ~v_56;
assign x_13733 = v_3206 | ~v_51;
assign x_13734 = v_3205 | ~v_889;
assign x_13735 = v_3205 | ~v_890;
assign x_13736 = v_3205 | ~v_3095;
assign x_13737 = v_3205 | ~v_3096;
assign x_13738 = v_3205 | ~v_751;
assign x_13739 = v_3205 | ~v_752;
assign x_13740 = v_3205 | ~v_753;
assign x_13741 = v_3205 | ~v_3097;
assign x_13742 = v_3205 | ~v_3098;
assign x_13743 = v_3205 | ~v_754;
assign x_13744 = v_3205 | ~v_755;
assign x_13745 = v_3205 | ~v_756;
assign x_13746 = v_3205 | ~v_1027;
assign x_13747 = v_3205 | ~v_1028;
assign x_13748 = v_3205 | ~v_1029;
assign x_13749 = v_3205 | ~v_1030;
assign x_13750 = v_3205 | ~v_3157;
assign x_13751 = v_3205 | ~v_3158;
assign x_13752 = v_3205 | ~v_897;
assign x_13753 = v_3205 | ~v_3159;
assign x_13754 = v_3205 | ~v_3160;
assign x_13755 = v_3205 | ~v_898;
assign x_13756 = v_3205 | ~v_3103;
assign x_13757 = v_3205 | ~v_3104;
assign x_13758 = v_3205 | ~v_773;
assign x_13759 = v_3205 | ~v_3105;
assign x_13760 = v_3205 | ~v_3106;
assign x_13761 = v_3205 | ~v_774;
assign x_13762 = v_3205 | ~v_901;
assign x_13763 = v_3205 | ~v_902;
assign x_13764 = v_3205 | ~v_182;
assign x_13765 = v_3205 | ~v_162;
assign x_13766 = v_3205 | ~v_138;
assign x_13767 = v_3205 | ~v_137;
assign x_13768 = v_3205 | ~v_136;
assign x_13769 = v_3205 | ~v_135;
assign x_13770 = v_3205 | ~v_134;
assign x_13771 = v_3205 | ~v_3107;
assign x_13772 = v_3205 | ~v_3108;
assign x_13773 = v_3205 | ~v_18;
assign x_13774 = v_3205 | ~v_16;
assign x_13775 = v_3205 | ~v_15;
assign x_13776 = v_3205 | ~v_13;
assign x_13777 = v_3205 | ~v_8;
assign x_13778 = ~v_3203 | ~v_3198 | ~v_3193 | v_3204;
assign x_13779 = v_3203 | ~v_1183;
assign x_13780 = v_3203 | ~v_1184;
assign x_13781 = v_3203 | ~v_1185;
assign x_13782 = v_3203 | ~v_1186;
assign x_13783 = v_3203 | ~v_3125;
assign x_13784 = v_3203 | ~v_3126;
assign x_13785 = v_3203 | ~v_817;
assign x_13786 = v_3203 | ~v_1011;
assign x_13787 = v_3203 | ~v_1012;
assign x_13788 = v_3203 | ~v_3127;
assign x_13789 = v_3203 | ~v_3128;
assign x_13790 = v_3203 | ~v_820;
assign x_13791 = v_3203 | ~v_1013;
assign x_13792 = v_3203 | ~v_1014;
assign x_13793 = v_3203 | ~v_3151;
assign x_13794 = v_3203 | ~v_3152;
assign x_13795 = v_3203 | ~v_1193;
assign x_13796 = v_3203 | ~v_1241;
assign x_13797 = v_3203 | ~v_3153;
assign x_13798 = v_3203 | ~v_3154;
assign x_13799 = v_3203 | ~v_1194;
assign x_13800 = v_3203 | ~v_1242;
assign x_13801 = v_3203 | ~v_3133;
assign x_13802 = v_3203 | ~v_3199;
assign x_13803 = v_3203 | ~v_3200;
assign x_13804 = v_3203 | ~v_1023;
assign x_13805 = v_3203 | ~v_3136;
assign x_13806 = v_3203 | ~v_3201;
assign x_13807 = v_3203 | ~v_3202;
assign x_13808 = v_3203 | ~v_1024;
assign x_13809 = v_3203 | ~v_1243;
assign x_13810 = v_3203 | ~v_1244;
assign x_13811 = v_3203 | ~v_184;
assign x_13812 = v_3203 | ~v_171;
assign x_13813 = v_3203 | ~v_170;
assign x_13814 = v_3203 | ~v_169;
assign x_13815 = v_3203 | ~v_149;
assign x_13816 = v_3203 | ~v_147;
assign x_13817 = v_3203 | ~v_103;
assign x_13818 = v_3203 | ~v_102;
assign x_13819 = v_3203 | ~v_101;
assign x_13820 = v_3203 | ~v_100;
assign x_13821 = v_3203 | ~v_99;
assign x_13822 = v_3203 | ~v_96;
assign x_13823 = ~v_19 | ~v_130 | v_3202;
assign x_13824 = ~v_19 | ~v_122 | v_3201;
assign x_13825 = v_19 | ~v_115 | v_3200;
assign x_13826 = v_19 | ~v_107 | v_3199;
assign x_13827 = v_3198 | ~v_1168;
assign x_13828 = v_3198 | ~v_1169;
assign x_13829 = v_3198 | ~v_1170;
assign x_13830 = v_3198 | ~v_1171;
assign x_13831 = v_3198 | ~v_3110;
assign x_13832 = v_3198 | ~v_3111;
assign x_13833 = v_3198 | ~v_784;
assign x_13834 = v_3198 | ~v_996;
assign x_13835 = v_3198 | ~v_997;
assign x_13836 = v_3198 | ~v_3112;
assign x_13837 = v_3198 | ~v_3113;
assign x_13838 = v_3198 | ~v_787;
assign x_13839 = v_3198 | ~v_998;
assign x_13840 = v_3198 | ~v_999;
assign x_13841 = v_3198 | ~v_3146;
assign x_13842 = v_3198 | ~v_3147;
assign x_13843 = v_3198 | ~v_1178;
assign x_13844 = v_3198 | ~v_1236;
assign x_13845 = v_3198 | ~v_3148;
assign x_13846 = v_3198 | ~v_3149;
assign x_13847 = v_3198 | ~v_1179;
assign x_13848 = v_3198 | ~v_1237;
assign x_13849 = v_3198 | ~v_3118;
assign x_13850 = v_3198 | ~v_3194;
assign x_13851 = v_3198 | ~v_3195;
assign x_13852 = v_3198 | ~v_1008;
assign x_13853 = v_3198 | ~v_3121;
assign x_13854 = v_3198 | ~v_1009;
assign x_13855 = v_3198 | ~v_3196;
assign x_13856 = v_3198 | ~v_1238;
assign x_13857 = v_3198 | ~v_1239;
assign x_13858 = v_3198 | ~v_183;
assign x_13859 = v_3198 | ~v_167;
assign x_13860 = v_3198 | ~v_166;
assign x_13861 = v_3198 | ~v_165;
assign x_13862 = v_3198 | ~v_144;
assign x_13863 = v_3198 | ~v_142;
assign x_13864 = v_3198 | ~v_3197;
assign x_13865 = v_3198 | ~v_61;
assign x_13866 = v_3198 | ~v_60;
assign x_13867 = v_3198 | ~v_59;
assign x_13868 = v_3198 | ~v_58;
assign x_13869 = v_3198 | ~v_57;
assign x_13870 = v_3198 | ~v_54;
assign x_13871 = ~v_19 | ~v_80 | v_3197;
assign x_13872 = ~v_19 | ~v_88 | v_3196;
assign x_13873 = v_19 | ~v_73 | v_3195;
assign x_13874 = v_19 | ~v_65 | v_3194;
assign x_13875 = v_3193 | ~v_1153;
assign x_13876 = v_3193 | ~v_1154;
assign x_13877 = v_3193 | ~v_1155;
assign x_13878 = v_3193 | ~v_1156;
assign x_13879 = v_3193 | ~v_3095;
assign x_13880 = v_3193 | ~v_3096;
assign x_13881 = v_3193 | ~v_751;
assign x_13882 = v_3193 | ~v_981;
assign x_13883 = v_3193 | ~v_982;
assign x_13884 = v_3193 | ~v_3097;
assign x_13885 = v_3193 | ~v_3098;
assign x_13886 = v_3193 | ~v_754;
assign x_13887 = v_3193 | ~v_983;
assign x_13888 = v_3193 | ~v_984;
assign x_13889 = v_3193 | ~v_3141;
assign x_13890 = v_3193 | ~v_3142;
assign x_13891 = v_3193 | ~v_1163;
assign x_13892 = v_3193 | ~v_1231;
assign x_13893 = v_3193 | ~v_3143;
assign x_13894 = v_3193 | ~v_3144;
assign x_13895 = v_3193 | ~v_1164;
assign x_13896 = v_3193 | ~v_1232;
assign x_13897 = v_3193 | ~v_3189;
assign x_13898 = v_3193 | ~v_3190;
assign x_13899 = v_3193 | ~v_3191;
assign x_13900 = v_3193 | ~v_3192;
assign x_13901 = v_3193 | ~v_1233;
assign x_13902 = v_3193 | ~v_1234;
assign x_13903 = v_3193 | ~v_182;
assign x_13904 = v_3193 | ~v_163;
assign x_13905 = v_3193 | ~v_162;
assign x_13906 = v_3193 | ~v_161;
assign x_13907 = v_3193 | ~v_136;
assign x_13908 = v_3193 | ~v_134;
assign x_13909 = v_3193 | ~v_3107;
assign x_13910 = v_3193 | ~v_993;
assign x_13911 = v_3193 | ~v_3108;
assign x_13912 = v_3193 | ~v_994;
assign x_13913 = v_3193 | ~v_18;
assign x_13914 = v_3193 | ~v_17;
assign x_13915 = v_3193 | ~v_16;
assign x_13916 = v_3193 | ~v_15;
assign x_13917 = v_3193 | ~v_14;
assign x_13918 = v_3193 | ~v_11;
assign x_13919 = ~v_19 | ~v_46 | v_3192;
assign x_13920 = ~v_19 | ~v_38 | v_3191;
assign x_13921 = ~v_31 | v_19 | v_3190;
assign x_13922 = ~v_23 | v_19 | v_3189;
assign x_13923 = ~v_3187 | ~v_3182 | ~v_3177 | v_3188;
assign x_13924 = v_3187 | ~v_1183;
assign x_13925 = v_3187 | ~v_1184;
assign x_13926 = v_3187 | ~v_1185;
assign x_13927 = v_3187 | ~v_1186;
assign x_13928 = v_3187 | ~v_813;
assign x_13929 = v_3187 | ~v_814;
assign x_13930 = v_3187 | ~v_815;
assign x_13931 = v_3187 | ~v_816;
assign x_13932 = v_3187 | ~v_3125;
assign x_13933 = v_3187 | ~v_3126;
assign x_13934 = v_3187 | ~v_817;
assign x_13935 = v_3187 | ~v_3127;
assign x_13936 = v_3187 | ~v_3128;
assign x_13937 = v_3187 | ~v_820;
assign x_13938 = v_3187 | ~v_1191;
assign x_13939 = v_3187 | ~v_1192;
assign x_13940 = v_3187 | ~v_3151;
assign x_13941 = v_3187 | ~v_3152;
assign x_13942 = v_3187 | ~v_1193;
assign x_13943 = v_3187 | ~v_3153;
assign x_13944 = v_3187 | ~v_3154;
assign x_13945 = v_3187 | ~v_1194;
assign x_13946 = v_3187 | ~v_3183;
assign x_13947 = v_3187 | ~v_3184;
assign x_13948 = v_3187 | ~v_837;
assign x_13949 = v_3187 | ~v_3185;
assign x_13950 = v_3187 | ~v_3186;
assign x_13951 = v_3187 | ~v_838;
assign x_13952 = v_3187 | ~v_3133;
assign x_13953 = v_3187 | ~v_3136;
assign x_13954 = v_3187 | ~v_1195;
assign x_13955 = v_3187 | ~v_1196;
assign x_13956 = v_3187 | ~v_184;
assign x_13957 = v_3187 | ~v_171;
assign x_13958 = v_3187 | ~v_170;
assign x_13959 = v_3187 | ~v_169;
assign x_13960 = v_3187 | ~v_160;
assign x_13961 = v_3187 | ~v_151;
assign x_13962 = v_3187 | ~v_150;
assign x_13963 = v_3187 | ~v_148;
assign x_13964 = v_3187 | ~v_147;
assign x_13965 = v_3187 | ~v_103;
assign x_13966 = v_3187 | ~v_100;
assign x_13967 = v_3187 | ~v_97;
assign x_13968 = ~v_130 | ~v_157 | v_3186;
assign x_13969 = ~v_122 | ~v_156 | v_3185;
assign x_13970 = ~v_115 | v_157 | v_3184;
assign x_13971 = ~v_107 | v_156 | v_3183;
assign x_13972 = v_3182 | ~v_1168;
assign x_13973 = v_3182 | ~v_1169;
assign x_13974 = v_3182 | ~v_1170;
assign x_13975 = v_3182 | ~v_1171;
assign x_13976 = v_3182 | ~v_780;
assign x_13977 = v_3182 | ~v_781;
assign x_13978 = v_3182 | ~v_782;
assign x_13979 = v_3182 | ~v_783;
assign x_13980 = v_3182 | ~v_3110;
assign x_13981 = v_3182 | ~v_3111;
assign x_13982 = v_3182 | ~v_784;
assign x_13983 = v_3182 | ~v_3112;
assign x_13984 = v_3182 | ~v_3113;
assign x_13985 = v_3182 | ~v_787;
assign x_13986 = v_3182 | ~v_1176;
assign x_13987 = v_3182 | ~v_1177;
assign x_13988 = v_3182 | ~v_3146;
assign x_13989 = v_3182 | ~v_3147;
assign x_13990 = v_3182 | ~v_1178;
assign x_13991 = v_3182 | ~v_3148;
assign x_13992 = v_3182 | ~v_3149;
assign x_13993 = v_3182 | ~v_1179;
assign x_13994 = v_3182 | ~v_3178;
assign x_13995 = v_3182 | ~v_3179;
assign x_13996 = v_3182 | ~v_804;
assign x_13997 = v_3182 | ~v_3180;
assign x_13998 = v_3182 | ~v_3181;
assign x_13999 = v_3182 | ~v_805;
assign x_14000 = v_3182 | ~v_3118;
assign x_14001 = v_3182 | ~v_3121;
assign x_14002 = v_3182 | ~v_1180;
assign x_14003 = v_3182 | ~v_1181;
assign x_14004 = v_3182 | ~v_183;
assign x_14005 = v_3182 | ~v_167;
assign x_14006 = v_3182 | ~v_166;
assign x_14007 = v_3182 | ~v_165;
assign x_14008 = v_3182 | ~v_159;
assign x_14009 = v_3182 | ~v_146;
assign x_14010 = v_3182 | ~v_145;
assign x_14011 = v_3182 | ~v_143;
assign x_14012 = v_3182 | ~v_142;
assign x_14013 = v_3182 | ~v_61;
assign x_14014 = v_3182 | ~v_58;
assign x_14015 = v_3182 | ~v_55;
assign x_14016 = ~v_88 | ~v_157 | v_3181;
assign x_14017 = ~v_80 | ~v_156 | v_3180;
assign x_14018 = ~v_73 | v_157 | v_3179;
assign x_14019 = ~v_65 | v_156 | v_3178;
assign x_14020 = v_3177 | ~v_1153;
assign x_14021 = v_3177 | ~v_1154;
assign x_14022 = v_3177 | ~v_1155;
assign x_14023 = v_3177 | ~v_1156;
assign x_14024 = v_3177 | ~v_747;
assign x_14025 = v_3177 | ~v_748;
assign x_14026 = v_3177 | ~v_749;
assign x_14027 = v_3177 | ~v_750;
assign x_14028 = v_3177 | ~v_3095;
assign x_14029 = v_3177 | ~v_3096;
assign x_14030 = v_3177 | ~v_751;
assign x_14031 = v_3177 | ~v_3097;
assign x_14032 = v_3177 | ~v_3098;
assign x_14033 = v_3177 | ~v_754;
assign x_14034 = v_3177 | ~v_1161;
assign x_14035 = v_3177 | ~v_1162;
assign x_14036 = v_3177 | ~v_3141;
assign x_14037 = v_3177 | ~v_3142;
assign x_14038 = v_3177 | ~v_1163;
assign x_14039 = v_3177 | ~v_3143;
assign x_14040 = v_3177 | ~v_3144;
assign x_14041 = v_3177 | ~v_1164;
assign x_14042 = v_3177 | ~v_3173;
assign x_14043 = v_3177 | ~v_3174;
assign x_14044 = v_3177 | ~v_771;
assign x_14045 = v_3177 | ~v_3175;
assign x_14046 = v_3177 | ~v_3176;
assign x_14047 = v_3177 | ~v_772;
assign x_14048 = v_3177 | ~v_1165;
assign x_14049 = v_3177 | ~v_1166;
assign x_14050 = v_3177 | ~v_182;
assign x_14051 = v_3177 | ~v_163;
assign x_14052 = v_3177 | ~v_162;
assign x_14053 = v_3177 | ~v_161;
assign x_14054 = v_3177 | ~v_155;
assign x_14055 = v_3177 | ~v_138;
assign x_14056 = v_3177 | ~v_137;
assign x_14057 = v_3177 | ~v_135;
assign x_14058 = v_3177 | ~v_134;
assign x_14059 = v_3177 | ~v_3107;
assign x_14060 = v_3177 | ~v_3108;
assign x_14061 = v_3177 | ~v_18;
assign x_14062 = v_3177 | ~v_15;
assign x_14063 = v_3177 | ~v_12;
assign x_14064 = ~v_46 | ~v_157 | v_3176;
assign x_14065 = ~v_38 | ~v_156 | v_3175;
assign x_14066 = ~v_31 | v_157 | v_3174;
assign x_14067 = ~v_23 | v_156 | v_3173;
assign x_14068 = ~v_3171 | ~v_3166 | ~v_3161 | v_3172;
assign x_14069 = v_3171 | ~v_1183;
assign x_14070 = v_3171 | ~v_1184;
assign x_14071 = v_3171 | ~v_1185;
assign x_14072 = v_3171 | ~v_1186;
assign x_14073 = v_3171 | ~v_919;
assign x_14074 = v_3171 | ~v_920;
assign x_14075 = v_3171 | ~v_3125;
assign x_14076 = v_3171 | ~v_3126;
assign x_14077 = v_3171 | ~v_817;
assign x_14078 = v_3171 | ~v_3127;
assign x_14079 = v_3171 | ~v_3128;
assign x_14080 = v_3171 | ~v_820;
assign x_14081 = v_3171 | ~v_1209;
assign x_14082 = v_3171 | ~v_1210;
assign x_14083 = v_3171 | ~v_3151;
assign x_14084 = v_3171 | ~v_3152;
assign x_14085 = v_3171 | ~v_1193;
assign x_14086 = v_3171 | ~v_3153;
assign x_14087 = v_3171 | ~v_3154;
assign x_14088 = v_3171 | ~v_1194;
assign x_14089 = v_3171 | ~v_3167;
assign x_14090 = v_3171 | ~v_3168;
assign x_14091 = v_3171 | ~v_927;
assign x_14092 = v_3171 | ~v_3169;
assign x_14093 = v_3171 | ~v_3170;
assign x_14094 = v_3171 | ~v_928;
assign x_14095 = v_3171 | ~v_3133;
assign x_14096 = v_3171 | ~v_3136;
assign x_14097 = v_3171 | ~v_931;
assign x_14098 = v_3171 | ~v_932;
assign x_14099 = v_3171 | ~v_1211;
assign x_14100 = v_3171 | ~v_1212;
assign x_14101 = v_3171 | ~v_184;
assign x_14102 = v_3171 | ~v_172;
assign x_14103 = v_3171 | ~v_171;
assign x_14104 = v_3171 | ~v_170;
assign x_14105 = v_3171 | ~v_169;
assign x_14106 = v_3171 | ~v_150;
assign x_14107 = v_3171 | ~v_149;
assign x_14108 = v_3171 | ~v_148;
assign x_14109 = v_3171 | ~v_147;
assign x_14110 = v_3171 | ~v_102;
assign x_14111 = v_3171 | ~v_101;
assign x_14112 = v_3171 | ~v_100;
assign x_14113 = ~v_130 | ~v_140 | v_3170;
assign x_14114 = ~v_122 | ~v_139 | v_3169;
assign x_14115 = ~v_115 | v_140 | v_3168;
assign x_14116 = ~v_107 | v_139 | v_3167;
assign x_14117 = v_3166 | ~v_1168;
assign x_14118 = v_3166 | ~v_1169;
assign x_14119 = v_3166 | ~v_1170;
assign x_14120 = v_3166 | ~v_1171;
assign x_14121 = v_3166 | ~v_904;
assign x_14122 = v_3166 | ~v_905;
assign x_14123 = v_3166 | ~v_3110;
assign x_14124 = v_3166 | ~v_3111;
assign x_14125 = v_3166 | ~v_784;
assign x_14126 = v_3166 | ~v_3112;
assign x_14127 = v_3166 | ~v_3113;
assign x_14128 = v_3166 | ~v_787;
assign x_14129 = v_3166 | ~v_1204;
assign x_14130 = v_3166 | ~v_1205;
assign x_14131 = v_3166 | ~v_3146;
assign x_14132 = v_3166 | ~v_3147;
assign x_14133 = v_3166 | ~v_1178;
assign x_14134 = v_3166 | ~v_3148;
assign x_14135 = v_3166 | ~v_3149;
assign x_14136 = v_3166 | ~v_1179;
assign x_14137 = v_3166 | ~v_3162;
assign x_14138 = v_3166 | ~v_3163;
assign x_14139 = v_3166 | ~v_912;
assign x_14140 = v_3166 | ~v_3164;
assign x_14141 = v_3166 | ~v_3165;
assign x_14142 = v_3166 | ~v_913;
assign x_14143 = v_3166 | ~v_3118;
assign x_14144 = v_3166 | ~v_3121;
assign x_14145 = v_3166 | ~v_916;
assign x_14146 = v_3166 | ~v_917;
assign x_14147 = v_3166 | ~v_1206;
assign x_14148 = v_3166 | ~v_1207;
assign x_14149 = v_3166 | ~v_183;
assign x_14150 = v_3166 | ~v_168;
assign x_14151 = v_3166 | ~v_167;
assign x_14152 = v_3166 | ~v_166;
assign x_14153 = v_3166 | ~v_165;
assign x_14154 = v_3166 | ~v_145;
assign x_14155 = v_3166 | ~v_144;
assign x_14156 = v_3166 | ~v_143;
assign x_14157 = v_3166 | ~v_142;
assign x_14158 = v_3166 | ~v_60;
assign x_14159 = v_3166 | ~v_59;
assign x_14160 = v_3166 | ~v_58;
assign x_14161 = ~v_88 | ~v_140 | v_3165;
assign x_14162 = ~v_80 | ~v_139 | v_3164;
assign x_14163 = ~v_73 | v_140 | v_3163;
assign x_14164 = ~v_65 | v_139 | v_3162;
assign x_14165 = v_3161 | ~v_1153;
assign x_14166 = v_3161 | ~v_1154;
assign x_14167 = v_3161 | ~v_1155;
assign x_14168 = v_3161 | ~v_1156;
assign x_14169 = v_3161 | ~v_889;
assign x_14170 = v_3161 | ~v_890;
assign x_14171 = v_3161 | ~v_3095;
assign x_14172 = v_3161 | ~v_3096;
assign x_14173 = v_3161 | ~v_751;
assign x_14174 = v_3161 | ~v_3097;
assign x_14175 = v_3161 | ~v_3098;
assign x_14176 = v_3161 | ~v_754;
assign x_14177 = v_3161 | ~v_1199;
assign x_14178 = v_3161 | ~v_1200;
assign x_14179 = v_3161 | ~v_3141;
assign x_14180 = v_3161 | ~v_3142;
assign x_14181 = v_3161 | ~v_1163;
assign x_14182 = v_3161 | ~v_3143;
assign x_14183 = v_3161 | ~v_3144;
assign x_14184 = v_3161 | ~v_1164;
assign x_14185 = v_3161 | ~v_3157;
assign x_14186 = v_3161 | ~v_3158;
assign x_14187 = v_3161 | ~v_897;
assign x_14188 = v_3161 | ~v_3159;
assign x_14189 = v_3161 | ~v_3160;
assign x_14190 = v_3161 | ~v_898;
assign x_14191 = v_3161 | ~v_901;
assign x_14192 = v_3161 | ~v_902;
assign x_14193 = v_3161 | ~v_1201;
assign x_14194 = v_3161 | ~v_1202;
assign x_14195 = v_3161 | ~v_182;
assign x_14196 = v_3161 | ~v_164;
assign x_14197 = v_3161 | ~v_163;
assign x_14198 = v_3161 | ~v_162;
assign x_14199 = v_3161 | ~v_161;
assign x_14200 = v_3161 | ~v_137;
assign x_14201 = v_3161 | ~v_136;
assign x_14202 = v_3161 | ~v_135;
assign x_14203 = v_3161 | ~v_134;
assign x_14204 = v_3161 | ~v_3107;
assign x_14205 = v_3161 | ~v_3108;
assign x_14206 = v_3161 | ~v_17;
assign x_14207 = v_3161 | ~v_16;
assign x_14208 = v_3161 | ~v_15;
assign x_14209 = ~v_46 | ~v_140 | v_3160;
assign x_14210 = ~v_38 | ~v_139 | v_3159;
assign x_14211 = ~v_31 | v_140 | v_3158;
assign x_14212 = ~v_23 | v_139 | v_3157;
assign x_14213 = ~v_3155 | ~v_3150 | ~v_3145 | v_3156;
assign x_14214 = v_3155 | ~v_1183;
assign x_14215 = v_3155 | ~v_1184;
assign x_14216 = v_3155 | ~v_1185;
assign x_14217 = v_3155 | ~v_1186;
assign x_14218 = v_3155 | ~v_965;
assign x_14219 = v_3155 | ~v_966;
assign x_14220 = v_3155 | ~v_967;
assign x_14221 = v_3155 | ~v_968;
assign x_14222 = v_3155 | ~v_3125;
assign x_14223 = v_3155 | ~v_3126;
assign x_14224 = v_3155 | ~v_817;
assign x_14225 = v_3155 | ~v_3127;
assign x_14226 = v_3155 | ~v_3128;
assign x_14227 = v_3155 | ~v_820;
assign x_14228 = v_3155 | ~v_1225;
assign x_14229 = v_3155 | ~v_1226;
assign x_14230 = v_3155 | ~v_1227;
assign x_14231 = v_3155 | ~v_1228;
assign x_14232 = v_3155 | ~v_3151;
assign x_14233 = v_3155 | ~v_3152;
assign x_14234 = v_3155 | ~v_1193;
assign x_14235 = v_3155 | ~v_3153;
assign x_14236 = v_3155 | ~v_3154;
assign x_14237 = v_3155 | ~v_1194;
assign x_14238 = v_3155 | ~v_3129;
assign x_14239 = v_3155 | ~v_3130;
assign x_14240 = v_3155 | ~v_975;
assign x_14241 = v_3155 | ~v_3131;
assign x_14242 = v_3155 | ~v_3132;
assign x_14243 = v_3155 | ~v_976;
assign x_14244 = v_3155 | ~v_3133;
assign x_14245 = v_3155 | ~v_3136;
assign x_14246 = v_3155 | ~v_184;
assign x_14247 = v_3155 | ~v_171;
assign x_14248 = v_3155 | ~v_170;
assign x_14249 = v_3155 | ~v_169;
assign x_14250 = v_3155 | ~v_150;
assign x_14251 = v_3155 | ~v_149;
assign x_14252 = v_3155 | ~v_148;
assign x_14253 = v_3155 | ~v_103;
assign x_14254 = v_3155 | ~v_102;
assign x_14255 = v_3155 | ~v_101;
assign x_14256 = v_3155 | ~v_100;
assign x_14257 = v_3155 | ~v_95;
assign x_14258 = ~v_127 | ~v_153 | v_3154;
assign x_14259 = ~v_121 | ~v_152 | v_3153;
assign x_14260 = ~v_112 | v_153 | v_3152;
assign x_14261 = ~v_106 | v_152 | v_3151;
assign x_14262 = v_3150 | ~v_1168;
assign x_14263 = v_3150 | ~v_1169;
assign x_14264 = v_3150 | ~v_1170;
assign x_14265 = v_3150 | ~v_1171;
assign x_14266 = v_3150 | ~v_950;
assign x_14267 = v_3150 | ~v_951;
assign x_14268 = v_3150 | ~v_952;
assign x_14269 = v_3150 | ~v_953;
assign x_14270 = v_3150 | ~v_3110;
assign x_14271 = v_3150 | ~v_3111;
assign x_14272 = v_3150 | ~v_784;
assign x_14273 = v_3150 | ~v_3112;
assign x_14274 = v_3150 | ~v_3113;
assign x_14275 = v_3150 | ~v_787;
assign x_14276 = v_3150 | ~v_1220;
assign x_14277 = v_3150 | ~v_1221;
assign x_14278 = v_3150 | ~v_1222;
assign x_14279 = v_3150 | ~v_1223;
assign x_14280 = v_3150 | ~v_3146;
assign x_14281 = v_3150 | ~v_3147;
assign x_14282 = v_3150 | ~v_1178;
assign x_14283 = v_3150 | ~v_3148;
assign x_14284 = v_3150 | ~v_3149;
assign x_14285 = v_3150 | ~v_1179;
assign x_14286 = v_3150 | ~v_3114;
assign x_14287 = v_3150 | ~v_3115;
assign x_14288 = v_3150 | ~v_960;
assign x_14289 = v_3150 | ~v_3116;
assign x_14290 = v_3150 | ~v_3117;
assign x_14291 = v_3150 | ~v_961;
assign x_14292 = v_3150 | ~v_3118;
assign x_14293 = v_3150 | ~v_3121;
assign x_14294 = v_3150 | ~v_183;
assign x_14295 = v_3150 | ~v_167;
assign x_14296 = v_3150 | ~v_166;
assign x_14297 = v_3150 | ~v_165;
assign x_14298 = v_3150 | ~v_145;
assign x_14299 = v_3150 | ~v_144;
assign x_14300 = v_3150 | ~v_143;
assign x_14301 = v_3150 | ~v_61;
assign x_14302 = v_3150 | ~v_60;
assign x_14303 = v_3150 | ~v_59;
assign x_14304 = v_3150 | ~v_58;
assign x_14305 = v_3150 | ~v_53;
assign x_14306 = ~v_85 | ~v_153 | v_3149;
assign x_14307 = ~v_79 | ~v_152 | v_3148;
assign x_14308 = ~v_70 | v_153 | v_3147;
assign x_14309 = ~v_64 | v_152 | v_3146;
assign x_14310 = v_3145 | ~v_1153;
assign x_14311 = v_3145 | ~v_1154;
assign x_14312 = v_3145 | ~v_1155;
assign x_14313 = v_3145 | ~v_1156;
assign x_14314 = v_3145 | ~v_935;
assign x_14315 = v_3145 | ~v_936;
assign x_14316 = v_3145 | ~v_937;
assign x_14317 = v_3145 | ~v_938;
assign x_14318 = v_3145 | ~v_3095;
assign x_14319 = v_3145 | ~v_3096;
assign x_14320 = v_3145 | ~v_751;
assign x_14321 = v_3145 | ~v_3097;
assign x_14322 = v_3145 | ~v_3098;
assign x_14323 = v_3145 | ~v_754;
assign x_14324 = v_3145 | ~v_1215;
assign x_14325 = v_3145 | ~v_1216;
assign x_14326 = v_3145 | ~v_1217;
assign x_14327 = v_3145 | ~v_1218;
assign x_14328 = v_3145 | ~v_3141;
assign x_14329 = v_3145 | ~v_3142;
assign x_14330 = v_3145 | ~v_1163;
assign x_14331 = v_3145 | ~v_3143;
assign x_14332 = v_3145 | ~v_3144;
assign x_14333 = v_3145 | ~v_1164;
assign x_14334 = v_3145 | ~v_3099;
assign x_14335 = v_3145 | ~v_3100;
assign x_14336 = v_3145 | ~v_945;
assign x_14337 = v_3145 | ~v_3101;
assign x_14338 = v_3145 | ~v_3102;
assign x_14339 = v_3145 | ~v_946;
assign x_14340 = v_3145 | ~v_182;
assign x_14341 = v_3145 | ~v_163;
assign x_14342 = v_3145 | ~v_162;
assign x_14343 = v_3145 | ~v_161;
assign x_14344 = v_3145 | ~v_137;
assign x_14345 = v_3145 | ~v_136;
assign x_14346 = v_3145 | ~v_135;
assign x_14347 = v_3145 | ~v_3107;
assign x_14348 = v_3145 | ~v_3108;
assign x_14349 = v_3145 | ~v_18;
assign x_14350 = v_3145 | ~v_17;
assign x_14351 = v_3145 | ~v_16;
assign x_14352 = v_3145 | ~v_15;
assign x_14353 = v_3145 | ~v_10;
assign x_14354 = ~v_43 | ~v_153 | v_3144;
assign x_14355 = ~v_37 | ~v_152 | v_3143;
assign x_14356 = ~v_28 | v_153 | v_3142;
assign x_14357 = ~v_22 | v_152 | v_3141;
assign x_14358 = ~v_3139 | ~v_3124 | ~v_3109 | v_3140;
assign x_14359 = v_3139 | ~v_965;
assign x_14360 = v_3139 | ~v_966;
assign x_14361 = v_3139 | ~v_967;
assign x_14362 = v_3139 | ~v_968;
assign x_14363 = v_3139 | ~v_3125;
assign x_14364 = v_3139 | ~v_3126;
assign x_14365 = v_3139 | ~v_817;
assign x_14366 = v_3139 | ~v_818;
assign x_14367 = v_3139 | ~v_819;
assign x_14368 = v_3139 | ~v_3127;
assign x_14369 = v_3139 | ~v_3128;
assign x_14370 = v_3139 | ~v_820;
assign x_14371 = v_3139 | ~v_821;
assign x_14372 = v_3139 | ~v_822;
assign x_14373 = v_3139 | ~v_1147;
assign x_14374 = v_3139 | ~v_1148;
assign x_14375 = v_3139 | ~v_3129;
assign x_14376 = v_3139 | ~v_3130;
assign x_14377 = v_3139 | ~v_975;
assign x_14378 = v_3139 | ~v_3131;
assign x_14379 = v_3139 | ~v_3132;
assign x_14380 = v_3139 | ~v_976;
assign x_14381 = v_3139 | ~v_3133;
assign x_14382 = v_3139 | ~v_3134;
assign x_14383 = v_3139 | ~v_3135;
assign x_14384 = v_3139 | ~v_839;
assign x_14385 = v_3139 | ~v_3136;
assign x_14386 = v_3139 | ~v_3137;
assign x_14387 = v_3139 | ~v_3138;
assign x_14388 = v_3139 | ~v_840;
assign x_14389 = v_3139 | ~v_1149;
assign x_14390 = v_3139 | ~v_1150;
assign x_14391 = v_3139 | ~v_184;
assign x_14392 = v_3139 | ~v_170;
assign x_14393 = v_3139 | ~v_150;
assign x_14394 = v_3139 | ~v_149;
assign x_14395 = v_3139 | ~v_148;
assign x_14396 = v_3139 | ~v_147;
assign x_14397 = v_3139 | ~v_103;
assign x_14398 = v_3139 | ~v_102;
assign x_14399 = v_3139 | ~v_101;
assign x_14400 = v_3139 | ~v_100;
assign x_14401 = v_3139 | ~v_98;
assign x_14402 = v_3139 | ~v_93;
assign x_14403 = ~v_19 | ~v_127 | v_3138;
assign x_14404 = ~v_19 | ~v_121 | v_3137;
assign x_14405 = ~v_19 | ~v_119 | v_3136;
assign x_14406 = v_19 | ~v_112 | v_3135;
assign x_14407 = v_19 | ~v_106 | v_3134;
assign x_14408 = v_19 | ~v_104 | v_3133;
assign x_14409 = ~v_130 | ~v_153 | v_3132;
assign x_14410 = ~v_122 | ~v_152 | v_3131;
assign x_14411 = ~v_115 | v_153 | v_3130;
assign x_14412 = ~v_107 | v_152 | v_3129;
assign x_14413 = ~v_123 | ~v_157 | v_3128;
assign x_14414 = ~v_120 | ~v_156 | v_3127;
assign x_14415 = ~v_108 | v_157 | v_3126;
assign x_14416 = ~v_105 | v_156 | v_3125;
assign x_14417 = v_3124 | ~v_950;
assign x_14418 = v_3124 | ~v_951;
assign x_14419 = v_3124 | ~v_952;
assign x_14420 = v_3124 | ~v_953;
assign x_14421 = v_3124 | ~v_3110;
assign x_14422 = v_3124 | ~v_3111;
assign x_14423 = v_3124 | ~v_784;
assign x_14424 = v_3124 | ~v_785;
assign x_14425 = v_3124 | ~v_786;
assign x_14426 = v_3124 | ~v_3112;
assign x_14427 = v_3124 | ~v_3113;
assign x_14428 = v_3124 | ~v_787;
assign x_14429 = v_3124 | ~v_788;
assign x_14430 = v_3124 | ~v_789;
assign x_14431 = v_3124 | ~v_1142;
assign x_14432 = v_3124 | ~v_1143;
assign x_14433 = v_3124 | ~v_3114;
assign x_14434 = v_3124 | ~v_3115;
assign x_14435 = v_3124 | ~v_960;
assign x_14436 = v_3124 | ~v_3116;
assign x_14437 = v_3124 | ~v_3117;
assign x_14438 = v_3124 | ~v_961;
assign x_14439 = v_3124 | ~v_3118;
assign x_14440 = v_3124 | ~v_3119;
assign x_14441 = v_3124 | ~v_3120;
assign x_14442 = v_3124 | ~v_806;
assign x_14443 = v_3124 | ~v_3121;
assign x_14444 = v_3124 | ~v_3122;
assign x_14445 = v_3124 | ~v_3123;
assign x_14446 = v_3124 | ~v_807;
assign x_14447 = v_3124 | ~v_1144;
assign x_14448 = v_3124 | ~v_1145;
assign x_14449 = v_3124 | ~v_183;
assign x_14450 = v_3124 | ~v_166;
assign x_14451 = v_3124 | ~v_145;
assign x_14452 = v_3124 | ~v_144;
assign x_14453 = v_3124 | ~v_143;
assign x_14454 = v_3124 | ~v_142;
assign x_14455 = v_3124 | ~v_61;
assign x_14456 = v_3124 | ~v_60;
assign x_14457 = v_3124 | ~v_59;
assign x_14458 = v_3124 | ~v_58;
assign x_14459 = v_3124 | ~v_56;
assign x_14460 = v_3124 | ~v_51;
assign x_14461 = ~v_19 | ~v_85 | v_3123;
assign x_14462 = ~v_19 | ~v_79 | v_3122;
assign x_14463 = ~v_19 | ~v_77 | v_3121;
assign x_14464 = v_19 | ~v_70 | v_3120;
assign x_14465 = v_19 | ~v_64 | v_3119;
assign x_14466 = v_19 | ~v_62 | v_3118;
assign x_14467 = ~v_88 | ~v_153 | v_3117;
assign x_14468 = ~v_80 | ~v_152 | v_3116;
assign x_14469 = ~v_73 | v_153 | v_3115;
assign x_14470 = ~v_65 | v_152 | v_3114;
assign x_14471 = ~v_81 | ~v_157 | v_3113;
assign x_14472 = ~v_78 | ~v_156 | v_3112;
assign x_14473 = ~v_66 | v_157 | v_3111;
assign x_14474 = ~v_63 | v_156 | v_3110;
assign x_14475 = v_3109 | ~v_935;
assign x_14476 = v_3109 | ~v_936;
assign x_14477 = v_3109 | ~v_937;
assign x_14478 = v_3109 | ~v_938;
assign x_14479 = v_3109 | ~v_3095;
assign x_14480 = v_3109 | ~v_3096;
assign x_14481 = v_3109 | ~v_751;
assign x_14482 = v_3109 | ~v_752;
assign x_14483 = v_3109 | ~v_753;
assign x_14484 = v_3109 | ~v_3097;
assign x_14485 = v_3109 | ~v_3098;
assign x_14486 = v_3109 | ~v_754;
assign x_14487 = v_3109 | ~v_755;
assign x_14488 = v_3109 | ~v_756;
assign x_14489 = v_3109 | ~v_1137;
assign x_14490 = v_3109 | ~v_1138;
assign x_14491 = v_3109 | ~v_3099;
assign x_14492 = v_3109 | ~v_3100;
assign x_14493 = v_3109 | ~v_945;
assign x_14494 = v_3109 | ~v_3101;
assign x_14495 = v_3109 | ~v_3102;
assign x_14496 = v_3109 | ~v_946;
assign x_14497 = v_3109 | ~v_3103;
assign x_14498 = v_3109 | ~v_3104;
assign x_14499 = v_3109 | ~v_773;
assign x_14500 = v_3109 | ~v_3105;
assign x_14501 = v_3109 | ~v_3106;
assign x_14502 = v_3109 | ~v_774;
assign x_14503 = v_3109 | ~v_1139;
assign x_14504 = v_3109 | ~v_1140;
assign x_14505 = v_3109 | ~v_182;
assign x_14506 = v_3109 | ~v_162;
assign x_14507 = v_3109 | ~v_137;
assign x_14508 = v_3109 | ~v_136;
assign x_14509 = v_3109 | ~v_135;
assign x_14510 = v_3109 | ~v_134;
assign x_14511 = v_3109 | ~v_3107;
assign x_14512 = v_3109 | ~v_3108;
assign x_14513 = v_3109 | ~v_18;
assign x_14514 = v_3109 | ~v_17;
assign x_14515 = v_3109 | ~v_16;
assign x_14516 = v_3109 | ~v_15;
assign x_14517 = v_3109 | ~v_13;
assign x_14518 = v_3109 | ~v_8;
assign x_14519 = ~v_19 | ~v_35 | v_3108;
assign x_14520 = ~v_20 | v_19 | v_3107;
assign x_14521 = ~v_19 | ~v_43 | v_3106;
assign x_14522 = ~v_19 | ~v_37 | v_3105;
assign x_14523 = ~v_28 | v_19 | v_3104;
assign x_14524 = ~v_22 | v_19 | v_3103;
assign x_14525 = ~v_46 | ~v_153 | v_3102;
assign x_14526 = ~v_38 | ~v_152 | v_3101;
assign x_14527 = ~v_31 | v_153 | v_3100;
assign x_14528 = ~v_23 | v_152 | v_3099;
assign x_14529 = ~v_39 | ~v_157 | v_3098;
assign x_14530 = ~v_36 | ~v_156 | v_3097;
assign x_14531 = ~v_24 | v_157 | v_3096;
assign x_14532 = ~v_21 | v_156 | v_3095;
assign x_14533 = v_3094 | ~v_733;
assign x_14534 = v_3094 | ~v_728;
assign x_14535 = v_3093 | ~v_2034;
assign x_14536 = v_3093 | ~v_737;
assign x_14537 = ~v_725 | ~v_724 | ~v_723 | ~v_722 | ~v_3091 | ~v_3087 | ~v_3083 | ~v_3079 | ~v_3075 | ~v_3059 | ~v_3055 | ~v_3051 | ~v_3047 | ~v_3043 | ~v_3027 | ~v_3023 | ~v_3007 | ~v_2991 | ~v_2975 | ~v_2959 | ~v_2913 | v_3092;
assign x_14538 = v_3091 | ~v_3088;
assign x_14539 = v_3091 | ~v_3089;
assign x_14540 = v_3091 | ~v_3090;
assign x_14541 = v_98 | v_103 | v_101 | v_96 | v_100 | v_95 | v_99 | v_93 | v_102 | ~v_719 | ~v_718 | v_170 | v_149 | v_184 | ~v_483 | ~v_717 | ~v_3021 | ~v_299 | ~v_2957 | ~v_3020 | ~v_2956 | ~v_2955 | ~v_482 | ~v_716 | ~v_3019 | ~v_298 | ~v_2954 | ~v_3018 | ~v_2953 | ~v_2952 | ~v_473 | ~v_281 | ~v_472 | ~v_280 | ~v_279 | ~v_2947 | ~v_2946 | ~v_471 | ~v_278 | ~v_470 | ~v_277 | ~v_276 | ~v_2945 | ~v_2944 | v_3090;
assign x_14542 = v_54 | v_53 | v_56 | v_61 | v_51 | v_60 | v_59 | v_58 | v_57 | ~v_714 | ~v_713 | ~v_3016 | v_144 | v_166 | v_183 | ~v_3015 | ~v_266 | ~v_2942 | ~v_468 | ~v_712 | ~v_2941 | ~v_2940 | ~v_467 | ~v_711 | ~v_3014 | ~v_265 | ~v_2939 | ~v_3013 | ~v_2938 | ~v_2937 | ~v_458 | ~v_248 | ~v_457 | ~v_247 | ~v_246 | ~v_2932 | ~v_2931 | ~v_456 | ~v_245 | ~v_455 | ~v_244 | ~v_243 | ~v_2930 | ~v_2929 | v_3089;
assign x_14543 = v_13 | v_18 | v_17 | v_16 | v_8 | v_15 | v_14 | v_11 | v_10 | ~v_453 | ~v_709 | ~v_2927 | ~v_452 | ~v_708 | ~v_2926 | v_136 | ~v_707 | ~v_706 | v_162 | v_182 | ~v_3011 | ~v_233 | ~v_2925 | ~v_3010 | ~v_2924 | ~v_3009 | ~v_232 | ~v_2923 | ~v_3008 | ~v_2922 | ~v_443 | ~v_215 | ~v_442 | ~v_214 | ~v_213 | ~v_2917 | ~v_2916 | ~v_441 | ~v_212 | ~v_440 | ~v_211 | ~v_210 | ~v_2915 | ~v_2914 | v_3088;
assign x_14544 = v_3087 | ~v_3084;
assign x_14545 = v_3087 | ~v_3085;
assign x_14546 = v_3087 | ~v_3086;
assign x_14547 = v_103 | v_101 | v_96 | v_94 | v_99 | v_102 | v_171 | v_169 | v_149 | v_147 | v_184 | v_181 | ~v_483 | ~v_3021 | ~v_3020 | ~v_2955 | ~v_482 | ~v_3019 | ~v_3018 | ~v_2952 | ~v_481 | ~v_480 | ~v_345 | ~v_3073 | ~v_3072 | ~v_479 | ~v_478 | ~v_344 | ~v_3071 | ~v_3070 | ~v_473 | ~v_472 | ~v_279 | ~v_2947 | ~v_2946 | ~v_471 | ~v_470 | ~v_276 | ~v_2945 | ~v_2944 | ~v_335 | ~v_334 | ~v_333 | ~v_332 | v_3086;
assign x_14548 = v_54 | v_61 | v_52 | v_60 | v_59 | v_57 | ~v_3016 | v_144 | v_180 | v_142 | v_167 | v_165 | v_183 | ~v_3015 | ~v_468 | ~v_2940 | ~v_467 | ~v_3014 | ~v_3013 | ~v_2937 | ~v_466 | ~v_465 | ~v_330 | ~v_3068 | ~v_3067 | ~v_464 | ~v_463 | ~v_329 | ~v_3066 | ~v_3065 | ~v_458 | ~v_457 | ~v_246 | ~v_2932 | ~v_2931 | ~v_456 | ~v_455 | ~v_243 | ~v_2930 | ~v_2929 | ~v_320 | ~v_319 | ~v_318 | ~v_317 | v_3085;
assign x_14549 = v_9 | v_18 | v_17 | v_16 | v_14 | v_11 | ~v_453 | ~v_2927 | ~v_452 | ~v_2926 | v_136 | v_134 | v_179 | v_163 | v_161 | v_182 | ~v_3011 | ~v_3010 | ~v_3009 | ~v_3008 | ~v_451 | ~v_450 | ~v_315 | ~v_3063 | ~v_3062 | ~v_449 | ~v_448 | ~v_314 | ~v_3061 | ~v_3060 | ~v_443 | ~v_442 | ~v_213 | ~v_2917 | ~v_2916 | ~v_441 | ~v_440 | ~v_210 | ~v_2915 | ~v_2914 | ~v_305 | ~v_304 | ~v_303 | ~v_302 | v_3084;
assign x_14550 = v_3083 | ~v_3080;
assign x_14551 = v_3083 | ~v_3081;
assign x_14552 = v_3083 | ~v_3082;
assign x_14553 = v_103 | v_97 | v_95 | v_94 | v_102 | v_171 | v_169 | v_160 | v_150 | v_148 | v_184 | v_181 | ~v_2955 | ~v_2952 | ~v_297 | ~v_3005 | ~v_3004 | ~v_296 | ~v_3003 | ~v_3002 | ~v_345 | ~v_3073 | ~v_3072 | ~v_344 | ~v_3071 | ~v_3070 | ~v_343 | ~v_342 | ~v_341 | ~v_340 | ~v_279 | ~v_2947 | ~v_2946 | ~v_276 | ~v_2945 | ~v_2944 | ~v_335 | ~v_334 | ~v_333 | ~v_332 | ~v_275 | ~v_274 | ~v_273 | ~v_272 | v_3082;
assign x_14554 = v_53 | v_55 | v_61 | v_52 | v_60 | v_180 | v_159 | v_145 | v_143 | v_167 | v_165 | v_183 | ~v_2940 | ~v_2937 | ~v_264 | ~v_3000 | ~v_2999 | ~v_263 | ~v_2998 | ~v_2997 | ~v_330 | ~v_3068 | ~v_3067 | ~v_329 | ~v_3066 | ~v_3065 | ~v_328 | ~v_327 | ~v_326 | ~v_325 | ~v_246 | ~v_2932 | ~v_2931 | ~v_243 | ~v_2930 | ~v_2929 | ~v_320 | ~v_319 | ~v_318 | ~v_317 | ~v_242 | ~v_241 | ~v_240 | ~v_239 | v_3081;
assign x_14555 = v_9 | v_18 | v_17 | v_12 | v_10 | ~v_2927 | ~v_2926 | v_135 | v_137 | v_179 | v_163 | v_161 | v_155 | v_182 | ~v_231 | ~v_2995 | ~v_2994 | ~v_230 | ~v_2993 | ~v_2992 | ~v_315 | ~v_3063 | ~v_3062 | ~v_314 | ~v_3061 | ~v_3060 | ~v_313 | ~v_312 | ~v_311 | ~v_310 | ~v_213 | ~v_2917 | ~v_2916 | ~v_210 | ~v_2915 | ~v_2914 | ~v_305 | ~v_304 | ~v_303 | ~v_302 | ~v_209 | ~v_208 | ~v_207 | ~v_206 | v_3080;
assign x_14556 = v_3079 | ~v_3076;
assign x_14557 = v_3079 | ~v_3077;
assign x_14558 = v_3079 | ~v_3078;
assign x_14559 = v_103 | v_101 | v_94 | v_102 | v_171 | v_169 | v_150 | v_149 | v_148 | v_147 | v_184 | v_181 | ~v_391 | ~v_390 | ~v_389 | ~v_388 | ~v_2955 | ~v_2952 | ~v_387 | ~v_2989 | ~v_2988 | ~v_386 | ~v_2987 | ~v_2986 | ~v_345 | ~v_3073 | ~v_3072 | ~v_344 | ~v_3071 | ~v_3070 | ~v_385 | ~v_384 | ~v_279 | ~v_2947 | ~v_2946 | ~v_276 | ~v_2945 | ~v_2944 | ~v_335 | ~v_334 | ~v_333 | ~v_332 | ~v_379 | ~v_378 | v_3078;
assign x_14560 = v_61 | v_52 | v_60 | v_59 | v_144 | v_180 | v_145 | v_143 | v_142 | v_167 | v_165 | v_183 | ~v_376 | ~v_375 | ~v_374 | ~v_373 | ~v_2940 | ~v_2937 | ~v_372 | ~v_2984 | ~v_2983 | ~v_371 | ~v_2982 | ~v_2981 | ~v_330 | ~v_3068 | ~v_3067 | ~v_329 | ~v_3066 | ~v_3065 | ~v_370 | ~v_369 | ~v_246 | ~v_2932 | ~v_2931 | ~v_243 | ~v_2930 | ~v_2929 | ~v_320 | ~v_319 | ~v_318 | ~v_317 | ~v_364 | ~v_363 | v_3077;
assign x_14561 = v_9 | v_18 | v_17 | v_16 | ~v_2927 | ~v_2926 | v_136 | v_135 | v_134 | v_137 | v_179 | v_163 | v_161 | v_182 | ~v_361 | ~v_360 | ~v_359 | ~v_358 | ~v_357 | ~v_2979 | ~v_2978 | ~v_356 | ~v_2977 | ~v_2976 | ~v_315 | ~v_3063 | ~v_3062 | ~v_314 | ~v_3061 | ~v_3060 | ~v_355 | ~v_354 | ~v_213 | ~v_2917 | ~v_2916 | ~v_210 | ~v_2915 | ~v_2914 | ~v_305 | ~v_304 | ~v_303 | ~v_302 | ~v_349 | ~v_348 | v_3076;
assign x_14562 = v_3075 | ~v_3064;
assign x_14563 = v_3075 | ~v_3069;
assign x_14564 = v_3075 | ~v_3074;
assign x_14565 = v_101 | v_94 | v_102 | v_172 | v_171 | v_169 | v_150 | v_149 | v_148 | v_147 | v_184 | v_181 | ~v_437 | ~v_436 | ~v_2955 | ~v_2952 | ~v_435 | ~v_2951 | ~v_2950 | ~v_434 | ~v_2949 | ~v_2948 | ~v_345 | ~v_3073 | ~v_3072 | ~v_344 | ~v_3071 | ~v_3070 | ~v_433 | ~v_432 | ~v_279 | ~v_2947 | ~v_2946 | ~v_276 | ~v_2945 | ~v_2944 | ~v_335 | ~v_334 | ~v_333 | ~v_332 | ~v_427 | ~v_426 | ~v_425 | ~v_424 | v_3074;
assign x_14566 = v_3073 | v_157;
assign x_14567 = v_3073 | v_127;
assign x_14568 = v_3072 | v_156;
assign x_14569 = v_3072 | v_121;
assign x_14570 = v_3071 | ~v_157;
assign x_14571 = v_3071 | v_112;
assign x_14572 = v_3070 | ~v_156;
assign x_14573 = v_3070 | v_106;
assign x_14574 = v_52 | v_60 | v_59 | v_144 | v_180 | v_145 | v_143 | v_142 | v_168 | v_167 | v_165 | v_183 | ~v_422 | ~v_421 | ~v_2940 | ~v_2937 | ~v_420 | ~v_2936 | ~v_2935 | ~v_419 | ~v_2934 | ~v_2933 | ~v_330 | ~v_3068 | ~v_3067 | ~v_329 | ~v_3066 | ~v_3065 | ~v_418 | ~v_417 | ~v_246 | ~v_2932 | ~v_2931 | ~v_243 | ~v_2930 | ~v_2929 | ~v_320 | ~v_319 | ~v_318 | ~v_317 | ~v_412 | ~v_411 | ~v_410 | ~v_409 | v_3069;
assign x_14575 = v_3068 | v_157;
assign x_14576 = v_3068 | v_85;
assign x_14577 = v_3067 | v_156;
assign x_14578 = v_3067 | v_79;
assign x_14579 = v_3066 | ~v_157;
assign x_14580 = v_3066 | v_70;
assign x_14581 = v_3065 | ~v_156;
assign x_14582 = v_3065 | v_64;
assign x_14583 = v_9 | v_17 | v_16 | ~v_2927 | ~v_2926 | v_136 | v_135 | v_134 | v_137 | v_179 | v_164 | v_163 | v_161 | v_182 | ~v_407 | ~v_406 | ~v_405 | ~v_2921 | ~v_2920 | ~v_404 | ~v_2919 | ~v_2918 | ~v_315 | ~v_3063 | ~v_3062 | ~v_314 | ~v_3061 | ~v_3060 | ~v_403 | ~v_402 | ~v_213 | ~v_2917 | ~v_2916 | ~v_210 | ~v_2915 | ~v_2914 | ~v_305 | ~v_304 | ~v_303 | ~v_302 | ~v_397 | ~v_396 | ~v_395 | ~v_394 | v_3064;
assign x_14584 = v_3063 | v_157;
assign x_14585 = v_3063 | v_43;
assign x_14586 = v_3062 | v_156;
assign x_14587 = v_3062 | v_37;
assign x_14588 = v_3061 | ~v_157;
assign x_14589 = v_3061 | v_28;
assign x_14590 = v_3060 | ~v_156;
assign x_14591 = v_3060 | v_22;
assign x_14592 = v_3059 | ~v_3056;
assign x_14593 = v_3059 | ~v_3057;
assign x_14594 = v_3059 | ~v_3058;
assign x_14595 = v_98 | v_103 | v_97 | v_100 | v_93 | v_102 | v_170 | v_160 | v_150 | v_148 | v_147 | v_184 | ~v_299 | ~v_2957 | ~v_2956 | ~v_2955 | ~v_298 | ~v_2954 | ~v_2953 | ~v_2952 | ~v_297 | ~v_3005 | ~v_3004 | ~v_296 | ~v_3003 | ~v_3002 | ~v_295 | ~v_294 | ~v_293 | ~v_292 | ~v_281 | ~v_280 | ~v_279 | ~v_2947 | ~v_2946 | ~v_278 | ~v_277 | ~v_276 | ~v_2945 | ~v_2944 | ~v_275 | ~v_274 | ~v_273 | ~v_272 | v_3058;
assign x_14596 = v_56 | v_55 | v_61 | v_51 | v_60 | v_58 | v_159 | v_145 | v_143 | v_142 | v_166 | v_183 | ~v_266 | ~v_2942 | ~v_2941 | ~v_2940 | ~v_265 | ~v_2939 | ~v_2938 | ~v_2937 | ~v_264 | ~v_3000 | ~v_2999 | ~v_263 | ~v_2998 | ~v_2997 | ~v_262 | ~v_261 | ~v_260 | ~v_259 | ~v_248 | ~v_247 | ~v_246 | ~v_2932 | ~v_2931 | ~v_245 | ~v_244 | ~v_243 | ~v_2930 | ~v_2929 | ~v_242 | ~v_241 | ~v_240 | ~v_239 | v_3057;
assign x_14597 = v_13 | v_18 | v_17 | v_8 | v_15 | v_12 | ~v_2927 | ~v_2926 | v_135 | v_134 | v_137 | v_162 | v_155 | v_182 | ~v_233 | ~v_2925 | ~v_2924 | ~v_232 | ~v_2923 | ~v_2922 | ~v_231 | ~v_2995 | ~v_2994 | ~v_230 | ~v_2993 | ~v_2992 | ~v_229 | ~v_228 | ~v_227 | ~v_226 | ~v_215 | ~v_214 | ~v_213 | ~v_2917 | ~v_2916 | ~v_212 | ~v_211 | ~v_210 | ~v_2915 | ~v_2914 | ~v_209 | ~v_208 | ~v_207 | ~v_206 | v_3056;
assign x_14598 = v_3055 | ~v_3052;
assign x_14599 = v_3055 | ~v_3053;
assign x_14600 = v_3055 | ~v_3054;
assign x_14601 = v_101 | v_96 | v_100 | v_99 | v_102 | v_172 | v_171 | v_170 | v_169 | v_149 | v_147 | v_184 | ~v_483 | ~v_3021 | ~v_3020 | ~v_2955 | ~v_482 | ~v_3019 | ~v_3018 | ~v_2952 | ~v_593 | ~v_592 | ~v_545 | ~v_3041 | ~v_3040 | ~v_591 | ~v_590 | ~v_544 | ~v_3039 | ~v_3038 | ~v_473 | ~v_472 | ~v_279 | ~v_2947 | ~v_2946 | ~v_471 | ~v_470 | ~v_276 | ~v_2945 | ~v_2944 | ~v_535 | ~v_534 | ~v_533 | ~v_532 | v_3054;
assign x_14602 = v_54 | v_60 | v_59 | v_58 | v_57 | ~v_3016 | v_144 | v_142 | v_168 | v_167 | v_166 | v_165 | v_183 | ~v_3015 | ~v_468 | ~v_2940 | ~v_467 | ~v_3014 | ~v_3013 | ~v_2937 | ~v_588 | ~v_587 | ~v_530 | ~v_3036 | ~v_3035 | ~v_586 | ~v_585 | ~v_529 | ~v_3034 | ~v_3033 | ~v_458 | ~v_457 | ~v_246 | ~v_2932 | ~v_2931 | ~v_456 | ~v_455 | ~v_243 | ~v_2930 | ~v_2929 | ~v_520 | ~v_519 | ~v_518 | ~v_517 | v_3053;
assign x_14603 = v_17 | v_16 | v_15 | v_14 | v_11 | ~v_453 | ~v_2927 | ~v_452 | ~v_2926 | v_136 | v_134 | v_164 | v_163 | v_162 | v_161 | v_182 | ~v_3011 | ~v_3010 | ~v_3009 | ~v_3008 | ~v_583 | ~v_582 | ~v_515 | ~v_3031 | ~v_3030 | ~v_581 | ~v_580 | ~v_514 | ~v_3029 | ~v_3028 | ~v_443 | ~v_442 | ~v_213 | ~v_2917 | ~v_2916 | ~v_441 | ~v_440 | ~v_210 | ~v_2915 | ~v_2914 | ~v_505 | ~v_504 | ~v_503 | ~v_502 | v_3052;
assign x_14604 = v_3051 | ~v_3048;
assign x_14605 = v_3051 | ~v_3049;
assign x_14606 = v_3051 | ~v_3050;
assign x_14607 = v_103 | v_97 | v_100 | v_102 | v_171 | v_170 | v_169 | v_160 | v_150 | v_148 | v_147 | v_184 | ~v_2955 | ~v_2952 | ~v_545 | ~v_3041 | ~v_3040 | ~v_544 | ~v_3039 | ~v_3038 | ~v_543 | ~v_542 | ~v_541 | ~v_540 | ~v_297 | ~v_3005 | ~v_3004 | ~v_296 | ~v_3003 | ~v_3002 | ~v_279 | ~v_2947 | ~v_2946 | ~v_276 | ~v_2945 | ~v_2944 | ~v_275 | ~v_274 | ~v_273 | ~v_272 | ~v_535 | ~v_534 | ~v_533 | ~v_532 | v_3050;
assign x_14608 = v_55 | v_61 | v_60 | v_58 | v_159 | v_145 | v_143 | v_142 | v_167 | v_166 | v_165 | v_183 | ~v_2940 | ~v_2937 | ~v_530 | ~v_3036 | ~v_3035 | ~v_529 | ~v_3034 | ~v_3033 | ~v_528 | ~v_527 | ~v_526 | ~v_525 | ~v_264 | ~v_3000 | ~v_2999 | ~v_263 | ~v_2998 | ~v_2997 | ~v_246 | ~v_2932 | ~v_2931 | ~v_243 | ~v_2930 | ~v_2929 | ~v_242 | ~v_241 | ~v_240 | ~v_239 | ~v_520 | ~v_519 | ~v_518 | ~v_517 | v_3049;
assign x_14609 = v_18 | v_17 | v_15 | v_12 | ~v_2927 | ~v_2926 | v_135 | v_134 | v_137 | v_163 | v_162 | v_161 | v_155 | v_182 | ~v_515 | ~v_3031 | ~v_3030 | ~v_514 | ~v_3029 | ~v_3028 | ~v_513 | ~v_512 | ~v_511 | ~v_510 | ~v_231 | ~v_2995 | ~v_2994 | ~v_230 | ~v_2993 | ~v_2992 | ~v_213 | ~v_2917 | ~v_2916 | ~v_210 | ~v_2915 | ~v_2914 | ~v_209 | ~v_208 | ~v_207 | ~v_206 | ~v_505 | ~v_504 | ~v_503 | ~v_502 | v_3048;
assign x_14610 = v_3047 | ~v_3044;
assign x_14611 = v_3047 | ~v_3045;
assign x_14612 = v_3047 | ~v_3046;
assign x_14613 = v_103 | v_101 | v_100 | v_95 | v_102 | v_171 | v_170 | v_169 | v_150 | v_149 | v_148 | v_184 | ~v_389 | ~v_388 | ~v_2955 | ~v_2952 | ~v_545 | ~v_3041 | ~v_3040 | ~v_544 | ~v_3039 | ~v_3038 | ~v_561 | ~v_560 | ~v_559 | ~v_558 | ~v_387 | ~v_2989 | ~v_2988 | ~v_386 | ~v_2987 | ~v_2986 | ~v_279 | ~v_2947 | ~v_2946 | ~v_276 | ~v_2945 | ~v_2944 | ~v_379 | ~v_378 | ~v_535 | ~v_534 | ~v_533 | ~v_532 | v_3046;
assign x_14614 = v_53 | v_61 | v_60 | v_59 | v_58 | v_144 | v_145 | v_143 | v_167 | v_166 | v_165 | v_183 | ~v_374 | ~v_373 | ~v_2940 | ~v_2937 | ~v_530 | ~v_3036 | ~v_3035 | ~v_529 | ~v_3034 | ~v_3033 | ~v_556 | ~v_555 | ~v_554 | ~v_553 | ~v_372 | ~v_2984 | ~v_2983 | ~v_371 | ~v_2982 | ~v_2981 | ~v_246 | ~v_2932 | ~v_2931 | ~v_243 | ~v_2930 | ~v_2929 | ~v_364 | ~v_363 | ~v_520 | ~v_519 | ~v_518 | ~v_517 | v_3045;
assign x_14615 = v_18 | v_17 | v_16 | v_15 | v_10 | ~v_2927 | ~v_2926 | v_136 | v_135 | v_137 | v_163 | v_162 | v_161 | v_182 | ~v_359 | ~v_358 | ~v_515 | ~v_3031 | ~v_3030 | ~v_514 | ~v_3029 | ~v_3028 | ~v_551 | ~v_550 | ~v_549 | ~v_548 | ~v_357 | ~v_2979 | ~v_2978 | ~v_356 | ~v_2977 | ~v_2976 | ~v_213 | ~v_2917 | ~v_2916 | ~v_210 | ~v_2915 | ~v_2914 | ~v_349 | ~v_348 | ~v_505 | ~v_504 | ~v_503 | ~v_502 | v_3044;
assign x_14616 = v_3043 | ~v_3032;
assign x_14617 = v_3043 | ~v_3037;
assign x_14618 = v_3043 | ~v_3042;
assign x_14619 = v_103 | v_101 | v_100 | v_151 | v_171 | v_170 | v_169 | v_150 | v_149 | v_148 | v_147 | v_184 | ~v_577 | ~v_576 | ~v_2955 | ~v_2952 | ~v_545 | ~v_3041 | ~v_3040 | ~v_544 | ~v_3039 | ~v_3038 | ~v_575 | ~v_574 | ~v_435 | ~v_2951 | ~v_2950 | ~v_434 | ~v_2949 | ~v_2948 | ~v_279 | ~v_2947 | ~v_2946 | ~v_276 | ~v_2945 | ~v_2944 | ~v_427 | ~v_426 | ~v_425 | ~v_424 | ~v_535 | ~v_534 | ~v_533 | ~v_532 | v_3042;
assign x_14620 = v_3041 | v_140;
assign x_14621 = v_3041 | v_127;
assign x_14622 = v_3040 | v_139;
assign x_14623 = v_3040 | v_121;
assign x_14624 = v_3039 | ~v_140;
assign x_14625 = v_3039 | v_112;
assign x_14626 = v_3038 | ~v_139;
assign x_14627 = v_3038 | v_106;
assign x_14628 = v_61 | v_59 | v_58 | v_144 | v_145 | v_143 | v_142 | v_167 | v_166 | v_165 | v_146 | v_183 | ~v_572 | ~v_571 | ~v_2940 | ~v_2937 | ~v_530 | ~v_3036 | ~v_3035 | ~v_529 | ~v_3034 | ~v_3033 | ~v_570 | ~v_569 | ~v_420 | ~v_2936 | ~v_2935 | ~v_419 | ~v_2934 | ~v_2933 | ~v_246 | ~v_2932 | ~v_2931 | ~v_243 | ~v_2930 | ~v_2929 | ~v_412 | ~v_411 | ~v_410 | ~v_409 | ~v_520 | ~v_519 | ~v_518 | ~v_517 | v_3037;
assign x_14629 = v_3036 | v_140;
assign x_14630 = v_3036 | v_85;
assign x_14631 = v_3035 | v_139;
assign x_14632 = v_3035 | v_79;
assign x_14633 = v_3034 | ~v_140;
assign x_14634 = v_3034 | v_70;
assign x_14635 = v_3033 | ~v_139;
assign x_14636 = v_3033 | v_64;
assign x_14637 = v_18 | v_16 | v_15 | ~v_2927 | ~v_2926 | v_136 | v_135 | v_134 | v_137 | v_138 | v_163 | v_162 | v_161 | v_182 | ~v_567 | ~v_566 | ~v_515 | ~v_3031 | ~v_3030 | ~v_514 | ~v_3029 | ~v_3028 | ~v_565 | ~v_564 | ~v_405 | ~v_2921 | ~v_2920 | ~v_404 | ~v_2919 | ~v_2918 | ~v_213 | ~v_2917 | ~v_2916 | ~v_210 | ~v_2915 | ~v_2914 | ~v_397 | ~v_396 | ~v_395 | ~v_394 | ~v_505 | ~v_504 | ~v_503 | ~v_502 | v_3032;
assign x_14638 = v_3031 | v_140;
assign x_14639 = v_3031 | v_43;
assign x_14640 = v_3030 | v_139;
assign x_14641 = v_3030 | v_37;
assign x_14642 = v_3029 | ~v_140;
assign x_14643 = v_3029 | v_28;
assign x_14644 = v_3028 | ~v_139;
assign x_14645 = v_3028 | v_22;
assign x_14646 = v_3027 | ~v_3024;
assign x_14647 = v_3027 | ~v_3025;
assign x_14648 = v_3027 | ~v_3026;
assign x_14649 = v_98 | v_103 | v_101 | v_100 | v_93 | v_151 | v_170 | v_150 | v_149 | v_148 | v_147 | v_184 | ~v_389 | ~v_388 | ~v_299 | ~v_2957 | ~v_2956 | ~v_2955 | ~v_298 | ~v_2954 | ~v_2953 | ~v_2952 | ~v_387 | ~v_2989 | ~v_2988 | ~v_386 | ~v_2987 | ~v_2986 | ~v_499 | ~v_498 | ~v_497 | ~v_496 | ~v_281 | ~v_280 | ~v_279 | ~v_2947 | ~v_2946 | ~v_278 | ~v_277 | ~v_276 | ~v_2945 | ~v_2944 | ~v_379 | ~v_378 | v_3026;
assign x_14650 = v_56 | v_61 | v_51 | v_59 | v_58 | v_144 | v_145 | v_143 | v_142 | v_166 | v_146 | v_183 | ~v_374 | ~v_373 | ~v_266 | ~v_2942 | ~v_2941 | ~v_2940 | ~v_265 | ~v_2939 | ~v_2938 | ~v_2937 | ~v_372 | ~v_2984 | ~v_2983 | ~v_371 | ~v_2982 | ~v_2981 | ~v_494 | ~v_493 | ~v_492 | ~v_491 | ~v_248 | ~v_247 | ~v_246 | ~v_2932 | ~v_2931 | ~v_245 | ~v_244 | ~v_243 | ~v_2930 | ~v_2929 | ~v_364 | ~v_363 | v_3025;
assign x_14651 = v_13 | v_18 | v_16 | v_8 | v_15 | ~v_2927 | ~v_2926 | v_136 | v_135 | v_134 | v_137 | v_138 | v_162 | v_182 | ~v_359 | ~v_358 | ~v_233 | ~v_2925 | ~v_2924 | ~v_232 | ~v_2923 | ~v_2922 | ~v_357 | ~v_2979 | ~v_2978 | ~v_356 | ~v_2977 | ~v_2976 | ~v_489 | ~v_488 | ~v_487 | ~v_486 | ~v_215 | ~v_214 | ~v_213 | ~v_2917 | ~v_2916 | ~v_212 | ~v_211 | ~v_210 | ~v_2915 | ~v_2914 | ~v_349 | ~v_348 | v_3024;
assign x_14652 = v_3023 | ~v_3012;
assign x_14653 = v_3023 | ~v_3017;
assign x_14654 = v_3023 | ~v_3022;
assign x_14655 = v_103 | v_101 | v_96 | v_100 | v_99 | v_102 | v_171 | v_170 | v_169 | v_149 | v_147 | v_184 | ~v_703 | ~v_702 | ~v_483 | ~v_3021 | ~v_3020 | ~v_2955 | ~v_482 | ~v_3019 | ~v_3018 | ~v_2952 | ~v_701 | ~v_653 | ~v_2973 | ~v_2972 | ~v_700 | ~v_652 | ~v_2971 | ~v_2970 | ~v_473 | ~v_472 | ~v_279 | ~v_2947 | ~v_2946 | ~v_471 | ~v_470 | ~v_276 | ~v_2945 | ~v_2944 | ~v_645 | ~v_644 | ~v_643 | ~v_642 | v_3022;
assign x_14656 = v_3021 | v_130;
assign x_14657 = v_3021 | v_19;
assign x_14658 = v_3020 | v_122;
assign x_14659 = v_3020 | v_19;
assign x_14660 = v_3019 | v_115;
assign x_14661 = v_3019 | ~v_19;
assign x_14662 = v_3018 | v_107;
assign x_14663 = v_3018 | ~v_19;
assign x_14664 = v_54 | v_61 | v_60 | v_59 | v_58 | v_57 | ~v_3016 | v_144 | v_142 | v_167 | v_166 | v_165 | v_183 | ~v_698 | ~v_697 | ~v_3015 | ~v_468 | ~v_2940 | ~v_467 | ~v_3014 | ~v_3013 | ~v_2937 | ~v_696 | ~v_638 | ~v_2968 | ~v_2967 | ~v_695 | ~v_637 | ~v_2966 | ~v_2965 | ~v_458 | ~v_457 | ~v_246 | ~v_2932 | ~v_2931 | ~v_456 | ~v_455 | ~v_243 | ~v_2930 | ~v_2929 | ~v_630 | ~v_629 | ~v_628 | ~v_627 | v_3017;
assign x_14665 = v_3016 | v_80;
assign x_14666 = v_3016 | v_19;
assign x_14667 = v_3015 | v_88;
assign x_14668 = v_3015 | v_19;
assign x_14669 = v_3014 | v_73;
assign x_14670 = v_3014 | ~v_19;
assign x_14671 = v_3013 | v_65;
assign x_14672 = v_3013 | ~v_19;
assign x_14673 = v_18 | v_17 | v_16 | v_15 | v_14 | v_11 | ~v_453 | ~v_2927 | ~v_452 | ~v_2926 | v_136 | v_134 | v_163 | v_162 | v_161 | v_182 | ~v_693 | ~v_692 | ~v_3011 | ~v_3010 | ~v_3009 | ~v_3008 | ~v_691 | ~v_623 | ~v_2963 | ~v_2962 | ~v_690 | ~v_622 | ~v_2961 | ~v_2960 | ~v_443 | ~v_442 | ~v_213 | ~v_2917 | ~v_2916 | ~v_441 | ~v_440 | ~v_210 | ~v_2915 | ~v_2914 | ~v_615 | ~v_614 | ~v_613 | ~v_612 | v_3012;
assign x_14674 = v_3011 | v_46;
assign x_14675 = v_3011 | v_19;
assign x_14676 = v_3010 | v_38;
assign x_14677 = v_3010 | v_19;
assign x_14678 = v_3009 | v_31;
assign x_14679 = v_3009 | ~v_19;
assign x_14680 = v_3008 | v_23;
assign x_14681 = v_3008 | ~v_19;
assign x_14682 = v_3007 | ~v_2996;
assign x_14683 = v_3007 | ~v_3001;
assign x_14684 = v_3007 | ~v_3006;
assign x_14685 = v_103 | v_97 | v_100 | v_151 | v_171 | v_170 | v_169 | v_160 | v_150 | v_148 | v_147 | v_184 | ~v_655 | ~v_654 | ~v_2955 | ~v_2952 | ~v_297 | ~v_3005 | ~v_3004 | ~v_296 | ~v_3003 | ~v_3002 | ~v_653 | ~v_2973 | ~v_2972 | ~v_652 | ~v_2971 | ~v_2970 | ~v_651 | ~v_650 | ~v_279 | ~v_2947 | ~v_2946 | ~v_276 | ~v_2945 | ~v_2944 | ~v_275 | ~v_274 | ~v_273 | ~v_272 | ~v_645 | ~v_644 | ~v_643 | ~v_642 | v_3006;
assign x_14686 = v_3005 | v_157;
assign x_14687 = v_3005 | v_130;
assign x_14688 = v_3004 | v_156;
assign x_14689 = v_3004 | v_122;
assign x_14690 = v_3003 | ~v_157;
assign x_14691 = v_3003 | v_115;
assign x_14692 = v_3002 | ~v_156;
assign x_14693 = v_3002 | v_107;
assign x_14694 = v_55 | v_61 | v_58 | v_159 | v_145 | v_143 | v_142 | v_167 | v_166 | v_165 | v_146 | v_183 | ~v_640 | ~v_639 | ~v_2940 | ~v_2937 | ~v_264 | ~v_3000 | ~v_2999 | ~v_263 | ~v_2998 | ~v_2997 | ~v_638 | ~v_2968 | ~v_2967 | ~v_637 | ~v_2966 | ~v_2965 | ~v_636 | ~v_635 | ~v_246 | ~v_2932 | ~v_2931 | ~v_243 | ~v_2930 | ~v_2929 | ~v_242 | ~v_241 | ~v_240 | ~v_239 | ~v_630 | ~v_629 | ~v_628 | ~v_627 | v_3001;
assign x_14695 = v_3000 | v_157;
assign x_14696 = v_3000 | v_88;
assign x_14697 = v_2999 | v_156;
assign x_14698 = v_2999 | v_80;
assign x_14699 = v_2998 | ~v_157;
assign x_14700 = v_2998 | v_73;
assign x_14701 = v_2997 | ~v_156;
assign x_14702 = v_2997 | v_65;
assign x_14703 = v_18 | v_15 | v_12 | ~v_2927 | ~v_2926 | v_135 | v_134 | v_137 | v_138 | v_163 | v_162 | v_161 | v_155 | v_182 | ~v_625 | ~v_624 | ~v_231 | ~v_2995 | ~v_2994 | ~v_230 | ~v_2993 | ~v_2992 | ~v_623 | ~v_2963 | ~v_2962 | ~v_622 | ~v_2961 | ~v_2960 | ~v_621 | ~v_620 | ~v_213 | ~v_2917 | ~v_2916 | ~v_210 | ~v_2915 | ~v_2914 | ~v_209 | ~v_208 | ~v_207 | ~v_206 | ~v_615 | ~v_614 | ~v_613 | ~v_612 | v_2996;
assign x_14704 = v_2995 | v_157;
assign x_14705 = v_2995 | v_46;
assign x_14706 = v_2994 | v_156;
assign x_14707 = v_2994 | v_38;
assign x_14708 = v_2993 | ~v_157;
assign x_14709 = v_2993 | v_31;
assign x_14710 = v_2992 | ~v_156;
assign x_14711 = v_2992 | v_23;
assign x_14712 = v_2991 | ~v_2980;
assign x_14713 = v_2991 | ~v_2985;
assign x_14714 = v_2991 | ~v_2990;
assign x_14715 = v_101 | v_100 | v_102 | v_172 | v_171 | v_170 | v_169 | v_150 | v_149 | v_148 | v_147 | v_184 | ~v_389 | ~v_388 | ~v_671 | ~v_670 | ~v_2955 | ~v_2952 | ~v_387 | ~v_2989 | ~v_2988 | ~v_386 | ~v_2987 | ~v_2986 | ~v_653 | ~v_2973 | ~v_2972 | ~v_652 | ~v_2971 | ~v_2970 | ~v_669 | ~v_668 | ~v_279 | ~v_2947 | ~v_2946 | ~v_276 | ~v_2945 | ~v_2944 | ~v_379 | ~v_378 | ~v_645 | ~v_644 | ~v_643 | ~v_642 | v_2990;
assign x_14716 = v_2989 | v_140;
assign x_14717 = v_2989 | v_130;
assign x_14718 = v_2988 | v_139;
assign x_14719 = v_2988 | v_122;
assign x_14720 = v_2987 | ~v_140;
assign x_14721 = v_2987 | v_115;
assign x_14722 = v_2986 | ~v_139;
assign x_14723 = v_2986 | v_107;
assign x_14724 = v_60 | v_59 | v_58 | v_144 | v_145 | v_143 | v_142 | v_168 | v_167 | v_166 | v_165 | v_183 | ~v_374 | ~v_373 | ~v_666 | ~v_665 | ~v_2940 | ~v_2937 | ~v_372 | ~v_2984 | ~v_2983 | ~v_371 | ~v_2982 | ~v_2981 | ~v_638 | ~v_2968 | ~v_2967 | ~v_637 | ~v_2966 | ~v_2965 | ~v_664 | ~v_663 | ~v_246 | ~v_2932 | ~v_2931 | ~v_243 | ~v_2930 | ~v_2929 | ~v_364 | ~v_363 | ~v_630 | ~v_629 | ~v_628 | ~v_627 | v_2985;
assign x_14725 = v_2984 | v_140;
assign x_14726 = v_2984 | v_88;
assign x_14727 = v_2983 | v_139;
assign x_14728 = v_2983 | v_80;
assign x_14729 = v_2982 | ~v_140;
assign x_14730 = v_2982 | v_73;
assign x_14731 = v_2981 | ~v_139;
assign x_14732 = v_2981 | v_65;
assign x_14733 = v_17 | v_16 | v_15 | ~v_2927 | ~v_2926 | v_136 | v_135 | v_134 | v_137 | v_164 | v_163 | v_162 | v_161 | v_182 | ~v_359 | ~v_358 | ~v_661 | ~v_660 | ~v_357 | ~v_2979 | ~v_2978 | ~v_356 | ~v_2977 | ~v_2976 | ~v_623 | ~v_2963 | ~v_2962 | ~v_622 | ~v_2961 | ~v_2960 | ~v_659 | ~v_658 | ~v_213 | ~v_2917 | ~v_2916 | ~v_210 | ~v_2915 | ~v_2914 | ~v_349 | ~v_348 | ~v_615 | ~v_614 | ~v_613 | ~v_612 | v_2980;
assign x_14734 = v_2979 | v_140;
assign x_14735 = v_2979 | v_46;
assign x_14736 = v_2978 | v_139;
assign x_14737 = v_2978 | v_38;
assign x_14738 = v_2977 | ~v_140;
assign x_14739 = v_2977 | v_31;
assign x_14740 = v_2976 | ~v_139;
assign x_14741 = v_2976 | v_23;
assign x_14742 = v_2975 | ~v_2964;
assign x_14743 = v_2975 | ~v_2969;
assign x_14744 = v_2975 | ~v_2974;
assign x_14745 = v_103 | v_101 | v_100 | v_95 | v_102 | v_171 | v_170 | v_169 | v_150 | v_149 | v_148 | v_184 | ~v_2955 | ~v_2952 | ~v_435 | ~v_2951 | ~v_2950 | ~v_434 | ~v_2949 | ~v_2948 | ~v_653 | ~v_2973 | ~v_2972 | ~v_652 | ~v_2971 | ~v_2970 | ~v_687 | ~v_686 | ~v_685 | ~v_684 | ~v_279 | ~v_2947 | ~v_2946 | ~v_276 | ~v_2945 | ~v_2944 | ~v_427 | ~v_426 | ~v_425 | ~v_424 | ~v_645 | ~v_644 | ~v_643 | ~v_642 | v_2974;
assign x_14746 = v_2973 | v_153;
assign x_14747 = v_2973 | v_127;
assign x_14748 = v_2972 | v_152;
assign x_14749 = v_2972 | v_121;
assign x_14750 = v_2971 | ~v_153;
assign x_14751 = v_2971 | v_112;
assign x_14752 = v_2970 | ~v_152;
assign x_14753 = v_2970 | v_106;
assign x_14754 = v_53 | v_61 | v_60 | v_59 | v_58 | v_144 | v_145 | v_143 | v_167 | v_166 | v_165 | v_183 | ~v_2940 | ~v_2937 | ~v_420 | ~v_2936 | ~v_2935 | ~v_419 | ~v_2934 | ~v_2933 | ~v_638 | ~v_2968 | ~v_2967 | ~v_637 | ~v_2966 | ~v_2965 | ~v_682 | ~v_681 | ~v_680 | ~v_679 | ~v_246 | ~v_2932 | ~v_2931 | ~v_243 | ~v_2930 | ~v_2929 | ~v_412 | ~v_411 | ~v_410 | ~v_409 | ~v_630 | ~v_629 | ~v_628 | ~v_627 | v_2969;
assign x_14755 = v_2968 | v_153;
assign x_14756 = v_2968 | v_85;
assign x_14757 = v_2967 | v_152;
assign x_14758 = v_2967 | v_79;
assign x_14759 = v_2966 | ~v_153;
assign x_14760 = v_2966 | v_70;
assign x_14761 = v_2965 | ~v_152;
assign x_14762 = v_2965 | v_64;
assign x_14763 = v_18 | v_17 | v_16 | v_15 | v_10 | ~v_2927 | ~v_2926 | v_136 | v_135 | v_137 | v_163 | v_162 | v_161 | v_182 | ~v_405 | ~v_2921 | ~v_2920 | ~v_404 | ~v_2919 | ~v_2918 | ~v_623 | ~v_2963 | ~v_2962 | ~v_622 | ~v_2961 | ~v_2960 | ~v_677 | ~v_676 | ~v_675 | ~v_674 | ~v_213 | ~v_2917 | ~v_2916 | ~v_210 | ~v_2915 | ~v_2914 | ~v_397 | ~v_396 | ~v_395 | ~v_394 | ~v_615 | ~v_614 | ~v_613 | ~v_612 | v_2964;
assign x_14764 = v_2963 | v_153;
assign x_14765 = v_2963 | v_43;
assign x_14766 = v_2962 | v_152;
assign x_14767 = v_2962 | v_37;
assign x_14768 = v_2961 | ~v_153;
assign x_14769 = v_2961 | v_28;
assign x_14770 = v_2960 | ~v_152;
assign x_14771 = v_2960 | v_22;
assign x_14772 = v_2959 | ~v_2928;
assign x_14773 = v_2959 | ~v_2943;
assign x_14774 = v_2959 | ~v_2958;
assign x_14775 = v_98 | v_103 | v_101 | v_100 | v_93 | v_102 | v_170 | v_150 | v_149 | v_148 | v_147 | v_184 | ~v_609 | ~v_608 | ~v_299 | ~v_2957 | ~v_2956 | ~v_2955 | ~v_298 | ~v_2954 | ~v_2953 | ~v_2952 | ~v_435 | ~v_2951 | ~v_2950 | ~v_434 | ~v_2949 | ~v_2948 | ~v_607 | ~v_606 | ~v_281 | ~v_280 | ~v_279 | ~v_2947 | ~v_2946 | ~v_278 | ~v_277 | ~v_276 | ~v_2945 | ~v_2944 | ~v_427 | ~v_426 | ~v_425 | ~v_424 | v_2958;
assign x_14776 = v_2957 | v_127;
assign x_14777 = v_2957 | v_19;
assign x_14778 = v_2956 | v_121;
assign x_14779 = v_2956 | v_19;
assign x_14780 = v_2955 | v_119;
assign x_14781 = v_2955 | v_19;
assign x_14782 = v_2954 | v_112;
assign x_14783 = v_2954 | ~v_19;
assign x_14784 = v_2953 | v_106;
assign x_14785 = v_2953 | ~v_19;
assign x_14786 = v_2952 | v_104;
assign x_14787 = v_2952 | ~v_19;
assign x_14788 = v_2951 | v_153;
assign x_14789 = v_2951 | v_130;
assign x_14790 = v_2950 | v_152;
assign x_14791 = v_2950 | v_122;
assign x_14792 = v_2949 | ~v_153;
assign x_14793 = v_2949 | v_115;
assign x_14794 = v_2948 | ~v_152;
assign x_14795 = v_2948 | v_107;
assign x_14796 = v_2947 | v_157;
assign x_14797 = v_2947 | v_123;
assign x_14798 = v_2946 | v_156;
assign x_14799 = v_2946 | v_120;
assign x_14800 = v_2945 | ~v_157;
assign x_14801 = v_2945 | v_108;
assign x_14802 = v_2944 | ~v_156;
assign x_14803 = v_2944 | v_105;
assign x_14804 = v_56 | v_61 | v_51 | v_60 | v_59 | v_58 | v_144 | v_145 | v_143 | v_142 | v_166 | v_183 | ~v_604 | ~v_603 | ~v_266 | ~v_2942 | ~v_2941 | ~v_2940 | ~v_265 | ~v_2939 | ~v_2938 | ~v_2937 | ~v_420 | ~v_2936 | ~v_2935 | ~v_419 | ~v_2934 | ~v_2933 | ~v_602 | ~v_601 | ~v_248 | ~v_247 | ~v_246 | ~v_2932 | ~v_2931 | ~v_245 | ~v_244 | ~v_243 | ~v_2930 | ~v_2929 | ~v_412 | ~v_411 | ~v_410 | ~v_409 | v_2943;
assign x_14805 = v_2942 | v_85;
assign x_14806 = v_2942 | v_19;
assign x_14807 = v_2941 | v_79;
assign x_14808 = v_2941 | v_19;
assign x_14809 = v_2940 | v_77;
assign x_14810 = v_2940 | v_19;
assign x_14811 = v_2939 | v_70;
assign x_14812 = v_2939 | ~v_19;
assign x_14813 = v_2938 | v_64;
assign x_14814 = v_2938 | ~v_19;
assign x_14815 = v_2937 | v_62;
assign x_14816 = v_2937 | ~v_19;
assign x_14817 = v_2936 | v_153;
assign x_14818 = v_2936 | v_88;
assign x_14819 = v_2935 | v_152;
assign x_14820 = v_2935 | v_80;
assign x_14821 = v_2934 | ~v_153;
assign x_14822 = v_2934 | v_73;
assign x_14823 = v_2933 | ~v_152;
assign x_14824 = v_2933 | v_65;
assign x_14825 = v_2932 | v_157;
assign x_14826 = v_2932 | v_81;
assign x_14827 = v_2931 | v_156;
assign x_14828 = v_2931 | v_78;
assign x_14829 = v_2930 | ~v_157;
assign x_14830 = v_2930 | v_66;
assign x_14831 = v_2929 | ~v_156;
assign x_14832 = v_2929 | v_63;
assign x_14833 = v_13 | v_18 | v_17 | v_16 | v_8 | v_15 | ~v_2927 | ~v_2926 | v_136 | v_135 | v_134 | v_137 | v_162 | v_182 | ~v_599 | ~v_598 | ~v_233 | ~v_2925 | ~v_2924 | ~v_232 | ~v_2923 | ~v_2922 | ~v_405 | ~v_2921 | ~v_2920 | ~v_404 | ~v_2919 | ~v_2918 | ~v_597 | ~v_596 | ~v_215 | ~v_214 | ~v_213 | ~v_2917 | ~v_2916 | ~v_212 | ~v_211 | ~v_210 | ~v_2915 | ~v_2914 | ~v_397 | ~v_396 | ~v_395 | ~v_394 | v_2928;
assign x_14834 = v_2927 | v_35;
assign x_14835 = v_2927 | v_19;
assign x_14836 = v_2926 | v_20;
assign x_14837 = v_2926 | ~v_19;
assign x_14838 = v_2925 | v_43;
assign x_14839 = v_2925 | v_19;
assign x_14840 = v_2924 | v_37;
assign x_14841 = v_2924 | v_19;
assign x_14842 = v_2923 | v_28;
assign x_14843 = v_2923 | ~v_19;
assign x_14844 = v_2922 | v_22;
assign x_14845 = v_2922 | ~v_19;
assign x_14846 = v_2921 | v_153;
assign x_14847 = v_2921 | v_46;
assign x_14848 = v_2920 | v_152;
assign x_14849 = v_2920 | v_38;
assign x_14850 = v_2919 | ~v_153;
assign x_14851 = v_2919 | v_31;
assign x_14852 = v_2918 | ~v_152;
assign x_14853 = v_2918 | v_23;
assign x_14854 = v_2917 | v_157;
assign x_14855 = v_2917 | v_39;
assign x_14856 = v_2916 | v_156;
assign x_14857 = v_2916 | v_36;
assign x_14858 = v_2915 | ~v_157;
assign x_14859 = v_2915 | v_24;
assign x_14860 = v_2914 | ~v_156;
assign x_14861 = v_2914 | v_21;
assign x_14862 = v_2913 | ~v_2911;
assign x_14863 = v_2913 | ~v_2912;
assign x_14864 = v_2913 | ~v_194;
assign x_14865 = v_2913 | ~v_196;
assign x_14866 = v_2913 | ~v_157;
assign x_14867 = v_2913 | ~v_156;
assign x_14868 = ~v_186 | ~v_191 | v_2912;
assign x_14869 = ~v_193 | ~v_1851 | v_2911;
assign x_14870 = v_2910 | ~v_2829;
assign x_14871 = v_2910 | ~v_2909;
assign x_14872 = v_174 | v_173 | ~v_2908 | ~v_1561 | ~v_1560 | ~v_2831 | ~v_2830 | v_2909;
assign x_14873 = v_2908 | ~v_2847;
assign x_14874 = v_2908 | ~v_2851;
assign x_14875 = v_2908 | ~v_2855;
assign x_14876 = v_2908 | ~v_2859;
assign x_14877 = v_2908 | ~v_2863;
assign x_14878 = v_2908 | ~v_2867;
assign x_14879 = v_2908 | ~v_2871;
assign x_14880 = v_2908 | ~v_2875;
assign x_14881 = v_2908 | ~v_2879;
assign x_14882 = v_2908 | ~v_2883;
assign x_14883 = v_2908 | ~v_2887;
assign x_14884 = v_2908 | ~v_2891;
assign x_14885 = v_2908 | ~v_2895;
assign x_14886 = v_2908 | ~v_2899;
assign x_14887 = v_2908 | ~v_2903;
assign x_14888 = v_2908 | ~v_2907;
assign x_14889 = v_2908 | ~v_1263;
assign x_14890 = v_2908 | ~v_1264;
assign x_14891 = v_2908 | ~v_1265;
assign x_14892 = v_2908 | ~v_1266;
assign x_14893 = ~v_2906 | ~v_2905 | ~v_2904 | v_2907;
assign x_14894 = v_2906 | ~v_2842;
assign x_14895 = v_2906 | ~v_2843;
assign x_14896 = v_2906 | ~v_2844;
assign x_14897 = v_2906 | ~v_2845;
assign x_14898 = v_2906 | ~v_827;
assign x_14899 = v_2906 | ~v_828;
assign x_14900 = v_2906 | ~v_1015;
assign x_14901 = v_2906 | ~v_829;
assign x_14902 = v_2906 | ~v_1016;
assign x_14903 = v_2906 | ~v_830;
assign x_14904 = v_2906 | ~v_831;
assign x_14905 = v_2906 | ~v_1017;
assign x_14906 = v_2906 | ~v_832;
assign x_14907 = v_2906 | ~v_1018;
assign x_14908 = v_2906 | ~v_839;
assign x_14909 = v_2906 | ~v_1257;
assign x_14910 = v_2906 | ~v_1023;
assign x_14911 = v_2906 | ~v_840;
assign x_14912 = v_2906 | ~v_1258;
assign x_14913 = v_2906 | ~v_1024;
assign x_14914 = v_2906 | ~v_2446;
assign x_14915 = v_2906 | ~v_2447;
assign x_14916 = v_2906 | ~v_2512;
assign x_14917 = v_2906 | ~v_2448;
assign x_14918 = v_2906 | ~v_2513;
assign x_14919 = v_2906 | ~v_2449;
assign x_14920 = v_2906 | ~v_2450;
assign x_14921 = v_2906 | ~v_2514;
assign x_14922 = v_2906 | ~v_2451;
assign x_14923 = v_2906 | ~v_2515;
assign x_14924 = v_2906 | ~v_184;
assign x_14925 = v_2906 | ~v_170;
assign x_14926 = v_2906 | ~v_169;
assign x_14927 = v_2906 | ~v_149;
assign x_14928 = v_2906 | ~v_148;
assign x_14929 = v_2906 | ~v_1259;
assign x_14930 = v_2906 | ~v_1260;
assign x_14931 = v_2906 | ~v_103;
assign x_14932 = v_2906 | ~v_102;
assign x_14933 = v_2906 | ~v_101;
assign x_14934 = v_2906 | ~v_100;
assign x_14935 = v_2906 | ~v_99;
assign x_14936 = v_2906 | ~v_98;
assign x_14937 = v_2906 | ~v_95;
assign x_14938 = v_2905 | ~v_2837;
assign x_14939 = v_2905 | ~v_2838;
assign x_14940 = v_2905 | ~v_2839;
assign x_14941 = v_2905 | ~v_2840;
assign x_14942 = v_2905 | ~v_794;
assign x_14943 = v_2905 | ~v_795;
assign x_14944 = v_2905 | ~v_1000;
assign x_14945 = v_2905 | ~v_796;
assign x_14946 = v_2905 | ~v_1001;
assign x_14947 = v_2905 | ~v_797;
assign x_14948 = v_2905 | ~v_798;
assign x_14949 = v_2905 | ~v_1002;
assign x_14950 = v_2905 | ~v_799;
assign x_14951 = v_2905 | ~v_1003;
assign x_14952 = v_2905 | ~v_806;
assign x_14953 = v_2905 | ~v_1252;
assign x_14954 = v_2905 | ~v_1008;
assign x_14955 = v_2905 | ~v_1253;
assign x_14956 = v_2905 | ~v_1009;
assign x_14957 = v_2905 | ~v_2431;
assign x_14958 = v_2905 | ~v_2432;
assign x_14959 = v_2905 | ~v_2507;
assign x_14960 = v_2905 | ~v_2433;
assign x_14961 = v_2905 | ~v_2508;
assign x_14962 = v_2905 | ~v_2434;
assign x_14963 = v_2905 | ~v_2435;
assign x_14964 = v_2905 | ~v_2509;
assign x_14965 = v_2905 | ~v_2436;
assign x_14966 = v_2905 | ~v_2510;
assign x_14967 = v_2905 | ~v_807;
assign x_14968 = v_2905 | ~v_183;
assign x_14969 = v_2905 | ~v_166;
assign x_14970 = v_2905 | ~v_165;
assign x_14971 = v_2905 | ~v_144;
assign x_14972 = v_2905 | ~v_143;
assign x_14973 = v_2905 | ~v_1254;
assign x_14974 = v_2905 | ~v_1255;
assign x_14975 = v_2905 | ~v_61;
assign x_14976 = v_2905 | ~v_60;
assign x_14977 = v_2905 | ~v_59;
assign x_14978 = v_2905 | ~v_58;
assign x_14979 = v_2905 | ~v_57;
assign x_14980 = v_2905 | ~v_56;
assign x_14981 = v_2905 | ~v_53;
assign x_14982 = v_2904 | ~v_2832;
assign x_14983 = v_2904 | ~v_2833;
assign x_14984 = v_2904 | ~v_2834;
assign x_14985 = v_2904 | ~v_2835;
assign x_14986 = v_2904 | ~v_761;
assign x_14987 = v_2904 | ~v_762;
assign x_14988 = v_2904 | ~v_985;
assign x_14989 = v_2904 | ~v_763;
assign x_14990 = v_2904 | ~v_986;
assign x_14991 = v_2904 | ~v_764;
assign x_14992 = v_2904 | ~v_765;
assign x_14993 = v_2904 | ~v_987;
assign x_14994 = v_2904 | ~v_766;
assign x_14995 = v_2904 | ~v_988;
assign x_14996 = v_2904 | ~v_773;
assign x_14997 = v_2904 | ~v_774;
assign x_14998 = v_2904 | ~v_2416;
assign x_14999 = v_2904 | ~v_2417;
assign x_15000 = v_2904 | ~v_2502;
assign x_15001 = v_2904 | ~v_2418;
assign x_15002 = v_2904 | ~v_2503;
assign x_15003 = v_2904 | ~v_2419;
assign x_15004 = v_2904 | ~v_2420;
assign x_15005 = v_2904 | ~v_2504;
assign x_15006 = v_2904 | ~v_2421;
assign x_15007 = v_2904 | ~v_2505;
assign x_15008 = v_2904 | ~v_182;
assign x_15009 = v_2904 | ~v_162;
assign x_15010 = v_2904 | ~v_161;
assign x_15011 = v_2904 | ~v_1247;
assign x_15012 = v_2904 | ~v_1248;
assign x_15013 = v_2904 | ~v_136;
assign x_15014 = v_2904 | ~v_135;
assign x_15015 = v_2904 | ~v_1249;
assign x_15016 = v_2904 | ~v_993;
assign x_15017 = v_2904 | ~v_1250;
assign x_15018 = v_2904 | ~v_994;
assign x_15019 = v_2904 | ~v_18;
assign x_15020 = v_2904 | ~v_17;
assign x_15021 = v_2904 | ~v_16;
assign x_15022 = v_2904 | ~v_15;
assign x_15023 = v_2904 | ~v_14;
assign x_15024 = v_2904 | ~v_13;
assign x_15025 = v_2904 | ~v_10;
assign x_15026 = ~v_2902 | ~v_2901 | ~v_2900 | v_2903;
assign x_15027 = v_2902 | ~v_2842;
assign x_15028 = v_2902 | ~v_2843;
assign x_15029 = v_2902 | ~v_2844;
assign x_15030 = v_2902 | ~v_2845;
assign x_15031 = v_2902 | ~v_1187;
assign x_15032 = v_2902 | ~v_1188;
assign x_15033 = v_2902 | ~v_1189;
assign x_15034 = v_2902 | ~v_1190;
assign x_15035 = v_2902 | ~v_827;
assign x_15036 = v_2902 | ~v_1015;
assign x_15037 = v_2902 | ~v_1016;
assign x_15038 = v_2902 | ~v_830;
assign x_15039 = v_2902 | ~v_1017;
assign x_15040 = v_2902 | ~v_1018;
assign x_15041 = v_2902 | ~v_1193;
assign x_15042 = v_2902 | ~v_1241;
assign x_15043 = v_2902 | ~v_1194;
assign x_15044 = v_2902 | ~v_1242;
assign x_15045 = v_2902 | ~v_2464;
assign x_15046 = v_2902 | ~v_2465;
assign x_15047 = v_2902 | ~v_2466;
assign x_15048 = v_2902 | ~v_2467;
assign x_15049 = v_2902 | ~v_1023;
assign x_15050 = v_2902 | ~v_1024;
assign x_15051 = v_2902 | ~v_2446;
assign x_15052 = v_2902 | ~v_2512;
assign x_15053 = v_2902 | ~v_2513;
assign x_15054 = v_2902 | ~v_2449;
assign x_15055 = v_2902 | ~v_2514;
assign x_15056 = v_2902 | ~v_2515;
assign x_15057 = v_2902 | ~v_1243;
assign x_15058 = v_2902 | ~v_1244;
assign x_15059 = v_2902 | ~v_184;
assign x_15060 = v_2902 | ~v_171;
assign x_15061 = v_2902 | ~v_170;
assign x_15062 = v_2902 | ~v_149;
assign x_15063 = v_2902 | ~v_148;
assign x_15064 = v_2902 | ~v_147;
assign x_15065 = v_2902 | ~v_103;
assign x_15066 = v_2902 | ~v_102;
assign x_15067 = v_2902 | ~v_101;
assign x_15068 = v_2902 | ~v_100;
assign x_15069 = v_2902 | ~v_99;
assign x_15070 = v_2902 | ~v_93;
assign x_15071 = v_2901 | ~v_2837;
assign x_15072 = v_2901 | ~v_2838;
assign x_15073 = v_2901 | ~v_2839;
assign x_15074 = v_2901 | ~v_2840;
assign x_15075 = v_2901 | ~v_1172;
assign x_15076 = v_2901 | ~v_1173;
assign x_15077 = v_2901 | ~v_1174;
assign x_15078 = v_2901 | ~v_1175;
assign x_15079 = v_2901 | ~v_794;
assign x_15080 = v_2901 | ~v_1000;
assign x_15081 = v_2901 | ~v_1001;
assign x_15082 = v_2901 | ~v_797;
assign x_15083 = v_2901 | ~v_1002;
assign x_15084 = v_2901 | ~v_1003;
assign x_15085 = v_2901 | ~v_1178;
assign x_15086 = v_2901 | ~v_1236;
assign x_15087 = v_2901 | ~v_1179;
assign x_15088 = v_2901 | ~v_1237;
assign x_15089 = v_2901 | ~v_2459;
assign x_15090 = v_2901 | ~v_2460;
assign x_15091 = v_2901 | ~v_2461;
assign x_15092 = v_2901 | ~v_2462;
assign x_15093 = v_2901 | ~v_1008;
assign x_15094 = v_2901 | ~v_1009;
assign x_15095 = v_2901 | ~v_2431;
assign x_15096 = v_2901 | ~v_2507;
assign x_15097 = v_2901 | ~v_2508;
assign x_15098 = v_2901 | ~v_2434;
assign x_15099 = v_2901 | ~v_2509;
assign x_15100 = v_2901 | ~v_2510;
assign x_15101 = v_2901 | ~v_1238;
assign x_15102 = v_2901 | ~v_1239;
assign x_15103 = v_2901 | ~v_183;
assign x_15104 = v_2901 | ~v_167;
assign x_15105 = v_2901 | ~v_166;
assign x_15106 = v_2901 | ~v_144;
assign x_15107 = v_2901 | ~v_143;
assign x_15108 = v_2901 | ~v_142;
assign x_15109 = v_2901 | ~v_61;
assign x_15110 = v_2901 | ~v_60;
assign x_15111 = v_2901 | ~v_59;
assign x_15112 = v_2901 | ~v_58;
assign x_15113 = v_2901 | ~v_57;
assign x_15114 = v_2901 | ~v_51;
assign x_15115 = v_2900 | ~v_2832;
assign x_15116 = v_2900 | ~v_2833;
assign x_15117 = v_2900 | ~v_2834;
assign x_15118 = v_2900 | ~v_2835;
assign x_15119 = v_2900 | ~v_1157;
assign x_15120 = v_2900 | ~v_1158;
assign x_15121 = v_2900 | ~v_1159;
assign x_15122 = v_2900 | ~v_1160;
assign x_15123 = v_2900 | ~v_761;
assign x_15124 = v_2900 | ~v_985;
assign x_15125 = v_2900 | ~v_986;
assign x_15126 = v_2900 | ~v_764;
assign x_15127 = v_2900 | ~v_987;
assign x_15128 = v_2900 | ~v_988;
assign x_15129 = v_2900 | ~v_1163;
assign x_15130 = v_2900 | ~v_1231;
assign x_15131 = v_2900 | ~v_1164;
assign x_15132 = v_2900 | ~v_1232;
assign x_15133 = v_2900 | ~v_2454;
assign x_15134 = v_2900 | ~v_2455;
assign x_15135 = v_2900 | ~v_2456;
assign x_15136 = v_2900 | ~v_2457;
assign x_15137 = v_2900 | ~v_2416;
assign x_15138 = v_2900 | ~v_2502;
assign x_15139 = v_2900 | ~v_2503;
assign x_15140 = v_2900 | ~v_2419;
assign x_15141 = v_2900 | ~v_2504;
assign x_15142 = v_2900 | ~v_2505;
assign x_15143 = v_2900 | ~v_1233;
assign x_15144 = v_2900 | ~v_1234;
assign x_15145 = v_2900 | ~v_182;
assign x_15146 = v_2900 | ~v_163;
assign x_15147 = v_2900 | ~v_162;
assign x_15148 = v_2900 | ~v_136;
assign x_15149 = v_2900 | ~v_135;
assign x_15150 = v_2900 | ~v_134;
assign x_15151 = v_2900 | ~v_993;
assign x_15152 = v_2900 | ~v_994;
assign x_15153 = v_2900 | ~v_18;
assign x_15154 = v_2900 | ~v_17;
assign x_15155 = v_2900 | ~v_16;
assign x_15156 = v_2900 | ~v_15;
assign x_15157 = v_2900 | ~v_14;
assign x_15158 = v_2900 | ~v_8;
assign x_15159 = ~v_2898 | ~v_2897 | ~v_2896 | v_2899;
assign x_15160 = v_2898 | ~v_2842;
assign x_15161 = v_2898 | ~v_2843;
assign x_15162 = v_2898 | ~v_2844;
assign x_15163 = v_2898 | ~v_2845;
assign x_15164 = v_2898 | ~v_969;
assign x_15165 = v_2898 | ~v_970;
assign x_15166 = v_2898 | ~v_971;
assign x_15167 = v_2898 | ~v_972;
assign x_15168 = v_2898 | ~v_1187;
assign x_15169 = v_2898 | ~v_1188;
assign x_15170 = v_2898 | ~v_1189;
assign x_15171 = v_2898 | ~v_1190;
assign x_15172 = v_2898 | ~v_827;
assign x_15173 = v_2898 | ~v_830;
assign x_15174 = v_2898 | ~v_1225;
assign x_15175 = v_2898 | ~v_1226;
assign x_15176 = v_2898 | ~v_1227;
assign x_15177 = v_2898 | ~v_1228;
assign x_15178 = v_2898 | ~v_1193;
assign x_15179 = v_2898 | ~v_1194;
assign x_15180 = v_2898 | ~v_2464;
assign x_15181 = v_2898 | ~v_2465;
assign x_15182 = v_2898 | ~v_2466;
assign x_15183 = v_2898 | ~v_2467;
assign x_15184 = v_2898 | ~v_975;
assign x_15185 = v_2898 | ~v_976;
assign x_15186 = v_2898 | ~v_2442;
assign x_15187 = v_2898 | ~v_2443;
assign x_15188 = v_2898 | ~v_2444;
assign x_15189 = v_2898 | ~v_2445;
assign x_15190 = v_2898 | ~v_2446;
assign x_15191 = v_2898 | ~v_2449;
assign x_15192 = v_2898 | ~v_184;
assign x_15193 = v_2898 | ~v_171;
assign x_15194 = v_2898 | ~v_170;
assign x_15195 = v_2898 | ~v_150;
assign x_15196 = v_2898 | ~v_149;
assign x_15197 = v_2898 | ~v_103;
assign x_15198 = v_2898 | ~v_102;
assign x_15199 = v_2898 | ~v_101;
assign x_15200 = v_2898 | ~v_100;
assign x_15201 = v_2898 | ~v_96;
assign x_15202 = v_2898 | ~v_95;
assign x_15203 = v_2898 | ~v_93;
assign x_15204 = v_2897 | ~v_2837;
assign x_15205 = v_2897 | ~v_2838;
assign x_15206 = v_2897 | ~v_2839;
assign x_15207 = v_2897 | ~v_2840;
assign x_15208 = v_2897 | ~v_954;
assign x_15209 = v_2897 | ~v_955;
assign x_15210 = v_2897 | ~v_956;
assign x_15211 = v_2897 | ~v_957;
assign x_15212 = v_2897 | ~v_1172;
assign x_15213 = v_2897 | ~v_1173;
assign x_15214 = v_2897 | ~v_1174;
assign x_15215 = v_2897 | ~v_1175;
assign x_15216 = v_2897 | ~v_794;
assign x_15217 = v_2897 | ~v_797;
assign x_15218 = v_2897 | ~v_1220;
assign x_15219 = v_2897 | ~v_1221;
assign x_15220 = v_2897 | ~v_1222;
assign x_15221 = v_2897 | ~v_1223;
assign x_15222 = v_2897 | ~v_1178;
assign x_15223 = v_2897 | ~v_1179;
assign x_15224 = v_2897 | ~v_2459;
assign x_15225 = v_2897 | ~v_2460;
assign x_15226 = v_2897 | ~v_2461;
assign x_15227 = v_2897 | ~v_2462;
assign x_15228 = v_2897 | ~v_960;
assign x_15229 = v_2897 | ~v_961;
assign x_15230 = v_2897 | ~v_2427;
assign x_15231 = v_2897 | ~v_2428;
assign x_15232 = v_2897 | ~v_2429;
assign x_15233 = v_2897 | ~v_2430;
assign x_15234 = v_2897 | ~v_2431;
assign x_15235 = v_2897 | ~v_2434;
assign x_15236 = v_2897 | ~v_183;
assign x_15237 = v_2897 | ~v_167;
assign x_15238 = v_2897 | ~v_166;
assign x_15239 = v_2897 | ~v_145;
assign x_15240 = v_2897 | ~v_144;
assign x_15241 = v_2897 | ~v_61;
assign x_15242 = v_2897 | ~v_60;
assign x_15243 = v_2897 | ~v_59;
assign x_15244 = v_2897 | ~v_58;
assign x_15245 = v_2897 | ~v_54;
assign x_15246 = v_2897 | ~v_53;
assign x_15247 = v_2897 | ~v_51;
assign x_15248 = v_2896 | ~v_2832;
assign x_15249 = v_2896 | ~v_2833;
assign x_15250 = v_2896 | ~v_2834;
assign x_15251 = v_2896 | ~v_2835;
assign x_15252 = v_2896 | ~v_939;
assign x_15253 = v_2896 | ~v_940;
assign x_15254 = v_2896 | ~v_941;
assign x_15255 = v_2896 | ~v_942;
assign x_15256 = v_2896 | ~v_1157;
assign x_15257 = v_2896 | ~v_1158;
assign x_15258 = v_2896 | ~v_1159;
assign x_15259 = v_2896 | ~v_1160;
assign x_15260 = v_2896 | ~v_761;
assign x_15261 = v_2896 | ~v_764;
assign x_15262 = v_2896 | ~v_1215;
assign x_15263 = v_2896 | ~v_1216;
assign x_15264 = v_2896 | ~v_1217;
assign x_15265 = v_2896 | ~v_1218;
assign x_15266 = v_2896 | ~v_1163;
assign x_15267 = v_2896 | ~v_1164;
assign x_15268 = v_2896 | ~v_2454;
assign x_15269 = v_2896 | ~v_2455;
assign x_15270 = v_2896 | ~v_2456;
assign x_15271 = v_2896 | ~v_2457;
assign x_15272 = v_2896 | ~v_945;
assign x_15273 = v_2896 | ~v_946;
assign x_15274 = v_2896 | ~v_2412;
assign x_15275 = v_2896 | ~v_2413;
assign x_15276 = v_2896 | ~v_2414;
assign x_15277 = v_2896 | ~v_2415;
assign x_15278 = v_2896 | ~v_2416;
assign x_15279 = v_2896 | ~v_2419;
assign x_15280 = v_2896 | ~v_182;
assign x_15281 = v_2896 | ~v_163;
assign x_15282 = v_2896 | ~v_162;
assign x_15283 = v_2896 | ~v_137;
assign x_15284 = v_2896 | ~v_136;
assign x_15285 = v_2896 | ~v_18;
assign x_15286 = v_2896 | ~v_17;
assign x_15287 = v_2896 | ~v_16;
assign x_15288 = v_2896 | ~v_15;
assign x_15289 = v_2896 | ~v_11;
assign x_15290 = v_2896 | ~v_10;
assign x_15291 = v_2896 | ~v_8;
assign x_15292 = ~v_2894 | ~v_2893 | ~v_2892 | v_2895;
assign x_15293 = v_2894 | ~v_2842;
assign x_15294 = v_2894 | ~v_2843;
assign x_15295 = v_2894 | ~v_2844;
assign x_15296 = v_2894 | ~v_2845;
assign x_15297 = v_2894 | ~v_921;
assign x_15298 = v_2894 | ~v_922;
assign x_15299 = v_2894 | ~v_923;
assign x_15300 = v_2894 | ~v_924;
assign x_15301 = v_2894 | ~v_1187;
assign x_15302 = v_2894 | ~v_1188;
assign x_15303 = v_2894 | ~v_1189;
assign x_15304 = v_2894 | ~v_1190;
assign x_15305 = v_2894 | ~v_827;
assign x_15306 = v_2894 | ~v_830;
assign x_15307 = v_2894 | ~v_1209;
assign x_15308 = v_2894 | ~v_1210;
assign x_15309 = v_2894 | ~v_1193;
assign x_15310 = v_2894 | ~v_1194;
assign x_15311 = v_2894 | ~v_2464;
assign x_15312 = v_2894 | ~v_2465;
assign x_15313 = v_2894 | ~v_2466;
assign x_15314 = v_2894 | ~v_2467;
assign x_15315 = v_2894 | ~v_927;
assign x_15316 = v_2894 | ~v_928;
assign x_15317 = v_2894 | ~v_2480;
assign x_15318 = v_2894 | ~v_2481;
assign x_15319 = v_2894 | ~v_2482;
assign x_15320 = v_2894 | ~v_2483;
assign x_15321 = v_2894 | ~v_2446;
assign x_15322 = v_2894 | ~v_2449;
assign x_15323 = v_2894 | ~v_1211;
assign x_15324 = v_2894 | ~v_1212;
assign x_15325 = v_2894 | ~v_184;
assign x_15326 = v_2894 | ~v_172;
assign x_15327 = v_2894 | ~v_171;
assign x_15328 = v_2894 | ~v_170;
assign x_15329 = v_2894 | ~v_150;
assign x_15330 = v_2894 | ~v_148;
assign x_15331 = v_2894 | ~v_147;
assign x_15332 = v_2894 | ~v_102;
assign x_15333 = v_2894 | ~v_101;
assign x_15334 = v_2894 | ~v_100;
assign x_15335 = v_2894 | ~v_97;
assign x_15336 = v_2894 | ~v_93;
assign x_15337 = v_2893 | ~v_2837;
assign x_15338 = v_2893 | ~v_2838;
assign x_15339 = v_2893 | ~v_2839;
assign x_15340 = v_2893 | ~v_2840;
assign x_15341 = v_2893 | ~v_906;
assign x_15342 = v_2893 | ~v_907;
assign x_15343 = v_2893 | ~v_908;
assign x_15344 = v_2893 | ~v_909;
assign x_15345 = v_2893 | ~v_1172;
assign x_15346 = v_2893 | ~v_1173;
assign x_15347 = v_2893 | ~v_1174;
assign x_15348 = v_2893 | ~v_1175;
assign x_15349 = v_2893 | ~v_794;
assign x_15350 = v_2893 | ~v_797;
assign x_15351 = v_2893 | ~v_1204;
assign x_15352 = v_2893 | ~v_1205;
assign x_15353 = v_2893 | ~v_1178;
assign x_15354 = v_2893 | ~v_1179;
assign x_15355 = v_2893 | ~v_2459;
assign x_15356 = v_2893 | ~v_2460;
assign x_15357 = v_2893 | ~v_2461;
assign x_15358 = v_2893 | ~v_2462;
assign x_15359 = v_2893 | ~v_912;
assign x_15360 = v_2893 | ~v_913;
assign x_15361 = v_2893 | ~v_2475;
assign x_15362 = v_2893 | ~v_2476;
assign x_15363 = v_2893 | ~v_2477;
assign x_15364 = v_2893 | ~v_2478;
assign x_15365 = v_2893 | ~v_2431;
assign x_15366 = v_2893 | ~v_2434;
assign x_15367 = v_2893 | ~v_1206;
assign x_15368 = v_2893 | ~v_1207;
assign x_15369 = v_2893 | ~v_183;
assign x_15370 = v_2893 | ~v_168;
assign x_15371 = v_2893 | ~v_167;
assign x_15372 = v_2893 | ~v_166;
assign x_15373 = v_2893 | ~v_145;
assign x_15374 = v_2893 | ~v_143;
assign x_15375 = v_2893 | ~v_142;
assign x_15376 = v_2893 | ~v_60;
assign x_15377 = v_2893 | ~v_59;
assign x_15378 = v_2893 | ~v_58;
assign x_15379 = v_2893 | ~v_55;
assign x_15380 = v_2893 | ~v_51;
assign x_15381 = v_2892 | ~v_2832;
assign x_15382 = v_2892 | ~v_2833;
assign x_15383 = v_2892 | ~v_2834;
assign x_15384 = v_2892 | ~v_2835;
assign x_15385 = v_2892 | ~v_891;
assign x_15386 = v_2892 | ~v_892;
assign x_15387 = v_2892 | ~v_893;
assign x_15388 = v_2892 | ~v_894;
assign x_15389 = v_2892 | ~v_1157;
assign x_15390 = v_2892 | ~v_1158;
assign x_15391 = v_2892 | ~v_1159;
assign x_15392 = v_2892 | ~v_1160;
assign x_15393 = v_2892 | ~v_761;
assign x_15394 = v_2892 | ~v_764;
assign x_15395 = v_2892 | ~v_1199;
assign x_15396 = v_2892 | ~v_1200;
assign x_15397 = v_2892 | ~v_1163;
assign x_15398 = v_2892 | ~v_1164;
assign x_15399 = v_2892 | ~v_2454;
assign x_15400 = v_2892 | ~v_2455;
assign x_15401 = v_2892 | ~v_2456;
assign x_15402 = v_2892 | ~v_2457;
assign x_15403 = v_2892 | ~v_897;
assign x_15404 = v_2892 | ~v_898;
assign x_15405 = v_2892 | ~v_2470;
assign x_15406 = v_2892 | ~v_2471;
assign x_15407 = v_2892 | ~v_2472;
assign x_15408 = v_2892 | ~v_2473;
assign x_15409 = v_2892 | ~v_2416;
assign x_15410 = v_2892 | ~v_2419;
assign x_15411 = v_2892 | ~v_1201;
assign x_15412 = v_2892 | ~v_1202;
assign x_15413 = v_2892 | ~v_182;
assign x_15414 = v_2892 | ~v_164;
assign x_15415 = v_2892 | ~v_163;
assign x_15416 = v_2892 | ~v_162;
assign x_15417 = v_2892 | ~v_137;
assign x_15418 = v_2892 | ~v_135;
assign x_15419 = v_2892 | ~v_134;
assign x_15420 = v_2892 | ~v_17;
assign x_15421 = v_2892 | ~v_16;
assign x_15422 = v_2892 | ~v_15;
assign x_15423 = v_2892 | ~v_12;
assign x_15424 = v_2892 | ~v_8;
assign x_15425 = ~v_2890 | ~v_2889 | ~v_2888 | v_2891;
assign x_15426 = v_2890 | ~v_2842;
assign x_15427 = v_2890 | ~v_2843;
assign x_15428 = v_2890 | ~v_2844;
assign x_15429 = v_2890 | ~v_2845;
assign x_15430 = v_2890 | ~v_823;
assign x_15431 = v_2890 | ~v_824;
assign x_15432 = v_2890 | ~v_825;
assign x_15433 = v_2890 | ~v_826;
assign x_15434 = v_2890 | ~v_1187;
assign x_15435 = v_2890 | ~v_1188;
assign x_15436 = v_2890 | ~v_1189;
assign x_15437 = v_2890 | ~v_1190;
assign x_15438 = v_2890 | ~v_827;
assign x_15439 = v_2890 | ~v_830;
assign x_15440 = v_2890 | ~v_1191;
assign x_15441 = v_2890 | ~v_1192;
assign x_15442 = v_2890 | ~v_1193;
assign x_15443 = v_2890 | ~v_1194;
assign x_15444 = v_2890 | ~v_2464;
assign x_15445 = v_2890 | ~v_2465;
assign x_15446 = v_2890 | ~v_2466;
assign x_15447 = v_2890 | ~v_2467;
assign x_15448 = v_2890 | ~v_837;
assign x_15449 = v_2890 | ~v_838;
assign x_15450 = v_2890 | ~v_2496;
assign x_15451 = v_2890 | ~v_2497;
assign x_15452 = v_2890 | ~v_2498;
assign x_15453 = v_2890 | ~v_2499;
assign x_15454 = v_2890 | ~v_2446;
assign x_15455 = v_2890 | ~v_2449;
assign x_15456 = v_2890 | ~v_1195;
assign x_15457 = v_2890 | ~v_1196;
assign x_15458 = v_2890 | ~v_184;
assign x_15459 = v_2890 | ~v_171;
assign x_15460 = v_2890 | ~v_170;
assign x_15461 = v_2890 | ~v_160;
assign x_15462 = v_2890 | ~v_151;
assign x_15463 = v_2890 | ~v_150;
assign x_15464 = v_2890 | ~v_149;
assign x_15465 = v_2890 | ~v_148;
assign x_15466 = v_2890 | ~v_147;
assign x_15467 = v_2890 | ~v_103;
assign x_15468 = v_2890 | ~v_100;
assign x_15469 = v_2890 | ~v_93;
assign x_15470 = v_2889 | ~v_2837;
assign x_15471 = v_2889 | ~v_2838;
assign x_15472 = v_2889 | ~v_2839;
assign x_15473 = v_2889 | ~v_2840;
assign x_15474 = v_2889 | ~v_790;
assign x_15475 = v_2889 | ~v_791;
assign x_15476 = v_2889 | ~v_792;
assign x_15477 = v_2889 | ~v_793;
assign x_15478 = v_2889 | ~v_1172;
assign x_15479 = v_2889 | ~v_1173;
assign x_15480 = v_2889 | ~v_1174;
assign x_15481 = v_2889 | ~v_1175;
assign x_15482 = v_2889 | ~v_794;
assign x_15483 = v_2889 | ~v_797;
assign x_15484 = v_2889 | ~v_1176;
assign x_15485 = v_2889 | ~v_1177;
assign x_15486 = v_2889 | ~v_1178;
assign x_15487 = v_2889 | ~v_1179;
assign x_15488 = v_2889 | ~v_2459;
assign x_15489 = v_2889 | ~v_2460;
assign x_15490 = v_2889 | ~v_2461;
assign x_15491 = v_2889 | ~v_2462;
assign x_15492 = v_2889 | ~v_804;
assign x_15493 = v_2889 | ~v_805;
assign x_15494 = v_2889 | ~v_2491;
assign x_15495 = v_2889 | ~v_2492;
assign x_15496 = v_2889 | ~v_2493;
assign x_15497 = v_2889 | ~v_2494;
assign x_15498 = v_2889 | ~v_2431;
assign x_15499 = v_2889 | ~v_2434;
assign x_15500 = v_2889 | ~v_1180;
assign x_15501 = v_2889 | ~v_1181;
assign x_15502 = v_2889 | ~v_183;
assign x_15503 = v_2889 | ~v_167;
assign x_15504 = v_2889 | ~v_166;
assign x_15505 = v_2889 | ~v_159;
assign x_15506 = v_2889 | ~v_146;
assign x_15507 = v_2889 | ~v_145;
assign x_15508 = v_2889 | ~v_144;
assign x_15509 = v_2889 | ~v_143;
assign x_15510 = v_2889 | ~v_142;
assign x_15511 = v_2889 | ~v_61;
assign x_15512 = v_2889 | ~v_58;
assign x_15513 = v_2889 | ~v_51;
assign x_15514 = v_2888 | ~v_2832;
assign x_15515 = v_2888 | ~v_2833;
assign x_15516 = v_2888 | ~v_2834;
assign x_15517 = v_2888 | ~v_2835;
assign x_15518 = v_2888 | ~v_757;
assign x_15519 = v_2888 | ~v_758;
assign x_15520 = v_2888 | ~v_759;
assign x_15521 = v_2888 | ~v_760;
assign x_15522 = v_2888 | ~v_1157;
assign x_15523 = v_2888 | ~v_1158;
assign x_15524 = v_2888 | ~v_1159;
assign x_15525 = v_2888 | ~v_1160;
assign x_15526 = v_2888 | ~v_761;
assign x_15527 = v_2888 | ~v_764;
assign x_15528 = v_2888 | ~v_1161;
assign x_15529 = v_2888 | ~v_1162;
assign x_15530 = v_2888 | ~v_1163;
assign x_15531 = v_2888 | ~v_1164;
assign x_15532 = v_2888 | ~v_2454;
assign x_15533 = v_2888 | ~v_2455;
assign x_15534 = v_2888 | ~v_2456;
assign x_15535 = v_2888 | ~v_2457;
assign x_15536 = v_2888 | ~v_771;
assign x_15537 = v_2888 | ~v_772;
assign x_15538 = v_2888 | ~v_2486;
assign x_15539 = v_2888 | ~v_2487;
assign x_15540 = v_2888 | ~v_2488;
assign x_15541 = v_2888 | ~v_2489;
assign x_15542 = v_2888 | ~v_2416;
assign x_15543 = v_2888 | ~v_2419;
assign x_15544 = v_2888 | ~v_1165;
assign x_15545 = v_2888 | ~v_1166;
assign x_15546 = v_2888 | ~v_182;
assign x_15547 = v_2888 | ~v_163;
assign x_15548 = v_2888 | ~v_162;
assign x_15549 = v_2888 | ~v_155;
assign x_15550 = v_2888 | ~v_138;
assign x_15551 = v_2888 | ~v_137;
assign x_15552 = v_2888 | ~v_136;
assign x_15553 = v_2888 | ~v_135;
assign x_15554 = v_2888 | ~v_134;
assign x_15555 = v_2888 | ~v_18;
assign x_15556 = v_2888 | ~v_15;
assign x_15557 = v_2888 | ~v_8;
assign x_15558 = ~v_2886 | ~v_2885 | ~v_2884 | v_2887;
assign x_15559 = v_2886 | ~v_2842;
assign x_15560 = v_2886 | ~v_2843;
assign x_15561 = v_2886 | ~v_2844;
assign x_15562 = v_2886 | ~v_2845;
assign x_15563 = v_2886 | ~v_969;
assign x_15564 = v_2886 | ~v_970;
assign x_15565 = v_2886 | ~v_971;
assign x_15566 = v_2886 | ~v_972;
assign x_15567 = v_2886 | ~v_827;
assign x_15568 = v_2886 | ~v_828;
assign x_15569 = v_2886 | ~v_829;
assign x_15570 = v_2886 | ~v_830;
assign x_15571 = v_2886 | ~v_831;
assign x_15572 = v_2886 | ~v_832;
assign x_15573 = v_2886 | ~v_1147;
assign x_15574 = v_2886 | ~v_1148;
assign x_15575 = v_2886 | ~v_975;
assign x_15576 = v_2886 | ~v_976;
assign x_15577 = v_2886 | ~v_2442;
assign x_15578 = v_2886 | ~v_2443;
assign x_15579 = v_2886 | ~v_2444;
assign x_15580 = v_2886 | ~v_2445;
assign x_15581 = v_2886 | ~v_839;
assign x_15582 = v_2886 | ~v_840;
assign x_15583 = v_2886 | ~v_2446;
assign x_15584 = v_2886 | ~v_2447;
assign x_15585 = v_2886 | ~v_2448;
assign x_15586 = v_2886 | ~v_2449;
assign x_15587 = v_2886 | ~v_2450;
assign x_15588 = v_2886 | ~v_2451;
assign x_15589 = v_2886 | ~v_1149;
assign x_15590 = v_2886 | ~v_1150;
assign x_15591 = v_2886 | ~v_184;
assign x_15592 = v_2886 | ~v_170;
assign x_15593 = v_2886 | ~v_169;
assign x_15594 = v_2886 | ~v_150;
assign x_15595 = v_2886 | ~v_149;
assign x_15596 = v_2886 | ~v_147;
assign x_15597 = v_2886 | ~v_103;
assign x_15598 = v_2886 | ~v_102;
assign x_15599 = v_2886 | ~v_101;
assign x_15600 = v_2886 | ~v_100;
assign x_15601 = v_2886 | ~v_98;
assign x_15602 = v_2886 | ~v_96;
assign x_15603 = v_2885 | ~v_2837;
assign x_15604 = v_2885 | ~v_2838;
assign x_15605 = v_2885 | ~v_2839;
assign x_15606 = v_2885 | ~v_2840;
assign x_15607 = v_2885 | ~v_954;
assign x_15608 = v_2885 | ~v_955;
assign x_15609 = v_2885 | ~v_956;
assign x_15610 = v_2885 | ~v_957;
assign x_15611 = v_2885 | ~v_794;
assign x_15612 = v_2885 | ~v_795;
assign x_15613 = v_2885 | ~v_796;
assign x_15614 = v_2885 | ~v_797;
assign x_15615 = v_2885 | ~v_798;
assign x_15616 = v_2885 | ~v_799;
assign x_15617 = v_2885 | ~v_1142;
assign x_15618 = v_2885 | ~v_1143;
assign x_15619 = v_2885 | ~v_960;
assign x_15620 = v_2885 | ~v_961;
assign x_15621 = v_2885 | ~v_2427;
assign x_15622 = v_2885 | ~v_2428;
assign x_15623 = v_2885 | ~v_2429;
assign x_15624 = v_2885 | ~v_2430;
assign x_15625 = v_2885 | ~v_806;
assign x_15626 = v_2885 | ~v_2431;
assign x_15627 = v_2885 | ~v_2432;
assign x_15628 = v_2885 | ~v_2433;
assign x_15629 = v_2885 | ~v_2434;
assign x_15630 = v_2885 | ~v_2435;
assign x_15631 = v_2885 | ~v_2436;
assign x_15632 = v_2885 | ~v_807;
assign x_15633 = v_2885 | ~v_1144;
assign x_15634 = v_2885 | ~v_1145;
assign x_15635 = v_2885 | ~v_183;
assign x_15636 = v_2885 | ~v_166;
assign x_15637 = v_2885 | ~v_165;
assign x_15638 = v_2885 | ~v_145;
assign x_15639 = v_2885 | ~v_144;
assign x_15640 = v_2885 | ~v_142;
assign x_15641 = v_2885 | ~v_61;
assign x_15642 = v_2885 | ~v_60;
assign x_15643 = v_2885 | ~v_59;
assign x_15644 = v_2885 | ~v_58;
assign x_15645 = v_2885 | ~v_56;
assign x_15646 = v_2885 | ~v_54;
assign x_15647 = v_2884 | ~v_2832;
assign x_15648 = v_2884 | ~v_2833;
assign x_15649 = v_2884 | ~v_2834;
assign x_15650 = v_2884 | ~v_2835;
assign x_15651 = v_2884 | ~v_939;
assign x_15652 = v_2884 | ~v_940;
assign x_15653 = v_2884 | ~v_941;
assign x_15654 = v_2884 | ~v_942;
assign x_15655 = v_2884 | ~v_761;
assign x_15656 = v_2884 | ~v_762;
assign x_15657 = v_2884 | ~v_763;
assign x_15658 = v_2884 | ~v_764;
assign x_15659 = v_2884 | ~v_765;
assign x_15660 = v_2884 | ~v_766;
assign x_15661 = v_2884 | ~v_1137;
assign x_15662 = v_2884 | ~v_1138;
assign x_15663 = v_2884 | ~v_945;
assign x_15664 = v_2884 | ~v_946;
assign x_15665 = v_2884 | ~v_2412;
assign x_15666 = v_2884 | ~v_2413;
assign x_15667 = v_2884 | ~v_2414;
assign x_15668 = v_2884 | ~v_2415;
assign x_15669 = v_2884 | ~v_773;
assign x_15670 = v_2884 | ~v_774;
assign x_15671 = v_2884 | ~v_2416;
assign x_15672 = v_2884 | ~v_2417;
assign x_15673 = v_2884 | ~v_2418;
assign x_15674 = v_2884 | ~v_2419;
assign x_15675 = v_2884 | ~v_2420;
assign x_15676 = v_2884 | ~v_2421;
assign x_15677 = v_2884 | ~v_1139;
assign x_15678 = v_2884 | ~v_1140;
assign x_15679 = v_2884 | ~v_182;
assign x_15680 = v_2884 | ~v_162;
assign x_15681 = v_2884 | ~v_161;
assign x_15682 = v_2884 | ~v_137;
assign x_15683 = v_2884 | ~v_136;
assign x_15684 = v_2884 | ~v_134;
assign x_15685 = v_2884 | ~v_18;
assign x_15686 = v_2884 | ~v_17;
assign x_15687 = v_2884 | ~v_16;
assign x_15688 = v_2884 | ~v_15;
assign x_15689 = v_2884 | ~v_13;
assign x_15690 = v_2884 | ~v_11;
assign x_15691 = ~v_2882 | ~v_2881 | ~v_2880 | v_2883;
assign x_15692 = v_2882 | ~v_2842;
assign x_15693 = v_2882 | ~v_2843;
assign x_15694 = v_2882 | ~v_2844;
assign x_15695 = v_2882 | ~v_2845;
assign x_15696 = v_2882 | ~v_1077;
assign x_15697 = v_2882 | ~v_1078;
assign x_15698 = v_2882 | ~v_1079;
assign x_15699 = v_2882 | ~v_1080;
assign x_15700 = v_2882 | ~v_827;
assign x_15701 = v_2882 | ~v_1015;
assign x_15702 = v_2882 | ~v_1016;
assign x_15703 = v_2882 | ~v_830;
assign x_15704 = v_2882 | ~v_1017;
assign x_15705 = v_2882 | ~v_1018;
assign x_15706 = v_2882 | ~v_1085;
assign x_15707 = v_2882 | ~v_1131;
assign x_15708 = v_2882 | ~v_1132;
assign x_15709 = v_2882 | ~v_1086;
assign x_15710 = v_2882 | ~v_1133;
assign x_15711 = v_2882 | ~v_1134;
assign x_15712 = v_2882 | ~v_2532;
assign x_15713 = v_2882 | ~v_2533;
assign x_15714 = v_2882 | ~v_2534;
assign x_15715 = v_2882 | ~v_2535;
assign x_15716 = v_2882 | ~v_1023;
assign x_15717 = v_2882 | ~v_1024;
assign x_15718 = v_2882 | ~v_2446;
assign x_15719 = v_2882 | ~v_2512;
assign x_15720 = v_2882 | ~v_2513;
assign x_15721 = v_2882 | ~v_2449;
assign x_15722 = v_2882 | ~v_2514;
assign x_15723 = v_2882 | ~v_2515;
assign x_15724 = v_2882 | ~v_184;
assign x_15725 = v_2882 | ~v_172;
assign x_15726 = v_2882 | ~v_171;
assign x_15727 = v_2882 | ~v_169;
assign x_15728 = v_2882 | ~v_149;
assign x_15729 = v_2882 | ~v_148;
assign x_15730 = v_2882 | ~v_147;
assign x_15731 = v_2882 | ~v_102;
assign x_15732 = v_2882 | ~v_101;
assign x_15733 = v_2882 | ~v_100;
assign x_15734 = v_2882 | ~v_99;
assign x_15735 = v_2882 | ~v_94;
assign x_15736 = v_2881 | ~v_2837;
assign x_15737 = v_2881 | ~v_2838;
assign x_15738 = v_2881 | ~v_2839;
assign x_15739 = v_2881 | ~v_2840;
assign x_15740 = v_2881 | ~v_1062;
assign x_15741 = v_2881 | ~v_1063;
assign x_15742 = v_2881 | ~v_1064;
assign x_15743 = v_2881 | ~v_1065;
assign x_15744 = v_2881 | ~v_794;
assign x_15745 = v_2881 | ~v_1000;
assign x_15746 = v_2881 | ~v_1001;
assign x_15747 = v_2881 | ~v_797;
assign x_15748 = v_2881 | ~v_1002;
assign x_15749 = v_2881 | ~v_1003;
assign x_15750 = v_2881 | ~v_1070;
assign x_15751 = v_2881 | ~v_1126;
assign x_15752 = v_2881 | ~v_1127;
assign x_15753 = v_2881 | ~v_1071;
assign x_15754 = v_2881 | ~v_1128;
assign x_15755 = v_2881 | ~v_1129;
assign x_15756 = v_2881 | ~v_2527;
assign x_15757 = v_2881 | ~v_2528;
assign x_15758 = v_2881 | ~v_2529;
assign x_15759 = v_2881 | ~v_2530;
assign x_15760 = v_2881 | ~v_1008;
assign x_15761 = v_2881 | ~v_1009;
assign x_15762 = v_2881 | ~v_2431;
assign x_15763 = v_2881 | ~v_2507;
assign x_15764 = v_2881 | ~v_2508;
assign x_15765 = v_2881 | ~v_2434;
assign x_15766 = v_2881 | ~v_2509;
assign x_15767 = v_2881 | ~v_2510;
assign x_15768 = v_2881 | ~v_183;
assign x_15769 = v_2881 | ~v_168;
assign x_15770 = v_2881 | ~v_167;
assign x_15771 = v_2881 | ~v_165;
assign x_15772 = v_2881 | ~v_144;
assign x_15773 = v_2881 | ~v_143;
assign x_15774 = v_2881 | ~v_142;
assign x_15775 = v_2881 | ~v_60;
assign x_15776 = v_2881 | ~v_59;
assign x_15777 = v_2881 | ~v_58;
assign x_15778 = v_2881 | ~v_57;
assign x_15779 = v_2881 | ~v_52;
assign x_15780 = v_2880 | ~v_2832;
assign x_15781 = v_2880 | ~v_2833;
assign x_15782 = v_2880 | ~v_2834;
assign x_15783 = v_2880 | ~v_2835;
assign x_15784 = v_2880 | ~v_1047;
assign x_15785 = v_2880 | ~v_1048;
assign x_15786 = v_2880 | ~v_1049;
assign x_15787 = v_2880 | ~v_1050;
assign x_15788 = v_2880 | ~v_761;
assign x_15789 = v_2880 | ~v_985;
assign x_15790 = v_2880 | ~v_986;
assign x_15791 = v_2880 | ~v_764;
assign x_15792 = v_2880 | ~v_987;
assign x_15793 = v_2880 | ~v_988;
assign x_15794 = v_2880 | ~v_1055;
assign x_15795 = v_2880 | ~v_1121;
assign x_15796 = v_2880 | ~v_1122;
assign x_15797 = v_2880 | ~v_1056;
assign x_15798 = v_2880 | ~v_1123;
assign x_15799 = v_2880 | ~v_1124;
assign x_15800 = v_2880 | ~v_2522;
assign x_15801 = v_2880 | ~v_2523;
assign x_15802 = v_2880 | ~v_2524;
assign x_15803 = v_2880 | ~v_2525;
assign x_15804 = v_2880 | ~v_2416;
assign x_15805 = v_2880 | ~v_2502;
assign x_15806 = v_2880 | ~v_2503;
assign x_15807 = v_2880 | ~v_2419;
assign x_15808 = v_2880 | ~v_2504;
assign x_15809 = v_2880 | ~v_2505;
assign x_15810 = v_2880 | ~v_182;
assign x_15811 = v_2880 | ~v_164;
assign x_15812 = v_2880 | ~v_163;
assign x_15813 = v_2880 | ~v_161;
assign x_15814 = v_2880 | ~v_136;
assign x_15815 = v_2880 | ~v_135;
assign x_15816 = v_2880 | ~v_134;
assign x_15817 = v_2880 | ~v_993;
assign x_15818 = v_2880 | ~v_994;
assign x_15819 = v_2880 | ~v_17;
assign x_15820 = v_2880 | ~v_16;
assign x_15821 = v_2880 | ~v_15;
assign x_15822 = v_2880 | ~v_14;
assign x_15823 = v_2880 | ~v_9;
assign x_15824 = ~v_2878 | ~v_2877 | ~v_2876 | v_2879;
assign x_15825 = v_2878 | ~v_2842;
assign x_15826 = v_2878 | ~v_2843;
assign x_15827 = v_2878 | ~v_2844;
assign x_15828 = v_2878 | ~v_2845;
assign x_15829 = v_2878 | ~v_1077;
assign x_15830 = v_2878 | ~v_1078;
assign x_15831 = v_2878 | ~v_1079;
assign x_15832 = v_2878 | ~v_1080;
assign x_15833 = v_2878 | ~v_969;
assign x_15834 = v_2878 | ~v_970;
assign x_15835 = v_2878 | ~v_971;
assign x_15836 = v_2878 | ~v_972;
assign x_15837 = v_2878 | ~v_827;
assign x_15838 = v_2878 | ~v_830;
assign x_15839 = v_2878 | ~v_975;
assign x_15840 = v_2878 | ~v_976;
assign x_15841 = v_2878 | ~v_1115;
assign x_15842 = v_2878 | ~v_1116;
assign x_15843 = v_2878 | ~v_2442;
assign x_15844 = v_2878 | ~v_2443;
assign x_15845 = v_2878 | ~v_2444;
assign x_15846 = v_2878 | ~v_2445;
assign x_15847 = v_2878 | ~v_1085;
assign x_15848 = v_2878 | ~v_1086;
assign x_15849 = v_2878 | ~v_2532;
assign x_15850 = v_2878 | ~v_2533;
assign x_15851 = v_2878 | ~v_2534;
assign x_15852 = v_2878 | ~v_2535;
assign x_15853 = v_2878 | ~v_2446;
assign x_15854 = v_2878 | ~v_2449;
assign x_15855 = v_2878 | ~v_1117;
assign x_15856 = v_2878 | ~v_1118;
assign x_15857 = v_2878 | ~v_184;
assign x_15858 = v_2878 | ~v_171;
assign x_15859 = v_2878 | ~v_169;
assign x_15860 = v_2878 | ~v_151;
assign x_15861 = v_2878 | ~v_150;
assign x_15862 = v_2878 | ~v_149;
assign x_15863 = v_2878 | ~v_147;
assign x_15864 = v_2878 | ~v_103;
assign x_15865 = v_2878 | ~v_101;
assign x_15866 = v_2878 | ~v_100;
assign x_15867 = v_2878 | ~v_96;
assign x_15868 = v_2878 | ~v_94;
assign x_15869 = v_2877 | ~v_2837;
assign x_15870 = v_2877 | ~v_2838;
assign x_15871 = v_2877 | ~v_2839;
assign x_15872 = v_2877 | ~v_2840;
assign x_15873 = v_2877 | ~v_1062;
assign x_15874 = v_2877 | ~v_1063;
assign x_15875 = v_2877 | ~v_1064;
assign x_15876 = v_2877 | ~v_1065;
assign x_15877 = v_2877 | ~v_954;
assign x_15878 = v_2877 | ~v_955;
assign x_15879 = v_2877 | ~v_956;
assign x_15880 = v_2877 | ~v_957;
assign x_15881 = v_2877 | ~v_794;
assign x_15882 = v_2877 | ~v_797;
assign x_15883 = v_2877 | ~v_960;
assign x_15884 = v_2877 | ~v_961;
assign x_15885 = v_2877 | ~v_1110;
assign x_15886 = v_2877 | ~v_1111;
assign x_15887 = v_2877 | ~v_2427;
assign x_15888 = v_2877 | ~v_2428;
assign x_15889 = v_2877 | ~v_2429;
assign x_15890 = v_2877 | ~v_2430;
assign x_15891 = v_2877 | ~v_1070;
assign x_15892 = v_2877 | ~v_1071;
assign x_15893 = v_2877 | ~v_2527;
assign x_15894 = v_2877 | ~v_2528;
assign x_15895 = v_2877 | ~v_2529;
assign x_15896 = v_2877 | ~v_2530;
assign x_15897 = v_2877 | ~v_2431;
assign x_15898 = v_2877 | ~v_2434;
assign x_15899 = v_2877 | ~v_1112;
assign x_15900 = v_2877 | ~v_1113;
assign x_15901 = v_2877 | ~v_183;
assign x_15902 = v_2877 | ~v_167;
assign x_15903 = v_2877 | ~v_165;
assign x_15904 = v_2877 | ~v_146;
assign x_15905 = v_2877 | ~v_145;
assign x_15906 = v_2877 | ~v_144;
assign x_15907 = v_2877 | ~v_142;
assign x_15908 = v_2877 | ~v_61;
assign x_15909 = v_2877 | ~v_59;
assign x_15910 = v_2877 | ~v_58;
assign x_15911 = v_2877 | ~v_54;
assign x_15912 = v_2877 | ~v_52;
assign x_15913 = v_2876 | ~v_2832;
assign x_15914 = v_2876 | ~v_2833;
assign x_15915 = v_2876 | ~v_2834;
assign x_15916 = v_2876 | ~v_2835;
assign x_15917 = v_2876 | ~v_1047;
assign x_15918 = v_2876 | ~v_1048;
assign x_15919 = v_2876 | ~v_1049;
assign x_15920 = v_2876 | ~v_1050;
assign x_15921 = v_2876 | ~v_939;
assign x_15922 = v_2876 | ~v_940;
assign x_15923 = v_2876 | ~v_941;
assign x_15924 = v_2876 | ~v_942;
assign x_15925 = v_2876 | ~v_761;
assign x_15926 = v_2876 | ~v_764;
assign x_15927 = v_2876 | ~v_945;
assign x_15928 = v_2876 | ~v_946;
assign x_15929 = v_2876 | ~v_1105;
assign x_15930 = v_2876 | ~v_1106;
assign x_15931 = v_2876 | ~v_2412;
assign x_15932 = v_2876 | ~v_2413;
assign x_15933 = v_2876 | ~v_2414;
assign x_15934 = v_2876 | ~v_2415;
assign x_15935 = v_2876 | ~v_1055;
assign x_15936 = v_2876 | ~v_1056;
assign x_15937 = v_2876 | ~v_2522;
assign x_15938 = v_2876 | ~v_2523;
assign x_15939 = v_2876 | ~v_2524;
assign x_15940 = v_2876 | ~v_2525;
assign x_15941 = v_2876 | ~v_2416;
assign x_15942 = v_2876 | ~v_2419;
assign x_15943 = v_2876 | ~v_1107;
assign x_15944 = v_2876 | ~v_1108;
assign x_15945 = v_2876 | ~v_182;
assign x_15946 = v_2876 | ~v_163;
assign x_15947 = v_2876 | ~v_161;
assign x_15948 = v_2876 | ~v_138;
assign x_15949 = v_2876 | ~v_137;
assign x_15950 = v_2876 | ~v_136;
assign x_15951 = v_2876 | ~v_134;
assign x_15952 = v_2876 | ~v_18;
assign x_15953 = v_2876 | ~v_16;
assign x_15954 = v_2876 | ~v_15;
assign x_15955 = v_2876 | ~v_11;
assign x_15956 = v_2876 | ~v_9;
assign x_15957 = ~v_2874 | ~v_2873 | ~v_2872 | v_2875;
assign x_15958 = v_2874 | ~v_2842;
assign x_15959 = v_2874 | ~v_2843;
assign x_15960 = v_2874 | ~v_2844;
assign x_15961 = v_2874 | ~v_2845;
assign x_15962 = v_2874 | ~v_1077;
assign x_15963 = v_2874 | ~v_1078;
assign x_15964 = v_2874 | ~v_1079;
assign x_15965 = v_2874 | ~v_1080;
assign x_15966 = v_2874 | ~v_921;
assign x_15967 = v_2874 | ~v_922;
assign x_15968 = v_2874 | ~v_923;
assign x_15969 = v_2874 | ~v_924;
assign x_15970 = v_2874 | ~v_827;
assign x_15971 = v_2874 | ~v_830;
assign x_15972 = v_2874 | ~v_927;
assign x_15973 = v_2874 | ~v_928;
assign x_15974 = v_2874 | ~v_1099;
assign x_15975 = v_2874 | ~v_1100;
assign x_15976 = v_2874 | ~v_1101;
assign x_15977 = v_2874 | ~v_1102;
assign x_15978 = v_2874 | ~v_2480;
assign x_15979 = v_2874 | ~v_2481;
assign x_15980 = v_2874 | ~v_2482;
assign x_15981 = v_2874 | ~v_2483;
assign x_15982 = v_2874 | ~v_1085;
assign x_15983 = v_2874 | ~v_1086;
assign x_15984 = v_2874 | ~v_2532;
assign x_15985 = v_2874 | ~v_2533;
assign x_15986 = v_2874 | ~v_2534;
assign x_15987 = v_2874 | ~v_2535;
assign x_15988 = v_2874 | ~v_2446;
assign x_15989 = v_2874 | ~v_2449;
assign x_15990 = v_2874 | ~v_184;
assign x_15991 = v_2874 | ~v_171;
assign x_15992 = v_2874 | ~v_169;
assign x_15993 = v_2874 | ~v_150;
assign x_15994 = v_2874 | ~v_148;
assign x_15995 = v_2874 | ~v_103;
assign x_15996 = v_2874 | ~v_102;
assign x_15997 = v_2874 | ~v_101;
assign x_15998 = v_2874 | ~v_100;
assign x_15999 = v_2874 | ~v_97;
assign x_16000 = v_2874 | ~v_95;
assign x_16001 = v_2874 | ~v_94;
assign x_16002 = v_2873 | ~v_2837;
assign x_16003 = v_2873 | ~v_2838;
assign x_16004 = v_2873 | ~v_2839;
assign x_16005 = v_2873 | ~v_2840;
assign x_16006 = v_2873 | ~v_1062;
assign x_16007 = v_2873 | ~v_1063;
assign x_16008 = v_2873 | ~v_1064;
assign x_16009 = v_2873 | ~v_1065;
assign x_16010 = v_2873 | ~v_906;
assign x_16011 = v_2873 | ~v_907;
assign x_16012 = v_2873 | ~v_908;
assign x_16013 = v_2873 | ~v_909;
assign x_16014 = v_2873 | ~v_794;
assign x_16015 = v_2873 | ~v_797;
assign x_16016 = v_2873 | ~v_912;
assign x_16017 = v_2873 | ~v_913;
assign x_16018 = v_2873 | ~v_1094;
assign x_16019 = v_2873 | ~v_1095;
assign x_16020 = v_2873 | ~v_1096;
assign x_16021 = v_2873 | ~v_1097;
assign x_16022 = v_2873 | ~v_2475;
assign x_16023 = v_2873 | ~v_2476;
assign x_16024 = v_2873 | ~v_2477;
assign x_16025 = v_2873 | ~v_2478;
assign x_16026 = v_2873 | ~v_1070;
assign x_16027 = v_2873 | ~v_1071;
assign x_16028 = v_2873 | ~v_2527;
assign x_16029 = v_2873 | ~v_2528;
assign x_16030 = v_2873 | ~v_2529;
assign x_16031 = v_2873 | ~v_2530;
assign x_16032 = v_2873 | ~v_2431;
assign x_16033 = v_2873 | ~v_2434;
assign x_16034 = v_2873 | ~v_183;
assign x_16035 = v_2873 | ~v_167;
assign x_16036 = v_2873 | ~v_165;
assign x_16037 = v_2873 | ~v_145;
assign x_16038 = v_2873 | ~v_143;
assign x_16039 = v_2873 | ~v_61;
assign x_16040 = v_2873 | ~v_60;
assign x_16041 = v_2873 | ~v_59;
assign x_16042 = v_2873 | ~v_58;
assign x_16043 = v_2873 | ~v_55;
assign x_16044 = v_2873 | ~v_53;
assign x_16045 = v_2873 | ~v_52;
assign x_16046 = v_2872 | ~v_2832;
assign x_16047 = v_2872 | ~v_2833;
assign x_16048 = v_2872 | ~v_2834;
assign x_16049 = v_2872 | ~v_2835;
assign x_16050 = v_2872 | ~v_1047;
assign x_16051 = v_2872 | ~v_1048;
assign x_16052 = v_2872 | ~v_1049;
assign x_16053 = v_2872 | ~v_1050;
assign x_16054 = v_2872 | ~v_891;
assign x_16055 = v_2872 | ~v_892;
assign x_16056 = v_2872 | ~v_893;
assign x_16057 = v_2872 | ~v_894;
assign x_16058 = v_2872 | ~v_761;
assign x_16059 = v_2872 | ~v_764;
assign x_16060 = v_2872 | ~v_897;
assign x_16061 = v_2872 | ~v_898;
assign x_16062 = v_2872 | ~v_1089;
assign x_16063 = v_2872 | ~v_1090;
assign x_16064 = v_2872 | ~v_1091;
assign x_16065 = v_2872 | ~v_1092;
assign x_16066 = v_2872 | ~v_2470;
assign x_16067 = v_2872 | ~v_2471;
assign x_16068 = v_2872 | ~v_2472;
assign x_16069 = v_2872 | ~v_2473;
assign x_16070 = v_2872 | ~v_1055;
assign x_16071 = v_2872 | ~v_1056;
assign x_16072 = v_2872 | ~v_2522;
assign x_16073 = v_2872 | ~v_2523;
assign x_16074 = v_2872 | ~v_2524;
assign x_16075 = v_2872 | ~v_2525;
assign x_16076 = v_2872 | ~v_2416;
assign x_16077 = v_2872 | ~v_2419;
assign x_16078 = v_2872 | ~v_182;
assign x_16079 = v_2872 | ~v_163;
assign x_16080 = v_2872 | ~v_161;
assign x_16081 = v_2872 | ~v_137;
assign x_16082 = v_2872 | ~v_135;
assign x_16083 = v_2872 | ~v_18;
assign x_16084 = v_2872 | ~v_17;
assign x_16085 = v_2872 | ~v_16;
assign x_16086 = v_2872 | ~v_15;
assign x_16087 = v_2872 | ~v_12;
assign x_16088 = v_2872 | ~v_10;
assign x_16089 = v_2872 | ~v_9;
assign x_16090 = ~v_2870 | ~v_2869 | ~v_2868 | v_2871;
assign x_16091 = v_2870 | ~v_2842;
assign x_16092 = v_2870 | ~v_2843;
assign x_16093 = v_2870 | ~v_2844;
assign x_16094 = v_2870 | ~v_2845;
assign x_16095 = v_2870 | ~v_1077;
assign x_16096 = v_2870 | ~v_1078;
assign x_16097 = v_2870 | ~v_1079;
assign x_16098 = v_2870 | ~v_1080;
assign x_16099 = v_2870 | ~v_823;
assign x_16100 = v_2870 | ~v_824;
assign x_16101 = v_2870 | ~v_825;
assign x_16102 = v_2870 | ~v_826;
assign x_16103 = v_2870 | ~v_827;
assign x_16104 = v_2870 | ~v_830;
assign x_16105 = v_2870 | ~v_837;
assign x_16106 = v_2870 | ~v_838;
assign x_16107 = v_2870 | ~v_1081;
assign x_16108 = v_2870 | ~v_1082;
assign x_16109 = v_2870 | ~v_1083;
assign x_16110 = v_2870 | ~v_1084;
assign x_16111 = v_2870 | ~v_2496;
assign x_16112 = v_2870 | ~v_2497;
assign x_16113 = v_2870 | ~v_2498;
assign x_16114 = v_2870 | ~v_2499;
assign x_16115 = v_2870 | ~v_1085;
assign x_16116 = v_2870 | ~v_1086;
assign x_16117 = v_2870 | ~v_2532;
assign x_16118 = v_2870 | ~v_2533;
assign x_16119 = v_2870 | ~v_2534;
assign x_16120 = v_2870 | ~v_2535;
assign x_16121 = v_2870 | ~v_2446;
assign x_16122 = v_2870 | ~v_2449;
assign x_16123 = v_2870 | ~v_184;
assign x_16124 = v_2870 | ~v_171;
assign x_16125 = v_2870 | ~v_169;
assign x_16126 = v_2870 | ~v_160;
assign x_16127 = v_2870 | ~v_150;
assign x_16128 = v_2870 | ~v_149;
assign x_16129 = v_2870 | ~v_148;
assign x_16130 = v_2870 | ~v_147;
assign x_16131 = v_2870 | ~v_103;
assign x_16132 = v_2870 | ~v_102;
assign x_16133 = v_2870 | ~v_100;
assign x_16134 = v_2870 | ~v_94;
assign x_16135 = v_2869 | ~v_2837;
assign x_16136 = v_2869 | ~v_2838;
assign x_16137 = v_2869 | ~v_2839;
assign x_16138 = v_2869 | ~v_2840;
assign x_16139 = v_2869 | ~v_1062;
assign x_16140 = v_2869 | ~v_1063;
assign x_16141 = v_2869 | ~v_1064;
assign x_16142 = v_2869 | ~v_1065;
assign x_16143 = v_2869 | ~v_790;
assign x_16144 = v_2869 | ~v_791;
assign x_16145 = v_2869 | ~v_792;
assign x_16146 = v_2869 | ~v_793;
assign x_16147 = v_2869 | ~v_794;
assign x_16148 = v_2869 | ~v_797;
assign x_16149 = v_2869 | ~v_804;
assign x_16150 = v_2869 | ~v_805;
assign x_16151 = v_2869 | ~v_1066;
assign x_16152 = v_2869 | ~v_1067;
assign x_16153 = v_2869 | ~v_1068;
assign x_16154 = v_2869 | ~v_1069;
assign x_16155 = v_2869 | ~v_2491;
assign x_16156 = v_2869 | ~v_2492;
assign x_16157 = v_2869 | ~v_2493;
assign x_16158 = v_2869 | ~v_2494;
assign x_16159 = v_2869 | ~v_1070;
assign x_16160 = v_2869 | ~v_1071;
assign x_16161 = v_2869 | ~v_2527;
assign x_16162 = v_2869 | ~v_2528;
assign x_16163 = v_2869 | ~v_2529;
assign x_16164 = v_2869 | ~v_2530;
assign x_16165 = v_2869 | ~v_2431;
assign x_16166 = v_2869 | ~v_2434;
assign x_16167 = v_2869 | ~v_183;
assign x_16168 = v_2869 | ~v_167;
assign x_16169 = v_2869 | ~v_165;
assign x_16170 = v_2869 | ~v_159;
assign x_16171 = v_2869 | ~v_145;
assign x_16172 = v_2869 | ~v_144;
assign x_16173 = v_2869 | ~v_143;
assign x_16174 = v_2869 | ~v_142;
assign x_16175 = v_2869 | ~v_61;
assign x_16176 = v_2869 | ~v_60;
assign x_16177 = v_2869 | ~v_58;
assign x_16178 = v_2869 | ~v_52;
assign x_16179 = v_2868 | ~v_2832;
assign x_16180 = v_2868 | ~v_2833;
assign x_16181 = v_2868 | ~v_2834;
assign x_16182 = v_2868 | ~v_2835;
assign x_16183 = v_2868 | ~v_1047;
assign x_16184 = v_2868 | ~v_1048;
assign x_16185 = v_2868 | ~v_1049;
assign x_16186 = v_2868 | ~v_1050;
assign x_16187 = v_2868 | ~v_757;
assign x_16188 = v_2868 | ~v_758;
assign x_16189 = v_2868 | ~v_759;
assign x_16190 = v_2868 | ~v_760;
assign x_16191 = v_2868 | ~v_761;
assign x_16192 = v_2868 | ~v_764;
assign x_16193 = v_2868 | ~v_771;
assign x_16194 = v_2868 | ~v_772;
assign x_16195 = v_2868 | ~v_1051;
assign x_16196 = v_2868 | ~v_1052;
assign x_16197 = v_2868 | ~v_1053;
assign x_16198 = v_2868 | ~v_1054;
assign x_16199 = v_2868 | ~v_2486;
assign x_16200 = v_2868 | ~v_2487;
assign x_16201 = v_2868 | ~v_2488;
assign x_16202 = v_2868 | ~v_2489;
assign x_16203 = v_2868 | ~v_1055;
assign x_16204 = v_2868 | ~v_1056;
assign x_16205 = v_2868 | ~v_2522;
assign x_16206 = v_2868 | ~v_2523;
assign x_16207 = v_2868 | ~v_2524;
assign x_16208 = v_2868 | ~v_2525;
assign x_16209 = v_2868 | ~v_2416;
assign x_16210 = v_2868 | ~v_2419;
assign x_16211 = v_2868 | ~v_182;
assign x_16212 = v_2868 | ~v_163;
assign x_16213 = v_2868 | ~v_161;
assign x_16214 = v_2868 | ~v_155;
assign x_16215 = v_2868 | ~v_137;
assign x_16216 = v_2868 | ~v_136;
assign x_16217 = v_2868 | ~v_135;
assign x_16218 = v_2868 | ~v_134;
assign x_16219 = v_2868 | ~v_18;
assign x_16220 = v_2868 | ~v_17;
assign x_16221 = v_2868 | ~v_15;
assign x_16222 = v_2868 | ~v_9;
assign x_16223 = ~v_2866 | ~v_2865 | ~v_2864 | v_2867;
assign x_16224 = v_2866 | ~v_2842;
assign x_16225 = v_2866 | ~v_2843;
assign x_16226 = v_2866 | ~v_2844;
assign x_16227 = v_2866 | ~v_2845;
assign x_16228 = v_2866 | ~v_921;
assign x_16229 = v_2866 | ~v_922;
assign x_16230 = v_2866 | ~v_923;
assign x_16231 = v_2866 | ~v_924;
assign x_16232 = v_2866 | ~v_827;
assign x_16233 = v_2866 | ~v_828;
assign x_16234 = v_2866 | ~v_829;
assign x_16235 = v_2866 | ~v_830;
assign x_16236 = v_2866 | ~v_831;
assign x_16237 = v_2866 | ~v_832;
assign x_16238 = v_2866 | ~v_1037;
assign x_16239 = v_2866 | ~v_1038;
assign x_16240 = v_2866 | ~v_1039;
assign x_16241 = v_2866 | ~v_1040;
assign x_16242 = v_2866 | ~v_927;
assign x_16243 = v_2866 | ~v_928;
assign x_16244 = v_2866 | ~v_2480;
assign x_16245 = v_2866 | ~v_2481;
assign x_16246 = v_2866 | ~v_2482;
assign x_16247 = v_2866 | ~v_2483;
assign x_16248 = v_2866 | ~v_839;
assign x_16249 = v_2866 | ~v_840;
assign x_16250 = v_2866 | ~v_2446;
assign x_16251 = v_2866 | ~v_2447;
assign x_16252 = v_2866 | ~v_2448;
assign x_16253 = v_2866 | ~v_2449;
assign x_16254 = v_2866 | ~v_2450;
assign x_16255 = v_2866 | ~v_2451;
assign x_16256 = v_2866 | ~v_184;
assign x_16257 = v_2866 | ~v_170;
assign x_16258 = v_2866 | ~v_169;
assign x_16259 = v_2866 | ~v_151;
assign x_16260 = v_2866 | ~v_150;
assign x_16261 = v_2866 | ~v_148;
assign x_16262 = v_2866 | ~v_147;
assign x_16263 = v_2866 | ~v_103;
assign x_16264 = v_2866 | ~v_101;
assign x_16265 = v_2866 | ~v_100;
assign x_16266 = v_2866 | ~v_98;
assign x_16267 = v_2866 | ~v_97;
assign x_16268 = v_2865 | ~v_2837;
assign x_16269 = v_2865 | ~v_2838;
assign x_16270 = v_2865 | ~v_2839;
assign x_16271 = v_2865 | ~v_2840;
assign x_16272 = v_2865 | ~v_906;
assign x_16273 = v_2865 | ~v_907;
assign x_16274 = v_2865 | ~v_908;
assign x_16275 = v_2865 | ~v_909;
assign x_16276 = v_2865 | ~v_794;
assign x_16277 = v_2865 | ~v_795;
assign x_16278 = v_2865 | ~v_796;
assign x_16279 = v_2865 | ~v_797;
assign x_16280 = v_2865 | ~v_798;
assign x_16281 = v_2865 | ~v_799;
assign x_16282 = v_2865 | ~v_1032;
assign x_16283 = v_2865 | ~v_1033;
assign x_16284 = v_2865 | ~v_1034;
assign x_16285 = v_2865 | ~v_1035;
assign x_16286 = v_2865 | ~v_912;
assign x_16287 = v_2865 | ~v_913;
assign x_16288 = v_2865 | ~v_2475;
assign x_16289 = v_2865 | ~v_2476;
assign x_16290 = v_2865 | ~v_2477;
assign x_16291 = v_2865 | ~v_2478;
assign x_16292 = v_2865 | ~v_806;
assign x_16293 = v_2865 | ~v_2431;
assign x_16294 = v_2865 | ~v_2432;
assign x_16295 = v_2865 | ~v_2433;
assign x_16296 = v_2865 | ~v_2434;
assign x_16297 = v_2865 | ~v_2435;
assign x_16298 = v_2865 | ~v_2436;
assign x_16299 = v_2865 | ~v_807;
assign x_16300 = v_2865 | ~v_183;
assign x_16301 = v_2865 | ~v_166;
assign x_16302 = v_2865 | ~v_165;
assign x_16303 = v_2865 | ~v_146;
assign x_16304 = v_2865 | ~v_145;
assign x_16305 = v_2865 | ~v_143;
assign x_16306 = v_2865 | ~v_142;
assign x_16307 = v_2865 | ~v_61;
assign x_16308 = v_2865 | ~v_59;
assign x_16309 = v_2865 | ~v_58;
assign x_16310 = v_2865 | ~v_56;
assign x_16311 = v_2865 | ~v_55;
assign x_16312 = v_2864 | ~v_2832;
assign x_16313 = v_2864 | ~v_2833;
assign x_16314 = v_2864 | ~v_2834;
assign x_16315 = v_2864 | ~v_2835;
assign x_16316 = v_2864 | ~v_891;
assign x_16317 = v_2864 | ~v_892;
assign x_16318 = v_2864 | ~v_893;
assign x_16319 = v_2864 | ~v_894;
assign x_16320 = v_2864 | ~v_761;
assign x_16321 = v_2864 | ~v_762;
assign x_16322 = v_2864 | ~v_763;
assign x_16323 = v_2864 | ~v_764;
assign x_16324 = v_2864 | ~v_765;
assign x_16325 = v_2864 | ~v_766;
assign x_16326 = v_2864 | ~v_1027;
assign x_16327 = v_2864 | ~v_1028;
assign x_16328 = v_2864 | ~v_1029;
assign x_16329 = v_2864 | ~v_1030;
assign x_16330 = v_2864 | ~v_897;
assign x_16331 = v_2864 | ~v_898;
assign x_16332 = v_2864 | ~v_2470;
assign x_16333 = v_2864 | ~v_2471;
assign x_16334 = v_2864 | ~v_2472;
assign x_16335 = v_2864 | ~v_2473;
assign x_16336 = v_2864 | ~v_773;
assign x_16337 = v_2864 | ~v_774;
assign x_16338 = v_2864 | ~v_2416;
assign x_16339 = v_2864 | ~v_2417;
assign x_16340 = v_2864 | ~v_2418;
assign x_16341 = v_2864 | ~v_2419;
assign x_16342 = v_2864 | ~v_2420;
assign x_16343 = v_2864 | ~v_2421;
assign x_16344 = v_2864 | ~v_182;
assign x_16345 = v_2864 | ~v_162;
assign x_16346 = v_2864 | ~v_161;
assign x_16347 = v_2864 | ~v_138;
assign x_16348 = v_2864 | ~v_137;
assign x_16349 = v_2864 | ~v_135;
assign x_16350 = v_2864 | ~v_134;
assign x_16351 = v_2864 | ~v_18;
assign x_16352 = v_2864 | ~v_16;
assign x_16353 = v_2864 | ~v_15;
assign x_16354 = v_2864 | ~v_13;
assign x_16355 = v_2864 | ~v_12;
assign x_16356 = ~v_2862 | ~v_2861 | ~v_2860 | v_2863;
assign x_16357 = v_2862 | ~v_2842;
assign x_16358 = v_2862 | ~v_2843;
assign x_16359 = v_2862 | ~v_2844;
assign x_16360 = v_2862 | ~v_2845;
assign x_16361 = v_2862 | ~v_877;
assign x_16362 = v_2862 | ~v_878;
assign x_16363 = v_2862 | ~v_879;
assign x_16364 = v_2862 | ~v_880;
assign x_16365 = v_2862 | ~v_827;
assign x_16366 = v_2862 | ~v_1015;
assign x_16367 = v_2862 | ~v_1016;
assign x_16368 = v_2862 | ~v_830;
assign x_16369 = v_2862 | ~v_1017;
assign x_16370 = v_2862 | ~v_1018;
assign x_16371 = v_2862 | ~v_885;
assign x_16372 = v_2862 | ~v_1019;
assign x_16373 = v_2862 | ~v_1020;
assign x_16374 = v_2862 | ~v_886;
assign x_16375 = v_2862 | ~v_1021;
assign x_16376 = v_2862 | ~v_1022;
assign x_16377 = v_2862 | ~v_2564;
assign x_16378 = v_2862 | ~v_2565;
assign x_16379 = v_2862 | ~v_2566;
assign x_16380 = v_2862 | ~v_2567;
assign x_16381 = v_2862 | ~v_1023;
assign x_16382 = v_2862 | ~v_1024;
assign x_16383 = v_2862 | ~v_2446;
assign x_16384 = v_2862 | ~v_2512;
assign x_16385 = v_2862 | ~v_2513;
assign x_16386 = v_2862 | ~v_2449;
assign x_16387 = v_2862 | ~v_2514;
assign x_16388 = v_2862 | ~v_2515;
assign x_16389 = v_2862 | ~v_184;
assign x_16390 = v_2862 | ~v_181;
assign x_16391 = v_2862 | ~v_171;
assign x_16392 = v_2862 | ~v_170;
assign x_16393 = v_2862 | ~v_169;
assign x_16394 = v_2862 | ~v_149;
assign x_16395 = v_2862 | ~v_148;
assign x_16396 = v_2862 | ~v_147;
assign x_16397 = v_2862 | ~v_103;
assign x_16398 = v_2862 | ~v_102;
assign x_16399 = v_2862 | ~v_101;
assign x_16400 = v_2862 | ~v_99;
assign x_16401 = v_2861 | ~v_2837;
assign x_16402 = v_2861 | ~v_2838;
assign x_16403 = v_2861 | ~v_2839;
assign x_16404 = v_2861 | ~v_2840;
assign x_16405 = v_2861 | ~v_862;
assign x_16406 = v_2861 | ~v_863;
assign x_16407 = v_2861 | ~v_864;
assign x_16408 = v_2861 | ~v_865;
assign x_16409 = v_2861 | ~v_794;
assign x_16410 = v_2861 | ~v_1000;
assign x_16411 = v_2861 | ~v_1001;
assign x_16412 = v_2861 | ~v_797;
assign x_16413 = v_2861 | ~v_1002;
assign x_16414 = v_2861 | ~v_1003;
assign x_16415 = v_2861 | ~v_870;
assign x_16416 = v_2861 | ~v_1004;
assign x_16417 = v_2861 | ~v_1005;
assign x_16418 = v_2861 | ~v_871;
assign x_16419 = v_2861 | ~v_1006;
assign x_16420 = v_2861 | ~v_1007;
assign x_16421 = v_2861 | ~v_2559;
assign x_16422 = v_2861 | ~v_2560;
assign x_16423 = v_2861 | ~v_2561;
assign x_16424 = v_2861 | ~v_2562;
assign x_16425 = v_2861 | ~v_1008;
assign x_16426 = v_2861 | ~v_1009;
assign x_16427 = v_2861 | ~v_2431;
assign x_16428 = v_2861 | ~v_2507;
assign x_16429 = v_2861 | ~v_2508;
assign x_16430 = v_2861 | ~v_2434;
assign x_16431 = v_2861 | ~v_2509;
assign x_16432 = v_2861 | ~v_2510;
assign x_16433 = v_2861 | ~v_183;
assign x_16434 = v_2861 | ~v_180;
assign x_16435 = v_2861 | ~v_167;
assign x_16436 = v_2861 | ~v_166;
assign x_16437 = v_2861 | ~v_165;
assign x_16438 = v_2861 | ~v_144;
assign x_16439 = v_2861 | ~v_143;
assign x_16440 = v_2861 | ~v_142;
assign x_16441 = v_2861 | ~v_61;
assign x_16442 = v_2861 | ~v_60;
assign x_16443 = v_2861 | ~v_59;
assign x_16444 = v_2861 | ~v_57;
assign x_16445 = v_2860 | ~v_2832;
assign x_16446 = v_2860 | ~v_2833;
assign x_16447 = v_2860 | ~v_2834;
assign x_16448 = v_2860 | ~v_2835;
assign x_16449 = v_2860 | ~v_847;
assign x_16450 = v_2860 | ~v_848;
assign x_16451 = v_2860 | ~v_849;
assign x_16452 = v_2860 | ~v_850;
assign x_16453 = v_2860 | ~v_761;
assign x_16454 = v_2860 | ~v_985;
assign x_16455 = v_2860 | ~v_986;
assign x_16456 = v_2860 | ~v_764;
assign x_16457 = v_2860 | ~v_987;
assign x_16458 = v_2860 | ~v_988;
assign x_16459 = v_2860 | ~v_855;
assign x_16460 = v_2860 | ~v_989;
assign x_16461 = v_2860 | ~v_990;
assign x_16462 = v_2860 | ~v_856;
assign x_16463 = v_2860 | ~v_991;
assign x_16464 = v_2860 | ~v_992;
assign x_16465 = v_2860 | ~v_2554;
assign x_16466 = v_2860 | ~v_2555;
assign x_16467 = v_2860 | ~v_2556;
assign x_16468 = v_2860 | ~v_2557;
assign x_16469 = v_2860 | ~v_2416;
assign x_16470 = v_2860 | ~v_2502;
assign x_16471 = v_2860 | ~v_2503;
assign x_16472 = v_2860 | ~v_2419;
assign x_16473 = v_2860 | ~v_2504;
assign x_16474 = v_2860 | ~v_2505;
assign x_16475 = v_2860 | ~v_182;
assign x_16476 = v_2860 | ~v_179;
assign x_16477 = v_2860 | ~v_163;
assign x_16478 = v_2860 | ~v_162;
assign x_16479 = v_2860 | ~v_161;
assign x_16480 = v_2860 | ~v_136;
assign x_16481 = v_2860 | ~v_135;
assign x_16482 = v_2860 | ~v_134;
assign x_16483 = v_2860 | ~v_993;
assign x_16484 = v_2860 | ~v_994;
assign x_16485 = v_2860 | ~v_18;
assign x_16486 = v_2860 | ~v_17;
assign x_16487 = v_2860 | ~v_16;
assign x_16488 = v_2860 | ~v_14;
assign x_16489 = ~v_2858 | ~v_2857 | ~v_2856 | v_2859;
assign x_16490 = v_2858 | ~v_2842;
assign x_16491 = v_2858 | ~v_2843;
assign x_16492 = v_2858 | ~v_2844;
assign x_16493 = v_2858 | ~v_2845;
assign x_16494 = v_2858 | ~v_877;
assign x_16495 = v_2858 | ~v_878;
assign x_16496 = v_2858 | ~v_879;
assign x_16497 = v_2858 | ~v_880;
assign x_16498 = v_2858 | ~v_969;
assign x_16499 = v_2858 | ~v_970;
assign x_16500 = v_2858 | ~v_971;
assign x_16501 = v_2858 | ~v_972;
assign x_16502 = v_2858 | ~v_827;
assign x_16503 = v_2858 | ~v_830;
assign x_16504 = v_2858 | ~v_973;
assign x_16505 = v_2858 | ~v_974;
assign x_16506 = v_2858 | ~v_885;
assign x_16507 = v_2858 | ~v_886;
assign x_16508 = v_2858 | ~v_2564;
assign x_16509 = v_2858 | ~v_2565;
assign x_16510 = v_2858 | ~v_2566;
assign x_16511 = v_2858 | ~v_2567;
assign x_16512 = v_2858 | ~v_975;
assign x_16513 = v_2858 | ~v_976;
assign x_16514 = v_2858 | ~v_2442;
assign x_16515 = v_2858 | ~v_2443;
assign x_16516 = v_2858 | ~v_2444;
assign x_16517 = v_2858 | ~v_2445;
assign x_16518 = v_2858 | ~v_2446;
assign x_16519 = v_2858 | ~v_2449;
assign x_16520 = v_2858 | ~v_977;
assign x_16521 = v_2858 | ~v_978;
assign x_16522 = v_2858 | ~v_184;
assign x_16523 = v_2858 | ~v_181;
assign x_16524 = v_2858 | ~v_172;
assign x_16525 = v_2858 | ~v_171;
assign x_16526 = v_2858 | ~v_170;
assign x_16527 = v_2858 | ~v_169;
assign x_16528 = v_2858 | ~v_150;
assign x_16529 = v_2858 | ~v_149;
assign x_16530 = v_2858 | ~v_147;
assign x_16531 = v_2858 | ~v_102;
assign x_16532 = v_2858 | ~v_101;
assign x_16533 = v_2858 | ~v_96;
assign x_16534 = v_2857 | ~v_2837;
assign x_16535 = v_2857 | ~v_2838;
assign x_16536 = v_2857 | ~v_2839;
assign x_16537 = v_2857 | ~v_2840;
assign x_16538 = v_2857 | ~v_862;
assign x_16539 = v_2857 | ~v_863;
assign x_16540 = v_2857 | ~v_864;
assign x_16541 = v_2857 | ~v_865;
assign x_16542 = v_2857 | ~v_954;
assign x_16543 = v_2857 | ~v_955;
assign x_16544 = v_2857 | ~v_956;
assign x_16545 = v_2857 | ~v_957;
assign x_16546 = v_2857 | ~v_794;
assign x_16547 = v_2857 | ~v_797;
assign x_16548 = v_2857 | ~v_958;
assign x_16549 = v_2857 | ~v_959;
assign x_16550 = v_2857 | ~v_870;
assign x_16551 = v_2857 | ~v_871;
assign x_16552 = v_2857 | ~v_2559;
assign x_16553 = v_2857 | ~v_2560;
assign x_16554 = v_2857 | ~v_2561;
assign x_16555 = v_2857 | ~v_2562;
assign x_16556 = v_2857 | ~v_960;
assign x_16557 = v_2857 | ~v_961;
assign x_16558 = v_2857 | ~v_2427;
assign x_16559 = v_2857 | ~v_2428;
assign x_16560 = v_2857 | ~v_2429;
assign x_16561 = v_2857 | ~v_2430;
assign x_16562 = v_2857 | ~v_2431;
assign x_16563 = v_2857 | ~v_2434;
assign x_16564 = v_2857 | ~v_962;
assign x_16565 = v_2857 | ~v_963;
assign x_16566 = v_2857 | ~v_183;
assign x_16567 = v_2857 | ~v_180;
assign x_16568 = v_2857 | ~v_168;
assign x_16569 = v_2857 | ~v_167;
assign x_16570 = v_2857 | ~v_166;
assign x_16571 = v_2857 | ~v_165;
assign x_16572 = v_2857 | ~v_145;
assign x_16573 = v_2857 | ~v_144;
assign x_16574 = v_2857 | ~v_142;
assign x_16575 = v_2857 | ~v_60;
assign x_16576 = v_2857 | ~v_59;
assign x_16577 = v_2857 | ~v_54;
assign x_16578 = v_2856 | ~v_2832;
assign x_16579 = v_2856 | ~v_2833;
assign x_16580 = v_2856 | ~v_2834;
assign x_16581 = v_2856 | ~v_2835;
assign x_16582 = v_2856 | ~v_847;
assign x_16583 = v_2856 | ~v_848;
assign x_16584 = v_2856 | ~v_849;
assign x_16585 = v_2856 | ~v_850;
assign x_16586 = v_2856 | ~v_939;
assign x_16587 = v_2856 | ~v_940;
assign x_16588 = v_2856 | ~v_941;
assign x_16589 = v_2856 | ~v_942;
assign x_16590 = v_2856 | ~v_761;
assign x_16591 = v_2856 | ~v_764;
assign x_16592 = v_2856 | ~v_943;
assign x_16593 = v_2856 | ~v_944;
assign x_16594 = v_2856 | ~v_855;
assign x_16595 = v_2856 | ~v_856;
assign x_16596 = v_2856 | ~v_2554;
assign x_16597 = v_2856 | ~v_2555;
assign x_16598 = v_2856 | ~v_2556;
assign x_16599 = v_2856 | ~v_2557;
assign x_16600 = v_2856 | ~v_945;
assign x_16601 = v_2856 | ~v_946;
assign x_16602 = v_2856 | ~v_2412;
assign x_16603 = v_2856 | ~v_2413;
assign x_16604 = v_2856 | ~v_2414;
assign x_16605 = v_2856 | ~v_2415;
assign x_16606 = v_2856 | ~v_2416;
assign x_16607 = v_2856 | ~v_2419;
assign x_16608 = v_2856 | ~v_947;
assign x_16609 = v_2856 | ~v_948;
assign x_16610 = v_2856 | ~v_182;
assign x_16611 = v_2856 | ~v_179;
assign x_16612 = v_2856 | ~v_164;
assign x_16613 = v_2856 | ~v_163;
assign x_16614 = v_2856 | ~v_162;
assign x_16615 = v_2856 | ~v_161;
assign x_16616 = v_2856 | ~v_137;
assign x_16617 = v_2856 | ~v_136;
assign x_16618 = v_2856 | ~v_134;
assign x_16619 = v_2856 | ~v_17;
assign x_16620 = v_2856 | ~v_16;
assign x_16621 = v_2856 | ~v_11;
assign x_16622 = ~v_2854 | ~v_2853 | ~v_2852 | v_2855;
assign x_16623 = v_2854 | ~v_2842;
assign x_16624 = v_2854 | ~v_2843;
assign x_16625 = v_2854 | ~v_2844;
assign x_16626 = v_2854 | ~v_2845;
assign x_16627 = v_2854 | ~v_877;
assign x_16628 = v_2854 | ~v_878;
assign x_16629 = v_2854 | ~v_879;
assign x_16630 = v_2854 | ~v_880;
assign x_16631 = v_2854 | ~v_921;
assign x_16632 = v_2854 | ~v_922;
assign x_16633 = v_2854 | ~v_923;
assign x_16634 = v_2854 | ~v_924;
assign x_16635 = v_2854 | ~v_827;
assign x_16636 = v_2854 | ~v_830;
assign x_16637 = v_2854 | ~v_925;
assign x_16638 = v_2854 | ~v_926;
assign x_16639 = v_2854 | ~v_885;
assign x_16640 = v_2854 | ~v_886;
assign x_16641 = v_2854 | ~v_2564;
assign x_16642 = v_2854 | ~v_2565;
assign x_16643 = v_2854 | ~v_2566;
assign x_16644 = v_2854 | ~v_2567;
assign x_16645 = v_2854 | ~v_927;
assign x_16646 = v_2854 | ~v_928;
assign x_16647 = v_2854 | ~v_2480;
assign x_16648 = v_2854 | ~v_2481;
assign x_16649 = v_2854 | ~v_2482;
assign x_16650 = v_2854 | ~v_2483;
assign x_16651 = v_2854 | ~v_2446;
assign x_16652 = v_2854 | ~v_2449;
assign x_16653 = v_2854 | ~v_929;
assign x_16654 = v_2854 | ~v_930;
assign x_16655 = v_2854 | ~v_184;
assign x_16656 = v_2854 | ~v_181;
assign x_16657 = v_2854 | ~v_171;
assign x_16658 = v_2854 | ~v_170;
assign x_16659 = v_2854 | ~v_169;
assign x_16660 = v_2854 | ~v_150;
assign x_16661 = v_2854 | ~v_148;
assign x_16662 = v_2854 | ~v_147;
assign x_16663 = v_2854 | ~v_103;
assign x_16664 = v_2854 | ~v_102;
assign x_16665 = v_2854 | ~v_101;
assign x_16666 = v_2854 | ~v_97;
assign x_16667 = v_2853 | ~v_2837;
assign x_16668 = v_2853 | ~v_2838;
assign x_16669 = v_2853 | ~v_2839;
assign x_16670 = v_2853 | ~v_2840;
assign x_16671 = v_2853 | ~v_862;
assign x_16672 = v_2853 | ~v_863;
assign x_16673 = v_2853 | ~v_864;
assign x_16674 = v_2853 | ~v_865;
assign x_16675 = v_2853 | ~v_906;
assign x_16676 = v_2853 | ~v_907;
assign x_16677 = v_2853 | ~v_908;
assign x_16678 = v_2853 | ~v_909;
assign x_16679 = v_2853 | ~v_794;
assign x_16680 = v_2853 | ~v_797;
assign x_16681 = v_2853 | ~v_910;
assign x_16682 = v_2853 | ~v_911;
assign x_16683 = v_2853 | ~v_870;
assign x_16684 = v_2853 | ~v_871;
assign x_16685 = v_2853 | ~v_2559;
assign x_16686 = v_2853 | ~v_2560;
assign x_16687 = v_2853 | ~v_2561;
assign x_16688 = v_2853 | ~v_2562;
assign x_16689 = v_2853 | ~v_912;
assign x_16690 = v_2853 | ~v_913;
assign x_16691 = v_2853 | ~v_2475;
assign x_16692 = v_2853 | ~v_2476;
assign x_16693 = v_2853 | ~v_2477;
assign x_16694 = v_2853 | ~v_2478;
assign x_16695 = v_2853 | ~v_2431;
assign x_16696 = v_2853 | ~v_2434;
assign x_16697 = v_2853 | ~v_914;
assign x_16698 = v_2853 | ~v_915;
assign x_16699 = v_2853 | ~v_183;
assign x_16700 = v_2853 | ~v_180;
assign x_16701 = v_2853 | ~v_167;
assign x_16702 = v_2853 | ~v_166;
assign x_16703 = v_2853 | ~v_165;
assign x_16704 = v_2853 | ~v_145;
assign x_16705 = v_2853 | ~v_143;
assign x_16706 = v_2853 | ~v_142;
assign x_16707 = v_2853 | ~v_61;
assign x_16708 = v_2853 | ~v_60;
assign x_16709 = v_2853 | ~v_59;
assign x_16710 = v_2853 | ~v_55;
assign x_16711 = v_2852 | ~v_2832;
assign x_16712 = v_2852 | ~v_2833;
assign x_16713 = v_2852 | ~v_2834;
assign x_16714 = v_2852 | ~v_2835;
assign x_16715 = v_2852 | ~v_847;
assign x_16716 = v_2852 | ~v_848;
assign x_16717 = v_2852 | ~v_849;
assign x_16718 = v_2852 | ~v_850;
assign x_16719 = v_2852 | ~v_891;
assign x_16720 = v_2852 | ~v_892;
assign x_16721 = v_2852 | ~v_893;
assign x_16722 = v_2852 | ~v_894;
assign x_16723 = v_2852 | ~v_761;
assign x_16724 = v_2852 | ~v_764;
assign x_16725 = v_2852 | ~v_895;
assign x_16726 = v_2852 | ~v_896;
assign x_16727 = v_2852 | ~v_855;
assign x_16728 = v_2852 | ~v_856;
assign x_16729 = v_2852 | ~v_2554;
assign x_16730 = v_2852 | ~v_2555;
assign x_16731 = v_2852 | ~v_2556;
assign x_16732 = v_2852 | ~v_2557;
assign x_16733 = v_2852 | ~v_897;
assign x_16734 = v_2852 | ~v_898;
assign x_16735 = v_2852 | ~v_2470;
assign x_16736 = v_2852 | ~v_2471;
assign x_16737 = v_2852 | ~v_2472;
assign x_16738 = v_2852 | ~v_2473;
assign x_16739 = v_2852 | ~v_2416;
assign x_16740 = v_2852 | ~v_2419;
assign x_16741 = v_2852 | ~v_899;
assign x_16742 = v_2852 | ~v_900;
assign x_16743 = v_2852 | ~v_182;
assign x_16744 = v_2852 | ~v_179;
assign x_16745 = v_2852 | ~v_163;
assign x_16746 = v_2852 | ~v_162;
assign x_16747 = v_2852 | ~v_161;
assign x_16748 = v_2852 | ~v_137;
assign x_16749 = v_2852 | ~v_135;
assign x_16750 = v_2852 | ~v_134;
assign x_16751 = v_2852 | ~v_18;
assign x_16752 = v_2852 | ~v_17;
assign x_16753 = v_2852 | ~v_16;
assign x_16754 = v_2852 | ~v_12;
assign x_16755 = ~v_2850 | ~v_2849 | ~v_2848 | v_2851;
assign x_16756 = v_2850 | ~v_2842;
assign x_16757 = v_2850 | ~v_2843;
assign x_16758 = v_2850 | ~v_2844;
assign x_16759 = v_2850 | ~v_2845;
assign x_16760 = v_2850 | ~v_877;
assign x_16761 = v_2850 | ~v_878;
assign x_16762 = v_2850 | ~v_879;
assign x_16763 = v_2850 | ~v_880;
assign x_16764 = v_2850 | ~v_823;
assign x_16765 = v_2850 | ~v_824;
assign x_16766 = v_2850 | ~v_825;
assign x_16767 = v_2850 | ~v_826;
assign x_16768 = v_2850 | ~v_827;
assign x_16769 = v_2850 | ~v_830;
assign x_16770 = v_2850 | ~v_881;
assign x_16771 = v_2850 | ~v_882;
assign x_16772 = v_2850 | ~v_883;
assign x_16773 = v_2850 | ~v_884;
assign x_16774 = v_2850 | ~v_885;
assign x_16775 = v_2850 | ~v_886;
assign x_16776 = v_2850 | ~v_2564;
assign x_16777 = v_2850 | ~v_2565;
assign x_16778 = v_2850 | ~v_2566;
assign x_16779 = v_2850 | ~v_2567;
assign x_16780 = v_2850 | ~v_837;
assign x_16781 = v_2850 | ~v_838;
assign x_16782 = v_2850 | ~v_2496;
assign x_16783 = v_2850 | ~v_2497;
assign x_16784 = v_2850 | ~v_2498;
assign x_16785 = v_2850 | ~v_2499;
assign x_16786 = v_2850 | ~v_2446;
assign x_16787 = v_2850 | ~v_2449;
assign x_16788 = v_2850 | ~v_184;
assign x_16789 = v_2850 | ~v_181;
assign x_16790 = v_2850 | ~v_171;
assign x_16791 = v_2850 | ~v_170;
assign x_16792 = v_2850 | ~v_169;
assign x_16793 = v_2850 | ~v_160;
assign x_16794 = v_2850 | ~v_150;
assign x_16795 = v_2850 | ~v_149;
assign x_16796 = v_2850 | ~v_148;
assign x_16797 = v_2850 | ~v_103;
assign x_16798 = v_2850 | ~v_102;
assign x_16799 = v_2850 | ~v_95;
assign x_16800 = v_2849 | ~v_2837;
assign x_16801 = v_2849 | ~v_2838;
assign x_16802 = v_2849 | ~v_2839;
assign x_16803 = v_2849 | ~v_2840;
assign x_16804 = v_2849 | ~v_862;
assign x_16805 = v_2849 | ~v_863;
assign x_16806 = v_2849 | ~v_864;
assign x_16807 = v_2849 | ~v_865;
assign x_16808 = v_2849 | ~v_790;
assign x_16809 = v_2849 | ~v_791;
assign x_16810 = v_2849 | ~v_792;
assign x_16811 = v_2849 | ~v_793;
assign x_16812 = v_2849 | ~v_794;
assign x_16813 = v_2849 | ~v_797;
assign x_16814 = v_2849 | ~v_866;
assign x_16815 = v_2849 | ~v_867;
assign x_16816 = v_2849 | ~v_868;
assign x_16817 = v_2849 | ~v_869;
assign x_16818 = v_2849 | ~v_870;
assign x_16819 = v_2849 | ~v_871;
assign x_16820 = v_2849 | ~v_2559;
assign x_16821 = v_2849 | ~v_2560;
assign x_16822 = v_2849 | ~v_2561;
assign x_16823 = v_2849 | ~v_2562;
assign x_16824 = v_2849 | ~v_804;
assign x_16825 = v_2849 | ~v_805;
assign x_16826 = v_2849 | ~v_2491;
assign x_16827 = v_2849 | ~v_2492;
assign x_16828 = v_2849 | ~v_2493;
assign x_16829 = v_2849 | ~v_2494;
assign x_16830 = v_2849 | ~v_2431;
assign x_16831 = v_2849 | ~v_2434;
assign x_16832 = v_2849 | ~v_183;
assign x_16833 = v_2849 | ~v_180;
assign x_16834 = v_2849 | ~v_167;
assign x_16835 = v_2849 | ~v_166;
assign x_16836 = v_2849 | ~v_165;
assign x_16837 = v_2849 | ~v_159;
assign x_16838 = v_2849 | ~v_145;
assign x_16839 = v_2849 | ~v_144;
assign x_16840 = v_2849 | ~v_143;
assign x_16841 = v_2849 | ~v_61;
assign x_16842 = v_2849 | ~v_60;
assign x_16843 = v_2849 | ~v_53;
assign x_16844 = v_2848 | ~v_2832;
assign x_16845 = v_2848 | ~v_2833;
assign x_16846 = v_2848 | ~v_2834;
assign x_16847 = v_2848 | ~v_2835;
assign x_16848 = v_2848 | ~v_847;
assign x_16849 = v_2848 | ~v_848;
assign x_16850 = v_2848 | ~v_849;
assign x_16851 = v_2848 | ~v_850;
assign x_16852 = v_2848 | ~v_757;
assign x_16853 = v_2848 | ~v_758;
assign x_16854 = v_2848 | ~v_759;
assign x_16855 = v_2848 | ~v_760;
assign x_16856 = v_2848 | ~v_761;
assign x_16857 = v_2848 | ~v_764;
assign x_16858 = v_2848 | ~v_851;
assign x_16859 = v_2848 | ~v_852;
assign x_16860 = v_2848 | ~v_853;
assign x_16861 = v_2848 | ~v_854;
assign x_16862 = v_2848 | ~v_855;
assign x_16863 = v_2848 | ~v_856;
assign x_16864 = v_2848 | ~v_2554;
assign x_16865 = v_2848 | ~v_2555;
assign x_16866 = v_2848 | ~v_2556;
assign x_16867 = v_2848 | ~v_2557;
assign x_16868 = v_2848 | ~v_771;
assign x_16869 = v_2848 | ~v_772;
assign x_16870 = v_2848 | ~v_2486;
assign x_16871 = v_2848 | ~v_2487;
assign x_16872 = v_2848 | ~v_2488;
assign x_16873 = v_2848 | ~v_2489;
assign x_16874 = v_2848 | ~v_2416;
assign x_16875 = v_2848 | ~v_2419;
assign x_16876 = v_2848 | ~v_182;
assign x_16877 = v_2848 | ~v_179;
assign x_16878 = v_2848 | ~v_163;
assign x_16879 = v_2848 | ~v_162;
assign x_16880 = v_2848 | ~v_161;
assign x_16881 = v_2848 | ~v_155;
assign x_16882 = v_2848 | ~v_137;
assign x_16883 = v_2848 | ~v_136;
assign x_16884 = v_2848 | ~v_135;
assign x_16885 = v_2848 | ~v_18;
assign x_16886 = v_2848 | ~v_17;
assign x_16887 = v_2848 | ~v_10;
assign x_16888 = ~v_2846 | ~v_2841 | ~v_2836 | v_2847;
assign x_16889 = v_2846 | ~v_2842;
assign x_16890 = v_2846 | ~v_2843;
assign x_16891 = v_2846 | ~v_2844;
assign x_16892 = v_2846 | ~v_2845;
assign x_16893 = v_2846 | ~v_823;
assign x_16894 = v_2846 | ~v_824;
assign x_16895 = v_2846 | ~v_825;
assign x_16896 = v_2846 | ~v_826;
assign x_16897 = v_2846 | ~v_827;
assign x_16898 = v_2846 | ~v_828;
assign x_16899 = v_2846 | ~v_829;
assign x_16900 = v_2846 | ~v_830;
assign x_16901 = v_2846 | ~v_831;
assign x_16902 = v_2846 | ~v_832;
assign x_16903 = v_2846 | ~v_833;
assign x_16904 = v_2846 | ~v_834;
assign x_16905 = v_2846 | ~v_835;
assign x_16906 = v_2846 | ~v_836;
assign x_16907 = v_2846 | ~v_837;
assign x_16908 = v_2846 | ~v_838;
assign x_16909 = v_2846 | ~v_2496;
assign x_16910 = v_2846 | ~v_2497;
assign x_16911 = v_2846 | ~v_2498;
assign x_16912 = v_2846 | ~v_2499;
assign x_16913 = v_2846 | ~v_839;
assign x_16914 = v_2846 | ~v_840;
assign x_16915 = v_2846 | ~v_2446;
assign x_16916 = v_2846 | ~v_2447;
assign x_16917 = v_2846 | ~v_2448;
assign x_16918 = v_2846 | ~v_2449;
assign x_16919 = v_2846 | ~v_2450;
assign x_16920 = v_2846 | ~v_2451;
assign x_16921 = v_2846 | ~v_184;
assign x_16922 = v_2846 | ~v_170;
assign x_16923 = v_2846 | ~v_169;
assign x_16924 = v_2846 | ~v_160;
assign x_16925 = v_2846 | ~v_150;
assign x_16926 = v_2846 | ~v_149;
assign x_16927 = v_2846 | ~v_148;
assign x_16928 = v_2846 | ~v_147;
assign x_16929 = v_2846 | ~v_103;
assign x_16930 = v_2846 | ~v_102;
assign x_16931 = v_2846 | ~v_100;
assign x_16932 = v_2846 | ~v_98;
assign x_16933 = ~v_123 | ~v_173 | v_2845;
assign x_16934 = ~v_120 | ~v_174 | v_2844;
assign x_16935 = ~v_108 | v_173 | v_2843;
assign x_16936 = ~v_105 | v_174 | v_2842;
assign x_16937 = v_2841 | ~v_2837;
assign x_16938 = v_2841 | ~v_2838;
assign x_16939 = v_2841 | ~v_2839;
assign x_16940 = v_2841 | ~v_2840;
assign x_16941 = v_2841 | ~v_790;
assign x_16942 = v_2841 | ~v_791;
assign x_16943 = v_2841 | ~v_792;
assign x_16944 = v_2841 | ~v_793;
assign x_16945 = v_2841 | ~v_794;
assign x_16946 = v_2841 | ~v_795;
assign x_16947 = v_2841 | ~v_796;
assign x_16948 = v_2841 | ~v_797;
assign x_16949 = v_2841 | ~v_798;
assign x_16950 = v_2841 | ~v_799;
assign x_16951 = v_2841 | ~v_800;
assign x_16952 = v_2841 | ~v_801;
assign x_16953 = v_2841 | ~v_802;
assign x_16954 = v_2841 | ~v_803;
assign x_16955 = v_2841 | ~v_804;
assign x_16956 = v_2841 | ~v_805;
assign x_16957 = v_2841 | ~v_2491;
assign x_16958 = v_2841 | ~v_2492;
assign x_16959 = v_2841 | ~v_2493;
assign x_16960 = v_2841 | ~v_2494;
assign x_16961 = v_2841 | ~v_806;
assign x_16962 = v_2841 | ~v_2431;
assign x_16963 = v_2841 | ~v_2432;
assign x_16964 = v_2841 | ~v_2433;
assign x_16965 = v_2841 | ~v_2434;
assign x_16966 = v_2841 | ~v_2435;
assign x_16967 = v_2841 | ~v_2436;
assign x_16968 = v_2841 | ~v_807;
assign x_16969 = v_2841 | ~v_183;
assign x_16970 = v_2841 | ~v_166;
assign x_16971 = v_2841 | ~v_165;
assign x_16972 = v_2841 | ~v_159;
assign x_16973 = v_2841 | ~v_145;
assign x_16974 = v_2841 | ~v_144;
assign x_16975 = v_2841 | ~v_143;
assign x_16976 = v_2841 | ~v_142;
assign x_16977 = v_2841 | ~v_61;
assign x_16978 = v_2841 | ~v_60;
assign x_16979 = v_2841 | ~v_58;
assign x_16980 = v_2841 | ~v_56;
assign x_16981 = ~v_81 | ~v_173 | v_2840;
assign x_16982 = ~v_78 | ~v_174 | v_2839;
assign x_16983 = ~v_66 | v_173 | v_2838;
assign x_16984 = ~v_63 | v_174 | v_2837;
assign x_16985 = v_2836 | ~v_2832;
assign x_16986 = v_2836 | ~v_2833;
assign x_16987 = v_2836 | ~v_2834;
assign x_16988 = v_2836 | ~v_2835;
assign x_16989 = v_2836 | ~v_757;
assign x_16990 = v_2836 | ~v_758;
assign x_16991 = v_2836 | ~v_759;
assign x_16992 = v_2836 | ~v_760;
assign x_16993 = v_2836 | ~v_761;
assign x_16994 = v_2836 | ~v_762;
assign x_16995 = v_2836 | ~v_763;
assign x_16996 = v_2836 | ~v_764;
assign x_16997 = v_2836 | ~v_765;
assign x_16998 = v_2836 | ~v_766;
assign x_16999 = v_2836 | ~v_767;
assign x_17000 = v_2836 | ~v_768;
assign x_17001 = v_2836 | ~v_769;
assign x_17002 = v_2836 | ~v_770;
assign x_17003 = v_2836 | ~v_771;
assign x_17004 = v_2836 | ~v_772;
assign x_17005 = v_2836 | ~v_2486;
assign x_17006 = v_2836 | ~v_2487;
assign x_17007 = v_2836 | ~v_2488;
assign x_17008 = v_2836 | ~v_2489;
assign x_17009 = v_2836 | ~v_773;
assign x_17010 = v_2836 | ~v_774;
assign x_17011 = v_2836 | ~v_2416;
assign x_17012 = v_2836 | ~v_2417;
assign x_17013 = v_2836 | ~v_2418;
assign x_17014 = v_2836 | ~v_2419;
assign x_17015 = v_2836 | ~v_2420;
assign x_17016 = v_2836 | ~v_2421;
assign x_17017 = v_2836 | ~v_182;
assign x_17018 = v_2836 | ~v_162;
assign x_17019 = v_2836 | ~v_161;
assign x_17020 = v_2836 | ~v_155;
assign x_17021 = v_2836 | ~v_137;
assign x_17022 = v_2836 | ~v_136;
assign x_17023 = v_2836 | ~v_135;
assign x_17024 = v_2836 | ~v_134;
assign x_17025 = v_2836 | ~v_18;
assign x_17026 = v_2836 | ~v_17;
assign x_17027 = v_2836 | ~v_15;
assign x_17028 = v_2836 | ~v_13;
assign x_17029 = ~v_39 | ~v_173 | v_2835;
assign x_17030 = ~v_36 | ~v_174 | v_2834;
assign x_17031 = ~v_24 | v_173 | v_2833;
assign x_17032 = ~v_21 | v_174 | v_2832;
assign x_17033 = v_2831 | ~v_2406;
assign x_17034 = v_2831 | ~v_737;
assign x_17035 = v_2830 | ~v_733;
assign x_17036 = v_2830 | ~v_730;
assign x_17037 = ~v_725 | ~v_724 | ~v_723 | ~v_722 | ~v_2828 | ~v_2824 | ~v_2820 | ~v_2816 | ~v_2812 | ~v_2808 | ~v_2804 | ~v_2800 | ~v_2796 | ~v_2792 | ~v_2788 | ~v_2784 | ~v_2780 | ~v_2776 | ~v_2772 | ~v_2768 | ~v_2752 | v_2829;
assign x_17038 = v_2828 | ~v_2825;
assign x_17039 = v_2828 | ~v_2826;
assign x_17040 = v_2828 | ~v_2827;
assign x_17041 = v_98 | v_103 | v_101 | v_100 | v_95 | v_99 | v_102 | ~v_719 | ~v_718 | v_170 | v_169 | v_149 | v_148 | v_184 | ~v_2331 | ~v_2267 | ~v_2330 | ~v_2266 | ~v_2265 | ~v_2329 | ~v_2264 | ~v_2328 | ~v_2263 | ~v_2262 | ~v_483 | ~v_717 | ~v_299 | ~v_482 | ~v_716 | ~v_298 | ~v_477 | ~v_291 | ~v_476 | ~v_290 | ~v_289 | ~v_475 | ~v_288 | ~v_474 | ~v_287 | ~v_286 | ~v_2766 | ~v_2765 | ~v_2764 | ~v_2763 | v_2827;
assign x_17042 = v_53 | v_56 | v_61 | v_60 | v_59 | v_58 | v_57 | ~v_714 | ~v_713 | v_144 | v_143 | v_166 | v_165 | v_183 | ~v_266 | ~v_2326 | ~v_2252 | ~v_2325 | ~v_2251 | ~v_2250 | ~v_2324 | ~v_2249 | ~v_2323 | ~v_2248 | ~v_2247 | ~v_468 | ~v_712 | ~v_467 | ~v_711 | ~v_265 | ~v_462 | ~v_258 | ~v_461 | ~v_257 | ~v_256 | ~v_460 | ~v_255 | ~v_459 | ~v_254 | ~v_253 | ~v_2761 | ~v_2760 | ~v_2759 | ~v_2758 | v_2826;
assign x_17043 = v_13 | v_18 | v_17 | v_16 | v_15 | v_14 | v_10 | ~v_453 | ~v_709 | ~v_452 | ~v_708 | v_136 | v_135 | ~v_707 | ~v_706 | v_162 | v_161 | v_182 | ~v_2321 | ~v_2237 | ~v_2320 | ~v_2236 | ~v_2235 | ~v_2319 | ~v_2234 | ~v_2318 | ~v_2233 | ~v_2232 | ~v_233 | ~v_232 | ~v_447 | ~v_225 | ~v_446 | ~v_224 | ~v_223 | ~v_445 | ~v_222 | ~v_444 | ~v_221 | ~v_220 | ~v_2756 | ~v_2755 | ~v_2754 | ~v_2753 | v_2825;
assign x_17044 = v_2824 | ~v_2821;
assign x_17045 = v_2824 | ~v_2822;
assign x_17046 = v_2824 | ~v_2823;
assign x_17047 = v_103 | v_101 | v_100 | v_99 | v_93 | v_102 | v_171 | v_170 | v_149 | v_148 | v_147 | v_184 | ~v_703 | ~v_702 | ~v_2331 | ~v_2330 | ~v_2265 | ~v_2329 | ~v_2328 | ~v_2262 | ~v_483 | ~v_482 | ~v_2283 | ~v_2282 | ~v_2281 | ~v_2280 | ~v_701 | ~v_653 | ~v_700 | ~v_652 | ~v_477 | ~v_476 | ~v_289 | ~v_475 | ~v_474 | ~v_286 | ~v_649 | ~v_648 | ~v_647 | ~v_646 | ~v_2766 | ~v_2765 | ~v_2764 | ~v_2763 | v_2823;
assign x_17048 = v_61 | v_51 | v_60 | v_59 | v_58 | v_57 | v_144 | v_143 | v_142 | v_167 | v_166 | v_183 | ~v_698 | ~v_697 | ~v_2326 | ~v_2325 | ~v_2250 | ~v_2324 | ~v_2323 | ~v_2247 | ~v_468 | ~v_467 | ~v_2278 | ~v_2277 | ~v_2276 | ~v_2275 | ~v_696 | ~v_638 | ~v_695 | ~v_637 | ~v_462 | ~v_461 | ~v_256 | ~v_460 | ~v_459 | ~v_253 | ~v_634 | ~v_633 | ~v_632 | ~v_631 | ~v_2761 | ~v_2760 | ~v_2759 | ~v_2758 | v_2822;
assign x_17049 = v_18 | v_17 | v_16 | v_8 | v_15 | v_14 | ~v_453 | ~v_452 | v_136 | v_135 | v_134 | v_163 | v_162 | v_182 | ~v_693 | ~v_692 | ~v_2321 | ~v_2320 | ~v_2235 | ~v_2319 | ~v_2318 | ~v_2232 | ~v_2273 | ~v_2272 | ~v_2271 | ~v_2270 | ~v_691 | ~v_623 | ~v_690 | ~v_622 | ~v_447 | ~v_446 | ~v_223 | ~v_445 | ~v_444 | ~v_220 | ~v_619 | ~v_618 | ~v_617 | ~v_616 | ~v_2756 | ~v_2755 | ~v_2754 | ~v_2753 | v_2821;
assign x_17050 = v_2820 | ~v_2817;
assign x_17051 = v_2820 | ~v_2818;
assign x_17052 = v_2820 | ~v_2819;
assign x_17053 = v_103 | v_101 | v_96 | v_100 | v_95 | v_93 | v_102 | v_171 | v_170 | v_150 | v_149 | v_184 | ~v_2265 | ~v_2262 | ~v_2261 | ~v_2260 | ~v_2259 | ~v_2258 | ~v_435 | ~v_434 | ~v_2283 | ~v_2282 | ~v_2281 | ~v_2280 | ~v_653 | ~v_652 | ~v_687 | ~v_686 | ~v_685 | ~v_684 | ~v_289 | ~v_286 | ~v_649 | ~v_648 | ~v_647 | ~v_646 | ~v_431 | ~v_430 | ~v_429 | ~v_428 | ~v_2766 | ~v_2765 | ~v_2764 | ~v_2763 | v_2819;
assign x_17054 = v_54 | v_53 | v_61 | v_51 | v_60 | v_59 | v_58 | v_144 | v_145 | v_167 | v_166 | v_183 | ~v_2250 | ~v_2247 | ~v_2246 | ~v_2245 | ~v_2244 | ~v_2243 | ~v_420 | ~v_419 | ~v_2278 | ~v_2277 | ~v_2276 | ~v_2275 | ~v_638 | ~v_637 | ~v_682 | ~v_681 | ~v_680 | ~v_679 | ~v_256 | ~v_253 | ~v_634 | ~v_633 | ~v_632 | ~v_631 | ~v_416 | ~v_415 | ~v_414 | ~v_413 | ~v_2761 | ~v_2760 | ~v_2759 | ~v_2758 | v_2818;
assign x_17055 = v_18 | v_17 | v_16 | v_8 | v_15 | v_11 | v_10 | v_136 | v_137 | v_163 | v_162 | v_182 | ~v_2235 | ~v_2232 | ~v_2231 | ~v_2230 | ~v_2229 | ~v_2228 | ~v_405 | ~v_404 | ~v_2273 | ~v_2272 | ~v_2271 | ~v_2270 | ~v_623 | ~v_622 | ~v_677 | ~v_676 | ~v_675 | ~v_674 | ~v_223 | ~v_220 | ~v_619 | ~v_618 | ~v_617 | ~v_616 | ~v_401 | ~v_400 | ~v_399 | ~v_398 | ~v_2756 | ~v_2755 | ~v_2754 | ~v_2753 | v_2817;
assign x_17056 = v_2816 | ~v_2813;
assign x_17057 = v_2816 | ~v_2814;
assign x_17058 = v_2816 | ~v_2815;
assign x_17059 = v_101 | v_97 | v_100 | v_93 | v_102 | v_172 | v_171 | v_170 | v_150 | v_148 | v_147 | v_184 | ~v_671 | ~v_670 | ~v_2265 | ~v_2262 | ~v_2299 | ~v_2298 | ~v_2297 | ~v_2296 | ~v_387 | ~v_386 | ~v_2283 | ~v_2282 | ~v_2281 | ~v_2280 | ~v_653 | ~v_652 | ~v_669 | ~v_668 | ~v_289 | ~v_286 | ~v_649 | ~v_648 | ~v_647 | ~v_646 | ~v_383 | ~v_382 | ~v_381 | ~v_380 | ~v_2766 | ~v_2765 | ~v_2764 | ~v_2763 | v_2815;
assign x_17060 = v_55 | v_51 | v_60 | v_59 | v_58 | v_145 | v_143 | v_142 | v_168 | v_167 | v_166 | v_183 | ~v_666 | ~v_665 | ~v_2250 | ~v_2247 | ~v_2294 | ~v_2293 | ~v_2292 | ~v_2291 | ~v_372 | ~v_371 | ~v_2278 | ~v_2277 | ~v_2276 | ~v_2275 | ~v_638 | ~v_637 | ~v_664 | ~v_663 | ~v_256 | ~v_253 | ~v_634 | ~v_633 | ~v_632 | ~v_631 | ~v_368 | ~v_367 | ~v_366 | ~v_365 | ~v_2761 | ~v_2760 | ~v_2759 | ~v_2758 | v_2814;
assign x_17061 = v_17 | v_16 | v_8 | v_15 | v_12 | v_135 | v_134 | v_137 | v_164 | v_163 | v_162 | v_182 | ~v_661 | ~v_660 | ~v_2235 | ~v_2232 | ~v_2289 | ~v_2288 | ~v_2287 | ~v_2286 | ~v_357 | ~v_356 | ~v_2273 | ~v_2272 | ~v_2271 | ~v_2270 | ~v_623 | ~v_622 | ~v_659 | ~v_658 | ~v_223 | ~v_220 | ~v_619 | ~v_618 | ~v_617 | ~v_616 | ~v_353 | ~v_352 | ~v_351 | ~v_350 | ~v_2756 | ~v_2755 | ~v_2754 | ~v_2753 | v_2813;
assign x_17062 = v_2812 | ~v_2809;
assign x_17063 = v_2812 | ~v_2810;
assign x_17064 = v_2812 | ~v_2811;
assign x_17065 = v_103 | v_100 | v_93 | v_151 | v_171 | v_170 | v_160 | v_150 | v_149 | v_148 | v_147 | v_184 | ~v_655 | ~v_654 | ~v_2265 | ~v_2262 | ~v_2315 | ~v_2314 | ~v_2313 | ~v_2312 | ~v_297 | ~v_296 | ~v_2283 | ~v_2282 | ~v_2281 | ~v_2280 | ~v_653 | ~v_652 | ~v_651 | ~v_650 | ~v_289 | ~v_286 | ~v_649 | ~v_648 | ~v_647 | ~v_646 | ~v_285 | ~v_284 | ~v_283 | ~v_282 | ~v_2766 | ~v_2765 | ~v_2764 | ~v_2763 | v_2811;
assign x_17066 = v_61 | v_51 | v_58 | v_144 | v_159 | v_145 | v_143 | v_142 | v_167 | v_166 | v_146 | v_183 | ~v_640 | ~v_639 | ~v_2250 | ~v_2247 | ~v_2310 | ~v_2309 | ~v_2308 | ~v_2307 | ~v_264 | ~v_263 | ~v_2278 | ~v_2277 | ~v_2276 | ~v_2275 | ~v_638 | ~v_637 | ~v_636 | ~v_635 | ~v_256 | ~v_253 | ~v_634 | ~v_633 | ~v_632 | ~v_631 | ~v_252 | ~v_251 | ~v_250 | ~v_249 | ~v_2761 | ~v_2760 | ~v_2759 | ~v_2758 | v_2810;
assign x_17067 = v_18 | v_8 | v_15 | v_136 | v_135 | v_134 | v_137 | v_138 | v_163 | v_162 | v_155 | v_182 | ~v_625 | ~v_624 | ~v_2235 | ~v_2232 | ~v_2305 | ~v_2304 | ~v_2303 | ~v_2302 | ~v_231 | ~v_230 | ~v_2273 | ~v_2272 | ~v_2271 | ~v_2270 | ~v_623 | ~v_622 | ~v_621 | ~v_620 | ~v_223 | ~v_220 | ~v_619 | ~v_618 | ~v_617 | ~v_616 | ~v_219 | ~v_218 | ~v_217 | ~v_216 | ~v_2756 | ~v_2755 | ~v_2754 | ~v_2753 | v_2809;
assign x_17068 = v_2808 | ~v_2805;
assign x_17069 = v_2808 | ~v_2806;
assign x_17070 = v_2808 | ~v_2807;
assign x_17071 = v_98 | v_103 | v_101 | v_96 | v_100 | v_102 | v_170 | v_169 | v_150 | v_149 | v_147 | v_184 | ~v_609 | ~v_608 | ~v_2267 | ~v_2266 | ~v_2265 | ~v_2264 | ~v_2263 | ~v_2262 | ~v_299 | ~v_298 | ~v_2261 | ~v_2260 | ~v_2259 | ~v_2258 | ~v_435 | ~v_434 | ~v_607 | ~v_606 | ~v_291 | ~v_290 | ~v_289 | ~v_288 | ~v_287 | ~v_286 | ~v_431 | ~v_430 | ~v_429 | ~v_428 | ~v_2766 | ~v_2765 | ~v_2764 | ~v_2763 | v_2807;
assign x_17072 = v_54 | v_56 | v_61 | v_60 | v_59 | v_58 | v_144 | v_145 | v_142 | v_166 | v_165 | v_183 | ~v_604 | ~v_603 | ~v_266 | ~v_2252 | ~v_2251 | ~v_2250 | ~v_2249 | ~v_2248 | ~v_2247 | ~v_265 | ~v_2246 | ~v_2245 | ~v_2244 | ~v_2243 | ~v_420 | ~v_419 | ~v_602 | ~v_601 | ~v_258 | ~v_257 | ~v_256 | ~v_255 | ~v_254 | ~v_253 | ~v_416 | ~v_415 | ~v_414 | ~v_413 | ~v_2761 | ~v_2760 | ~v_2759 | ~v_2758 | v_2806;
assign x_17073 = v_13 | v_18 | v_17 | v_16 | v_15 | v_11 | v_136 | v_134 | v_137 | v_162 | v_161 | v_182 | ~v_599 | ~v_598 | ~v_2237 | ~v_2236 | ~v_2235 | ~v_2234 | ~v_2233 | ~v_2232 | ~v_233 | ~v_232 | ~v_2231 | ~v_2230 | ~v_2229 | ~v_2228 | ~v_405 | ~v_404 | ~v_597 | ~v_596 | ~v_225 | ~v_224 | ~v_223 | ~v_222 | ~v_221 | ~v_220 | ~v_401 | ~v_400 | ~v_399 | ~v_398 | ~v_2756 | ~v_2755 | ~v_2754 | ~v_2753 | v_2805;
assign x_17074 = v_2804 | ~v_2801;
assign x_17075 = v_2804 | ~v_2802;
assign x_17076 = v_2804 | ~v_2803;
assign x_17077 = v_101 | v_100 | v_94 | v_99 | v_102 | v_172 | v_171 | v_169 | v_149 | v_148 | v_147 | v_184 | ~v_2331 | ~v_2330 | ~v_2265 | ~v_2329 | ~v_2328 | ~v_2262 | ~v_483 | ~v_482 | ~v_2351 | ~v_2350 | ~v_2349 | ~v_2348 | ~v_593 | ~v_592 | ~v_545 | ~v_591 | ~v_590 | ~v_544 | ~v_477 | ~v_476 | ~v_289 | ~v_475 | ~v_474 | ~v_286 | ~v_539 | ~v_538 | ~v_537 | ~v_536 | ~v_2766 | ~v_2765 | ~v_2764 | ~v_2763 | v_2803;
assign x_17078 = v_52 | v_60 | v_59 | v_58 | v_57 | v_144 | v_143 | v_142 | v_168 | v_167 | v_165 | v_183 | ~v_2326 | ~v_2325 | ~v_2250 | ~v_2324 | ~v_2323 | ~v_2247 | ~v_468 | ~v_467 | ~v_2346 | ~v_2345 | ~v_2344 | ~v_2343 | ~v_588 | ~v_587 | ~v_530 | ~v_586 | ~v_585 | ~v_529 | ~v_462 | ~v_461 | ~v_256 | ~v_460 | ~v_459 | ~v_253 | ~v_524 | ~v_523 | ~v_522 | ~v_521 | ~v_2761 | ~v_2760 | ~v_2759 | ~v_2758 | v_2802;
assign x_17079 = v_9 | v_17 | v_16 | v_15 | v_14 | ~v_453 | ~v_452 | v_136 | v_135 | v_134 | v_164 | v_163 | v_161 | v_182 | ~v_2321 | ~v_2320 | ~v_2235 | ~v_2319 | ~v_2318 | ~v_2232 | ~v_2341 | ~v_2340 | ~v_2339 | ~v_2338 | ~v_583 | ~v_582 | ~v_515 | ~v_581 | ~v_580 | ~v_514 | ~v_447 | ~v_446 | ~v_223 | ~v_445 | ~v_444 | ~v_220 | ~v_509 | ~v_508 | ~v_507 | ~v_506 | ~v_2756 | ~v_2755 | ~v_2754 | ~v_2753 | v_2801;
assign x_17080 = v_2800 | ~v_2797;
assign x_17081 = v_2800 | ~v_2798;
assign x_17082 = v_2800 | ~v_2799;
assign x_17083 = v_103 | v_101 | v_96 | v_100 | v_94 | v_151 | v_171 | v_169 | v_150 | v_149 | v_147 | v_184 | ~v_577 | ~v_576 | ~v_2265 | ~v_2262 | ~v_2351 | ~v_2350 | ~v_2349 | ~v_2348 | ~v_545 | ~v_544 | ~v_2261 | ~v_2260 | ~v_2259 | ~v_2258 | ~v_575 | ~v_574 | ~v_435 | ~v_434 | ~v_289 | ~v_286 | ~v_431 | ~v_430 | ~v_429 | ~v_428 | ~v_539 | ~v_538 | ~v_537 | ~v_536 | ~v_2766 | ~v_2765 | ~v_2764 | ~v_2763 | v_2799;
assign x_17084 = v_54 | v_61 | v_52 | v_59 | v_58 | v_144 | v_145 | v_142 | v_167 | v_165 | v_146 | v_183 | ~v_572 | ~v_571 | ~v_2250 | ~v_2247 | ~v_2346 | ~v_2345 | ~v_2344 | ~v_2343 | ~v_530 | ~v_529 | ~v_2246 | ~v_2245 | ~v_2244 | ~v_2243 | ~v_570 | ~v_569 | ~v_420 | ~v_419 | ~v_256 | ~v_253 | ~v_416 | ~v_415 | ~v_414 | ~v_413 | ~v_524 | ~v_523 | ~v_522 | ~v_521 | ~v_2761 | ~v_2760 | ~v_2759 | ~v_2758 | v_2798;
assign x_17085 = v_9 | v_18 | v_16 | v_15 | v_11 | v_136 | v_134 | v_137 | v_138 | v_163 | v_161 | v_182 | ~v_567 | ~v_566 | ~v_2235 | ~v_2232 | ~v_2341 | ~v_2340 | ~v_2339 | ~v_2338 | ~v_515 | ~v_514 | ~v_2231 | ~v_2230 | ~v_2229 | ~v_2228 | ~v_565 | ~v_564 | ~v_405 | ~v_404 | ~v_223 | ~v_220 | ~v_401 | ~v_400 | ~v_399 | ~v_398 | ~v_509 | ~v_508 | ~v_507 | ~v_506 | ~v_2756 | ~v_2755 | ~v_2754 | ~v_2753 | v_2797;
assign x_17086 = v_2796 | ~v_2793;
assign x_17087 = v_2796 | ~v_2794;
assign x_17088 = v_2796 | ~v_2795;
assign x_17089 = v_103 | v_101 | v_97 | v_100 | v_95 | v_94 | v_102 | v_171 | v_169 | v_150 | v_148 | v_184 | ~v_2265 | ~v_2262 | ~v_2351 | ~v_2350 | ~v_2349 | ~v_2348 | ~v_545 | ~v_544 | ~v_2299 | ~v_2298 | ~v_2297 | ~v_2296 | ~v_561 | ~v_560 | ~v_559 | ~v_558 | ~v_387 | ~v_386 | ~v_289 | ~v_286 | ~v_383 | ~v_382 | ~v_381 | ~v_380 | ~v_539 | ~v_538 | ~v_537 | ~v_536 | ~v_2766 | ~v_2765 | ~v_2764 | ~v_2763 | v_2795;
assign x_17090 = v_53 | v_55 | v_61 | v_52 | v_60 | v_59 | v_58 | v_145 | v_143 | v_167 | v_165 | v_183 | ~v_2250 | ~v_2247 | ~v_2346 | ~v_2345 | ~v_2344 | ~v_2343 | ~v_530 | ~v_529 | ~v_2294 | ~v_2293 | ~v_2292 | ~v_2291 | ~v_556 | ~v_555 | ~v_554 | ~v_553 | ~v_372 | ~v_371 | ~v_256 | ~v_253 | ~v_368 | ~v_367 | ~v_366 | ~v_365 | ~v_524 | ~v_523 | ~v_522 | ~v_521 | ~v_2761 | ~v_2760 | ~v_2759 | ~v_2758 | v_2794;
assign x_17091 = v_9 | v_18 | v_17 | v_16 | v_15 | v_12 | v_10 | v_135 | v_137 | v_163 | v_161 | v_182 | ~v_2235 | ~v_2232 | ~v_2341 | ~v_2340 | ~v_2339 | ~v_2338 | ~v_515 | ~v_514 | ~v_2289 | ~v_2288 | ~v_2287 | ~v_2286 | ~v_551 | ~v_550 | ~v_549 | ~v_548 | ~v_357 | ~v_356 | ~v_223 | ~v_220 | ~v_353 | ~v_352 | ~v_351 | ~v_350 | ~v_509 | ~v_508 | ~v_507 | ~v_506 | ~v_2756 | ~v_2755 | ~v_2754 | ~v_2753 | v_2793;
assign x_17092 = v_2792 | ~v_2789;
assign x_17093 = v_2792 | ~v_2790;
assign x_17094 = v_2792 | ~v_2791;
assign x_17095 = v_103 | v_100 | v_94 | v_102 | v_171 | v_169 | v_160 | v_150 | v_149 | v_148 | v_147 | v_184 | ~v_2265 | ~v_2262 | ~v_2351 | ~v_2350 | ~v_2349 | ~v_2348 | ~v_545 | ~v_544 | ~v_2315 | ~v_2314 | ~v_2313 | ~v_2312 | ~v_543 | ~v_542 | ~v_541 | ~v_540 | ~v_297 | ~v_296 | ~v_289 | ~v_286 | ~v_285 | ~v_284 | ~v_283 | ~v_282 | ~v_539 | ~v_538 | ~v_537 | ~v_536 | ~v_2766 | ~v_2765 | ~v_2764 | ~v_2763 | v_2791;
assign x_17096 = v_61 | v_52 | v_60 | v_58 | v_144 | v_159 | v_145 | v_143 | v_142 | v_167 | v_165 | v_183 | ~v_2250 | ~v_2247 | ~v_2346 | ~v_2345 | ~v_2344 | ~v_2343 | ~v_530 | ~v_529 | ~v_2310 | ~v_2309 | ~v_2308 | ~v_2307 | ~v_528 | ~v_527 | ~v_526 | ~v_525 | ~v_264 | ~v_263 | ~v_256 | ~v_253 | ~v_252 | ~v_251 | ~v_250 | ~v_249 | ~v_524 | ~v_523 | ~v_522 | ~v_521 | ~v_2761 | ~v_2760 | ~v_2759 | ~v_2758 | v_2790;
assign x_17097 = v_9 | v_18 | v_17 | v_15 | v_136 | v_135 | v_134 | v_137 | v_163 | v_161 | v_155 | v_182 | ~v_2235 | ~v_2232 | ~v_2341 | ~v_2340 | ~v_2339 | ~v_2338 | ~v_515 | ~v_514 | ~v_2305 | ~v_2304 | ~v_2303 | ~v_2302 | ~v_513 | ~v_512 | ~v_511 | ~v_510 | ~v_231 | ~v_230 | ~v_223 | ~v_220 | ~v_219 | ~v_218 | ~v_217 | ~v_216 | ~v_509 | ~v_508 | ~v_507 | ~v_506 | ~v_2756 | ~v_2755 | ~v_2754 | ~v_2753 | v_2789;
assign x_17098 = v_2788 | ~v_2785;
assign x_17099 = v_2788 | ~v_2786;
assign x_17100 = v_2788 | ~v_2787;
assign x_17101 = v_98 | v_103 | v_101 | v_97 | v_100 | v_151 | v_170 | v_169 | v_150 | v_148 | v_147 | v_184 | ~v_2267 | ~v_2266 | ~v_2265 | ~v_2264 | ~v_2263 | ~v_2262 | ~v_299 | ~v_298 | ~v_2299 | ~v_2298 | ~v_2297 | ~v_2296 | ~v_387 | ~v_386 | ~v_499 | ~v_498 | ~v_497 | ~v_496 | ~v_291 | ~v_290 | ~v_289 | ~v_288 | ~v_287 | ~v_286 | ~v_383 | ~v_382 | ~v_381 | ~v_380 | ~v_2766 | ~v_2765 | ~v_2764 | ~v_2763 | v_2787;
assign x_17102 = v_56 | v_55 | v_61 | v_59 | v_58 | v_145 | v_143 | v_142 | v_166 | v_165 | v_146 | v_183 | ~v_266 | ~v_2252 | ~v_2251 | ~v_2250 | ~v_2249 | ~v_2248 | ~v_2247 | ~v_265 | ~v_2294 | ~v_2293 | ~v_2292 | ~v_2291 | ~v_372 | ~v_371 | ~v_494 | ~v_493 | ~v_492 | ~v_491 | ~v_258 | ~v_257 | ~v_256 | ~v_255 | ~v_254 | ~v_253 | ~v_368 | ~v_367 | ~v_366 | ~v_365 | ~v_2761 | ~v_2760 | ~v_2759 | ~v_2758 | v_2786;
assign x_17103 = v_13 | v_18 | v_16 | v_15 | v_12 | v_135 | v_134 | v_137 | v_138 | v_162 | v_161 | v_182 | ~v_2237 | ~v_2236 | ~v_2235 | ~v_2234 | ~v_2233 | ~v_2232 | ~v_233 | ~v_232 | ~v_2289 | ~v_2288 | ~v_2287 | ~v_2286 | ~v_357 | ~v_356 | ~v_489 | ~v_488 | ~v_487 | ~v_486 | ~v_225 | ~v_224 | ~v_223 | ~v_222 | ~v_221 | ~v_220 | ~v_353 | ~v_352 | ~v_351 | ~v_350 | ~v_2756 | ~v_2755 | ~v_2754 | ~v_2753 | v_2785;
assign x_17104 = v_2784 | ~v_2781;
assign x_17105 = v_2784 | ~v_2782;
assign x_17106 = v_2784 | ~v_2783;
assign x_17107 = v_103 | v_101 | v_99 | v_102 | v_171 | v_170 | v_169 | v_149 | v_148 | v_147 | v_184 | v_181 | ~v_2331 | ~v_2330 | ~v_2265 | ~v_2329 | ~v_2328 | ~v_2262 | ~v_483 | ~v_482 | ~v_2383 | ~v_2382 | ~v_2381 | ~v_2380 | ~v_481 | ~v_480 | ~v_345 | ~v_479 | ~v_478 | ~v_344 | ~v_477 | ~v_476 | ~v_289 | ~v_475 | ~v_474 | ~v_286 | ~v_339 | ~v_338 | ~v_337 | ~v_336 | ~v_2766 | ~v_2765 | ~v_2764 | ~v_2763 | v_2783;
assign x_17108 = v_61 | v_60 | v_59 | v_57 | v_144 | v_180 | v_143 | v_142 | v_167 | v_166 | v_165 | v_183 | ~v_2326 | ~v_2325 | ~v_2250 | ~v_2324 | ~v_2323 | ~v_2247 | ~v_468 | ~v_467 | ~v_2378 | ~v_2377 | ~v_2376 | ~v_2375 | ~v_466 | ~v_465 | ~v_330 | ~v_464 | ~v_463 | ~v_329 | ~v_462 | ~v_461 | ~v_256 | ~v_460 | ~v_459 | ~v_253 | ~v_324 | ~v_323 | ~v_322 | ~v_321 | ~v_2761 | ~v_2760 | ~v_2759 | ~v_2758 | v_2782;
assign x_17109 = v_18 | v_17 | v_16 | v_14 | ~v_453 | ~v_452 | v_136 | v_135 | v_134 | v_179 | v_163 | v_162 | v_161 | v_182 | ~v_2321 | ~v_2320 | ~v_2235 | ~v_2319 | ~v_2318 | ~v_2232 | ~v_2373 | ~v_2372 | ~v_2371 | ~v_2370 | ~v_451 | ~v_450 | ~v_315 | ~v_449 | ~v_448 | ~v_314 | ~v_447 | ~v_446 | ~v_223 | ~v_445 | ~v_444 | ~v_220 | ~v_309 | ~v_308 | ~v_307 | ~v_306 | ~v_2756 | ~v_2755 | ~v_2754 | ~v_2753 | v_2781;
assign x_17110 = v_2780 | ~v_2777;
assign x_17111 = v_2780 | ~v_2778;
assign x_17112 = v_2780 | ~v_2779;
assign x_17113 = v_101 | v_96 | v_102 | v_172 | v_171 | v_170 | v_169 | v_150 | v_149 | v_147 | v_184 | v_181 | ~v_437 | ~v_436 | ~v_2265 | ~v_2262 | ~v_2261 | ~v_2260 | ~v_2259 | ~v_2258 | ~v_435 | ~v_434 | ~v_2383 | ~v_2382 | ~v_2381 | ~v_2380 | ~v_345 | ~v_344 | ~v_433 | ~v_432 | ~v_289 | ~v_286 | ~v_431 | ~v_430 | ~v_429 | ~v_428 | ~v_339 | ~v_338 | ~v_337 | ~v_336 | ~v_2766 | ~v_2765 | ~v_2764 | ~v_2763 | v_2779;
assign x_17114 = v_54 | v_60 | v_59 | v_144 | v_180 | v_145 | v_142 | v_168 | v_167 | v_166 | v_165 | v_183 | ~v_422 | ~v_421 | ~v_2250 | ~v_2247 | ~v_2246 | ~v_2245 | ~v_2244 | ~v_2243 | ~v_420 | ~v_419 | ~v_2378 | ~v_2377 | ~v_2376 | ~v_2375 | ~v_330 | ~v_329 | ~v_418 | ~v_417 | ~v_256 | ~v_253 | ~v_416 | ~v_415 | ~v_414 | ~v_413 | ~v_324 | ~v_323 | ~v_322 | ~v_321 | ~v_2761 | ~v_2760 | ~v_2759 | ~v_2758 | v_2778;
assign x_17115 = v_17 | v_16 | v_11 | v_136 | v_134 | v_137 | v_179 | v_164 | v_163 | v_162 | v_161 | v_182 | ~v_407 | ~v_406 | ~v_2235 | ~v_2232 | ~v_2231 | ~v_2230 | ~v_2229 | ~v_2228 | ~v_405 | ~v_404 | ~v_2373 | ~v_2372 | ~v_2371 | ~v_2370 | ~v_315 | ~v_314 | ~v_403 | ~v_402 | ~v_223 | ~v_220 | ~v_401 | ~v_400 | ~v_399 | ~v_398 | ~v_309 | ~v_308 | ~v_307 | ~v_306 | ~v_2756 | ~v_2755 | ~v_2754 | ~v_2753 | v_2777;
assign x_17116 = v_2776 | ~v_2773;
assign x_17117 = v_2776 | ~v_2774;
assign x_17118 = v_2776 | ~v_2775;
assign x_17119 = v_103 | v_101 | v_97 | v_102 | v_171 | v_170 | v_169 | v_150 | v_148 | v_147 | v_184 | v_181 | ~v_391 | ~v_390 | ~v_2265 | ~v_2262 | ~v_2299 | ~v_2298 | ~v_2297 | ~v_2296 | ~v_387 | ~v_386 | ~v_2383 | ~v_2382 | ~v_2381 | ~v_2380 | ~v_345 | ~v_344 | ~v_385 | ~v_384 | ~v_289 | ~v_286 | ~v_383 | ~v_382 | ~v_381 | ~v_380 | ~v_339 | ~v_338 | ~v_337 | ~v_336 | ~v_2766 | ~v_2765 | ~v_2764 | ~v_2763 | v_2775;
assign x_17120 = v_55 | v_61 | v_60 | v_59 | v_180 | v_145 | v_143 | v_142 | v_167 | v_166 | v_165 | v_183 | ~v_376 | ~v_375 | ~v_2250 | ~v_2247 | ~v_2294 | ~v_2293 | ~v_2292 | ~v_2291 | ~v_372 | ~v_371 | ~v_2378 | ~v_2377 | ~v_2376 | ~v_2375 | ~v_330 | ~v_329 | ~v_370 | ~v_369 | ~v_256 | ~v_253 | ~v_368 | ~v_367 | ~v_366 | ~v_365 | ~v_324 | ~v_323 | ~v_322 | ~v_321 | ~v_2761 | ~v_2760 | ~v_2759 | ~v_2758 | v_2774;
assign x_17121 = v_18 | v_17 | v_16 | v_12 | v_135 | v_134 | v_137 | v_179 | v_163 | v_162 | v_161 | v_182 | ~v_361 | ~v_360 | ~v_2235 | ~v_2232 | ~v_2289 | ~v_2288 | ~v_2287 | ~v_2286 | ~v_357 | ~v_356 | ~v_2373 | ~v_2372 | ~v_2371 | ~v_2370 | ~v_315 | ~v_314 | ~v_355 | ~v_354 | ~v_223 | ~v_220 | ~v_353 | ~v_352 | ~v_351 | ~v_350 | ~v_309 | ~v_308 | ~v_307 | ~v_306 | ~v_2756 | ~v_2755 | ~v_2754 | ~v_2753 | v_2773;
assign x_17122 = v_2772 | ~v_2769;
assign x_17123 = v_2772 | ~v_2770;
assign x_17124 = v_2772 | ~v_2771;
assign x_17125 = v_103 | v_95 | v_102 | v_171 | v_170 | v_169 | v_160 | v_150 | v_149 | v_148 | v_184 | v_181 | ~v_2265 | ~v_2262 | ~v_2315 | ~v_2314 | ~v_2313 | ~v_2312 | ~v_297 | ~v_296 | ~v_2383 | ~v_2382 | ~v_2381 | ~v_2380 | ~v_345 | ~v_344 | ~v_343 | ~v_342 | ~v_341 | ~v_340 | ~v_289 | ~v_286 | ~v_285 | ~v_284 | ~v_283 | ~v_282 | ~v_339 | ~v_338 | ~v_337 | ~v_336 | ~v_2766 | ~v_2765 | ~v_2764 | ~v_2763 | v_2771;
assign x_17126 = v_53 | v_61 | v_60 | v_144 | v_180 | v_159 | v_145 | v_143 | v_167 | v_166 | v_165 | v_183 | ~v_2250 | ~v_2247 | ~v_2310 | ~v_2309 | ~v_2308 | ~v_2307 | ~v_264 | ~v_263 | ~v_2378 | ~v_2377 | ~v_2376 | ~v_2375 | ~v_330 | ~v_329 | ~v_328 | ~v_327 | ~v_326 | ~v_325 | ~v_256 | ~v_253 | ~v_252 | ~v_251 | ~v_250 | ~v_249 | ~v_324 | ~v_323 | ~v_322 | ~v_321 | ~v_2761 | ~v_2760 | ~v_2759 | ~v_2758 | v_2770;
assign x_17127 = v_18 | v_17 | v_10 | v_136 | v_135 | v_137 | v_179 | v_163 | v_162 | v_161 | v_155 | v_182 | ~v_2235 | ~v_2232 | ~v_2305 | ~v_2304 | ~v_2303 | ~v_2302 | ~v_231 | ~v_230 | ~v_2373 | ~v_2372 | ~v_2371 | ~v_2370 | ~v_315 | ~v_314 | ~v_313 | ~v_312 | ~v_311 | ~v_310 | ~v_223 | ~v_220 | ~v_219 | ~v_218 | ~v_217 | ~v_216 | ~v_309 | ~v_308 | ~v_307 | ~v_306 | ~v_2756 | ~v_2755 | ~v_2754 | ~v_2753 | v_2769;
assign x_17128 = v_2768 | ~v_2757;
assign x_17129 = v_2768 | ~v_2762;
assign x_17130 = v_2768 | ~v_2767;
assign x_17131 = v_98 | v_103 | v_100 | v_102 | v_170 | v_169 | v_160 | v_150 | v_149 | v_148 | v_147 | v_184 | ~v_2267 | ~v_2266 | ~v_2265 | ~v_2264 | ~v_2263 | ~v_2262 | ~v_299 | ~v_298 | ~v_2315 | ~v_2314 | ~v_2313 | ~v_2312 | ~v_297 | ~v_296 | ~v_295 | ~v_294 | ~v_293 | ~v_292 | ~v_291 | ~v_290 | ~v_289 | ~v_288 | ~v_287 | ~v_286 | ~v_285 | ~v_284 | ~v_283 | ~v_282 | ~v_2766 | ~v_2765 | ~v_2764 | ~v_2763 | v_2767;
assign x_17132 = v_2766 | v_173;
assign x_17133 = v_2766 | v_123;
assign x_17134 = v_2765 | v_174;
assign x_17135 = v_2765 | v_120;
assign x_17136 = v_2764 | ~v_173;
assign x_17137 = v_2764 | v_108;
assign x_17138 = v_2763 | ~v_174;
assign x_17139 = v_2763 | v_105;
assign x_17140 = v_56 | v_61 | v_60 | v_58 | v_144 | v_159 | v_145 | v_143 | v_142 | v_166 | v_165 | v_183 | ~v_266 | ~v_2252 | ~v_2251 | ~v_2250 | ~v_2249 | ~v_2248 | ~v_2247 | ~v_265 | ~v_2310 | ~v_2309 | ~v_2308 | ~v_2307 | ~v_264 | ~v_263 | ~v_262 | ~v_261 | ~v_260 | ~v_259 | ~v_258 | ~v_257 | ~v_256 | ~v_255 | ~v_254 | ~v_253 | ~v_252 | ~v_251 | ~v_250 | ~v_249 | ~v_2761 | ~v_2760 | ~v_2759 | ~v_2758 | v_2762;
assign x_17141 = v_2761 | v_173;
assign x_17142 = v_2761 | v_81;
assign x_17143 = v_2760 | v_174;
assign x_17144 = v_2760 | v_78;
assign x_17145 = v_2759 | ~v_173;
assign x_17146 = v_2759 | v_66;
assign x_17147 = v_2758 | ~v_174;
assign x_17148 = v_2758 | v_63;
assign x_17149 = v_13 | v_18 | v_17 | v_15 | v_136 | v_135 | v_134 | v_137 | v_162 | v_161 | v_155 | v_182 | ~v_2237 | ~v_2236 | ~v_2235 | ~v_2234 | ~v_2233 | ~v_2232 | ~v_233 | ~v_232 | ~v_2305 | ~v_2304 | ~v_2303 | ~v_2302 | ~v_231 | ~v_230 | ~v_229 | ~v_228 | ~v_227 | ~v_226 | ~v_225 | ~v_224 | ~v_223 | ~v_222 | ~v_221 | ~v_220 | ~v_219 | ~v_218 | ~v_217 | ~v_216 | ~v_2756 | ~v_2755 | ~v_2754 | ~v_2753 | v_2757;
assign x_17150 = v_2756 | v_173;
assign x_17151 = v_2756 | v_39;
assign x_17152 = v_2755 | v_174;
assign x_17153 = v_2755 | v_36;
assign x_17154 = v_2754 | ~v_173;
assign x_17155 = v_2754 | v_24;
assign x_17156 = v_2753 | ~v_174;
assign x_17157 = v_2753 | v_21;
assign x_17158 = v_2752 | ~v_2750;
assign x_17159 = v_2752 | ~v_2751;
assign x_17160 = v_2752 | ~v_1270;
assign x_17161 = v_2752 | ~v_1271;
assign x_17162 = v_2752 | ~v_174;
assign x_17163 = v_2752 | ~v_173;
assign x_17164 = ~v_193 | ~v_2221 | v_2751;
assign x_17165 = ~v_188 | ~v_191 | v_2750;
assign x_17166 = v_2749 | ~v_2668;
assign x_17167 = v_2749 | ~v_2748;
assign x_17168 = v_174 | v_173 | ~v_2747 | ~v_1561 | ~v_1560 | ~v_2670 | ~v_2669 | v_2748;
assign x_17169 = v_2747 | ~v_2686;
assign x_17170 = v_2747 | ~v_2690;
assign x_17171 = v_2747 | ~v_2694;
assign x_17172 = v_2747 | ~v_2698;
assign x_17173 = v_2747 | ~v_2702;
assign x_17174 = v_2747 | ~v_2706;
assign x_17175 = v_2747 | ~v_2710;
assign x_17176 = v_2747 | ~v_2714;
assign x_17177 = v_2747 | ~v_2718;
assign x_17178 = v_2747 | ~v_2722;
assign x_17179 = v_2747 | ~v_2726;
assign x_17180 = v_2747 | ~v_2730;
assign x_17181 = v_2747 | ~v_2734;
assign x_17182 = v_2747 | ~v_2738;
assign x_17183 = v_2747 | ~v_2742;
assign x_17184 = v_2747 | ~v_2746;
assign x_17185 = v_2747 | ~v_1263;
assign x_17186 = v_2747 | ~v_1264;
assign x_17187 = v_2747 | ~v_1265;
assign x_17188 = v_2747 | ~v_1266;
assign x_17189 = ~v_2745 | ~v_2744 | ~v_2743 | v_2746;
assign x_17190 = v_2745 | ~v_2681;
assign x_17191 = v_2745 | ~v_2682;
assign x_17192 = v_2745 | ~v_2683;
assign x_17193 = v_2745 | ~v_2684;
assign x_17194 = v_2745 | ~v_1636;
assign x_17195 = v_2745 | ~v_1637;
assign x_17196 = v_2745 | ~v_1750;
assign x_17197 = v_2745 | ~v_1638;
assign x_17198 = v_2745 | ~v_1751;
assign x_17199 = v_2745 | ~v_1639;
assign x_17200 = v_2745 | ~v_1640;
assign x_17201 = v_2745 | ~v_1752;
assign x_17202 = v_2745 | ~v_1641;
assign x_17203 = v_2745 | ~v_1753;
assign x_17204 = v_2745 | ~v_2075;
assign x_17205 = v_2745 | ~v_2076;
assign x_17206 = v_2745 | ~v_2141;
assign x_17207 = v_2745 | ~v_2077;
assign x_17208 = v_2745 | ~v_2142;
assign x_17209 = v_2745 | ~v_2078;
assign x_17210 = v_2745 | ~v_2079;
assign x_17211 = v_2745 | ~v_2143;
assign x_17212 = v_2745 | ~v_2080;
assign x_17213 = v_2745 | ~v_2144;
assign x_17214 = v_2745 | ~v_839;
assign x_17215 = v_2745 | ~v_1257;
assign x_17216 = v_2745 | ~v_1023;
assign x_17217 = v_2745 | ~v_840;
assign x_17218 = v_2745 | ~v_1258;
assign x_17219 = v_2745 | ~v_1024;
assign x_17220 = v_2745 | ~v_184;
assign x_17221 = v_2745 | ~v_170;
assign x_17222 = v_2745 | ~v_169;
assign x_17223 = v_2745 | ~v_149;
assign x_17224 = v_2745 | ~v_148;
assign x_17225 = v_2745 | ~v_1259;
assign x_17226 = v_2745 | ~v_1260;
assign x_17227 = v_2745 | ~v_103;
assign x_17228 = v_2745 | ~v_102;
assign x_17229 = v_2745 | ~v_101;
assign x_17230 = v_2745 | ~v_100;
assign x_17231 = v_2745 | ~v_99;
assign x_17232 = v_2745 | ~v_98;
assign x_17233 = v_2745 | ~v_95;
assign x_17234 = v_2744 | ~v_2676;
assign x_17235 = v_2744 | ~v_2677;
assign x_17236 = v_2744 | ~v_2678;
assign x_17237 = v_2744 | ~v_2679;
assign x_17238 = v_2744 | ~v_1611;
assign x_17239 = v_2744 | ~v_1612;
assign x_17240 = v_2744 | ~v_1741;
assign x_17241 = v_2744 | ~v_1613;
assign x_17242 = v_2744 | ~v_1742;
assign x_17243 = v_2744 | ~v_1614;
assign x_17244 = v_2744 | ~v_1615;
assign x_17245 = v_2744 | ~v_1743;
assign x_17246 = v_2744 | ~v_1616;
assign x_17247 = v_2744 | ~v_1744;
assign x_17248 = v_2744 | ~v_2060;
assign x_17249 = v_2744 | ~v_2061;
assign x_17250 = v_2744 | ~v_2136;
assign x_17251 = v_2744 | ~v_2062;
assign x_17252 = v_2744 | ~v_2137;
assign x_17253 = v_2744 | ~v_2063;
assign x_17254 = v_2744 | ~v_2064;
assign x_17255 = v_2744 | ~v_2138;
assign x_17256 = v_2744 | ~v_2065;
assign x_17257 = v_2744 | ~v_2139;
assign x_17258 = v_2744 | ~v_806;
assign x_17259 = v_2744 | ~v_1252;
assign x_17260 = v_2744 | ~v_1008;
assign x_17261 = v_2744 | ~v_1253;
assign x_17262 = v_2744 | ~v_1009;
assign x_17263 = v_2744 | ~v_807;
assign x_17264 = v_2744 | ~v_183;
assign x_17265 = v_2744 | ~v_166;
assign x_17266 = v_2744 | ~v_165;
assign x_17267 = v_2744 | ~v_144;
assign x_17268 = v_2744 | ~v_143;
assign x_17269 = v_2744 | ~v_1254;
assign x_17270 = v_2744 | ~v_1255;
assign x_17271 = v_2744 | ~v_61;
assign x_17272 = v_2744 | ~v_60;
assign x_17273 = v_2744 | ~v_59;
assign x_17274 = v_2744 | ~v_58;
assign x_17275 = v_2744 | ~v_57;
assign x_17276 = v_2744 | ~v_56;
assign x_17277 = v_2744 | ~v_53;
assign x_17278 = v_2743 | ~v_2671;
assign x_17279 = v_2743 | ~v_2672;
assign x_17280 = v_2743 | ~v_2673;
assign x_17281 = v_2743 | ~v_2674;
assign x_17282 = v_2743 | ~v_1586;
assign x_17283 = v_2743 | ~v_1587;
assign x_17284 = v_2743 | ~v_1732;
assign x_17285 = v_2743 | ~v_1588;
assign x_17286 = v_2743 | ~v_1733;
assign x_17287 = v_2743 | ~v_1589;
assign x_17288 = v_2743 | ~v_1590;
assign x_17289 = v_2743 | ~v_1734;
assign x_17290 = v_2743 | ~v_1591;
assign x_17291 = v_2743 | ~v_1735;
assign x_17292 = v_2743 | ~v_2045;
assign x_17293 = v_2743 | ~v_2046;
assign x_17294 = v_2743 | ~v_2131;
assign x_17295 = v_2743 | ~v_2047;
assign x_17296 = v_2743 | ~v_2132;
assign x_17297 = v_2743 | ~v_2048;
assign x_17298 = v_2743 | ~v_2049;
assign x_17299 = v_2743 | ~v_2133;
assign x_17300 = v_2743 | ~v_2050;
assign x_17301 = v_2743 | ~v_2134;
assign x_17302 = v_2743 | ~v_773;
assign x_17303 = v_2743 | ~v_774;
assign x_17304 = v_2743 | ~v_182;
assign x_17305 = v_2743 | ~v_162;
assign x_17306 = v_2743 | ~v_161;
assign x_17307 = v_2743 | ~v_1247;
assign x_17308 = v_2743 | ~v_1248;
assign x_17309 = v_2743 | ~v_136;
assign x_17310 = v_2743 | ~v_135;
assign x_17311 = v_2743 | ~v_1249;
assign x_17312 = v_2743 | ~v_993;
assign x_17313 = v_2743 | ~v_1250;
assign x_17314 = v_2743 | ~v_994;
assign x_17315 = v_2743 | ~v_18;
assign x_17316 = v_2743 | ~v_17;
assign x_17317 = v_2743 | ~v_16;
assign x_17318 = v_2743 | ~v_15;
assign x_17319 = v_2743 | ~v_14;
assign x_17320 = v_2743 | ~v_13;
assign x_17321 = v_2743 | ~v_10;
assign x_17322 = ~v_2741 | ~v_2740 | ~v_2739 | v_2742;
assign x_17323 = v_2741 | ~v_2681;
assign x_17324 = v_2741 | ~v_2682;
assign x_17325 = v_2741 | ~v_2683;
assign x_17326 = v_2741 | ~v_2684;
assign x_17327 = v_2741 | ~v_1782;
assign x_17328 = v_2741 | ~v_1783;
assign x_17329 = v_2741 | ~v_1784;
assign x_17330 = v_2741 | ~v_1785;
assign x_17331 = v_2741 | ~v_1636;
assign x_17332 = v_2741 | ~v_1750;
assign x_17333 = v_2741 | ~v_1751;
assign x_17334 = v_2741 | ~v_1639;
assign x_17335 = v_2741 | ~v_1752;
assign x_17336 = v_2741 | ~v_1753;
assign x_17337 = v_2741 | ~v_2193;
assign x_17338 = v_2741 | ~v_2194;
assign x_17339 = v_2741 | ~v_2195;
assign x_17340 = v_2741 | ~v_2196;
assign x_17341 = v_2741 | ~v_2075;
assign x_17342 = v_2741 | ~v_2141;
assign x_17343 = v_2741 | ~v_2142;
assign x_17344 = v_2741 | ~v_2078;
assign x_17345 = v_2741 | ~v_2143;
assign x_17346 = v_2741 | ~v_2144;
assign x_17347 = v_2741 | ~v_1085;
assign x_17348 = v_2741 | ~v_1131;
assign x_17349 = v_2741 | ~v_1132;
assign x_17350 = v_2741 | ~v_1086;
assign x_17351 = v_2741 | ~v_1133;
assign x_17352 = v_2741 | ~v_1134;
assign x_17353 = v_2741 | ~v_1023;
assign x_17354 = v_2741 | ~v_1024;
assign x_17355 = v_2741 | ~v_184;
assign x_17356 = v_2741 | ~v_172;
assign x_17357 = v_2741 | ~v_171;
assign x_17358 = v_2741 | ~v_170;
assign x_17359 = v_2741 | ~v_149;
assign x_17360 = v_2741 | ~v_148;
assign x_17361 = v_2741 | ~v_147;
assign x_17362 = v_2741 | ~v_102;
assign x_17363 = v_2741 | ~v_101;
assign x_17364 = v_2741 | ~v_100;
assign x_17365 = v_2741 | ~v_99;
assign x_17366 = v_2741 | ~v_93;
assign x_17367 = v_2740 | ~v_2676;
assign x_17368 = v_2740 | ~v_2677;
assign x_17369 = v_2740 | ~v_2678;
assign x_17370 = v_2740 | ~v_2679;
assign x_17371 = v_2740 | ~v_1773;
assign x_17372 = v_2740 | ~v_1774;
assign x_17373 = v_2740 | ~v_1775;
assign x_17374 = v_2740 | ~v_1776;
assign x_17375 = v_2740 | ~v_1611;
assign x_17376 = v_2740 | ~v_1741;
assign x_17377 = v_2740 | ~v_1742;
assign x_17378 = v_2740 | ~v_1614;
assign x_17379 = v_2740 | ~v_1743;
assign x_17380 = v_2740 | ~v_1744;
assign x_17381 = v_2740 | ~v_2188;
assign x_17382 = v_2740 | ~v_2189;
assign x_17383 = v_2740 | ~v_2190;
assign x_17384 = v_2740 | ~v_2191;
assign x_17385 = v_2740 | ~v_2060;
assign x_17386 = v_2740 | ~v_2136;
assign x_17387 = v_2740 | ~v_2137;
assign x_17388 = v_2740 | ~v_2063;
assign x_17389 = v_2740 | ~v_2138;
assign x_17390 = v_2740 | ~v_2139;
assign x_17391 = v_2740 | ~v_1070;
assign x_17392 = v_2740 | ~v_1126;
assign x_17393 = v_2740 | ~v_1127;
assign x_17394 = v_2740 | ~v_1071;
assign x_17395 = v_2740 | ~v_1128;
assign x_17396 = v_2740 | ~v_1129;
assign x_17397 = v_2740 | ~v_1008;
assign x_17398 = v_2740 | ~v_1009;
assign x_17399 = v_2740 | ~v_183;
assign x_17400 = v_2740 | ~v_168;
assign x_17401 = v_2740 | ~v_167;
assign x_17402 = v_2740 | ~v_166;
assign x_17403 = v_2740 | ~v_144;
assign x_17404 = v_2740 | ~v_143;
assign x_17405 = v_2740 | ~v_142;
assign x_17406 = v_2740 | ~v_60;
assign x_17407 = v_2740 | ~v_59;
assign x_17408 = v_2740 | ~v_58;
assign x_17409 = v_2740 | ~v_57;
assign x_17410 = v_2740 | ~v_51;
assign x_17411 = v_2739 | ~v_2671;
assign x_17412 = v_2739 | ~v_2672;
assign x_17413 = v_2739 | ~v_2673;
assign x_17414 = v_2739 | ~v_2674;
assign x_17415 = v_2739 | ~v_1764;
assign x_17416 = v_2739 | ~v_1765;
assign x_17417 = v_2739 | ~v_1766;
assign x_17418 = v_2739 | ~v_1767;
assign x_17419 = v_2739 | ~v_1586;
assign x_17420 = v_2739 | ~v_1732;
assign x_17421 = v_2739 | ~v_1733;
assign x_17422 = v_2739 | ~v_1589;
assign x_17423 = v_2739 | ~v_1734;
assign x_17424 = v_2739 | ~v_1735;
assign x_17425 = v_2739 | ~v_2183;
assign x_17426 = v_2739 | ~v_2184;
assign x_17427 = v_2739 | ~v_2185;
assign x_17428 = v_2739 | ~v_2186;
assign x_17429 = v_2739 | ~v_2045;
assign x_17430 = v_2739 | ~v_2131;
assign x_17431 = v_2739 | ~v_2132;
assign x_17432 = v_2739 | ~v_2048;
assign x_17433 = v_2739 | ~v_2133;
assign x_17434 = v_2739 | ~v_2134;
assign x_17435 = v_2739 | ~v_1055;
assign x_17436 = v_2739 | ~v_1121;
assign x_17437 = v_2739 | ~v_1122;
assign x_17438 = v_2739 | ~v_1056;
assign x_17439 = v_2739 | ~v_1123;
assign x_17440 = v_2739 | ~v_1124;
assign x_17441 = v_2739 | ~v_182;
assign x_17442 = v_2739 | ~v_164;
assign x_17443 = v_2739 | ~v_163;
assign x_17444 = v_2739 | ~v_162;
assign x_17445 = v_2739 | ~v_136;
assign x_17446 = v_2739 | ~v_135;
assign x_17447 = v_2739 | ~v_134;
assign x_17448 = v_2739 | ~v_993;
assign x_17449 = v_2739 | ~v_994;
assign x_17450 = v_2739 | ~v_17;
assign x_17451 = v_2739 | ~v_16;
assign x_17452 = v_2739 | ~v_15;
assign x_17453 = v_2739 | ~v_14;
assign x_17454 = v_2739 | ~v_8;
assign x_17455 = ~v_2737 | ~v_2736 | ~v_2735 | v_2738;
assign x_17456 = v_2737 | ~v_2681;
assign x_17457 = v_2737 | ~v_2682;
assign x_17458 = v_2737 | ~v_2683;
assign x_17459 = v_2737 | ~v_2684;
assign x_17460 = v_2737 | ~v_1782;
assign x_17461 = v_2737 | ~v_1783;
assign x_17462 = v_2737 | ~v_1784;
assign x_17463 = v_2737 | ~v_1785;
assign x_17464 = v_2737 | ~v_1694;
assign x_17465 = v_2737 | ~v_1695;
assign x_17466 = v_2737 | ~v_1696;
assign x_17467 = v_2737 | ~v_1697;
assign x_17468 = v_2737 | ~v_1636;
assign x_17469 = v_2737 | ~v_1639;
assign x_17470 = v_2737 | ~v_2125;
assign x_17471 = v_2737 | ~v_2126;
assign x_17472 = v_2737 | ~v_2127;
assign x_17473 = v_2737 | ~v_2128;
assign x_17474 = v_2737 | ~v_2193;
assign x_17475 = v_2737 | ~v_2194;
assign x_17476 = v_2737 | ~v_2195;
assign x_17477 = v_2737 | ~v_2196;
assign x_17478 = v_2737 | ~v_2075;
assign x_17479 = v_2737 | ~v_2078;
assign x_17480 = v_2737 | ~v_927;
assign x_17481 = v_2737 | ~v_928;
assign x_17482 = v_2737 | ~v_1099;
assign x_17483 = v_2737 | ~v_1100;
assign x_17484 = v_2737 | ~v_1101;
assign x_17485 = v_2737 | ~v_1102;
assign x_17486 = v_2737 | ~v_1085;
assign x_17487 = v_2737 | ~v_1086;
assign x_17488 = v_2737 | ~v_184;
assign x_17489 = v_2737 | ~v_171;
assign x_17490 = v_2737 | ~v_170;
assign x_17491 = v_2737 | ~v_150;
assign x_17492 = v_2737 | ~v_149;
assign x_17493 = v_2737 | ~v_103;
assign x_17494 = v_2737 | ~v_102;
assign x_17495 = v_2737 | ~v_101;
assign x_17496 = v_2737 | ~v_100;
assign x_17497 = v_2737 | ~v_96;
assign x_17498 = v_2737 | ~v_95;
assign x_17499 = v_2737 | ~v_93;
assign x_17500 = v_2736 | ~v_2676;
assign x_17501 = v_2736 | ~v_2677;
assign x_17502 = v_2736 | ~v_2678;
assign x_17503 = v_2736 | ~v_2679;
assign x_17504 = v_2736 | ~v_1773;
assign x_17505 = v_2736 | ~v_1774;
assign x_17506 = v_2736 | ~v_1775;
assign x_17507 = v_2736 | ~v_1776;
assign x_17508 = v_2736 | ~v_1685;
assign x_17509 = v_2736 | ~v_1686;
assign x_17510 = v_2736 | ~v_1687;
assign x_17511 = v_2736 | ~v_1688;
assign x_17512 = v_2736 | ~v_1611;
assign x_17513 = v_2736 | ~v_1614;
assign x_17514 = v_2736 | ~v_2120;
assign x_17515 = v_2736 | ~v_2121;
assign x_17516 = v_2736 | ~v_2122;
assign x_17517 = v_2736 | ~v_2123;
assign x_17518 = v_2736 | ~v_2188;
assign x_17519 = v_2736 | ~v_2189;
assign x_17520 = v_2736 | ~v_2190;
assign x_17521 = v_2736 | ~v_2191;
assign x_17522 = v_2736 | ~v_2060;
assign x_17523 = v_2736 | ~v_2063;
assign x_17524 = v_2736 | ~v_912;
assign x_17525 = v_2736 | ~v_913;
assign x_17526 = v_2736 | ~v_1094;
assign x_17527 = v_2736 | ~v_1095;
assign x_17528 = v_2736 | ~v_1096;
assign x_17529 = v_2736 | ~v_1097;
assign x_17530 = v_2736 | ~v_1070;
assign x_17531 = v_2736 | ~v_1071;
assign x_17532 = v_2736 | ~v_183;
assign x_17533 = v_2736 | ~v_167;
assign x_17534 = v_2736 | ~v_166;
assign x_17535 = v_2736 | ~v_145;
assign x_17536 = v_2736 | ~v_144;
assign x_17537 = v_2736 | ~v_61;
assign x_17538 = v_2736 | ~v_60;
assign x_17539 = v_2736 | ~v_59;
assign x_17540 = v_2736 | ~v_58;
assign x_17541 = v_2736 | ~v_54;
assign x_17542 = v_2736 | ~v_53;
assign x_17543 = v_2736 | ~v_51;
assign x_17544 = v_2735 | ~v_2671;
assign x_17545 = v_2735 | ~v_2672;
assign x_17546 = v_2735 | ~v_2673;
assign x_17547 = v_2735 | ~v_2674;
assign x_17548 = v_2735 | ~v_1764;
assign x_17549 = v_2735 | ~v_1765;
assign x_17550 = v_2735 | ~v_1766;
assign x_17551 = v_2735 | ~v_1767;
assign x_17552 = v_2735 | ~v_1676;
assign x_17553 = v_2735 | ~v_1677;
assign x_17554 = v_2735 | ~v_1678;
assign x_17555 = v_2735 | ~v_1679;
assign x_17556 = v_2735 | ~v_1586;
assign x_17557 = v_2735 | ~v_1589;
assign x_17558 = v_2735 | ~v_2115;
assign x_17559 = v_2735 | ~v_2116;
assign x_17560 = v_2735 | ~v_2117;
assign x_17561 = v_2735 | ~v_2118;
assign x_17562 = v_2735 | ~v_2183;
assign x_17563 = v_2735 | ~v_2184;
assign x_17564 = v_2735 | ~v_2185;
assign x_17565 = v_2735 | ~v_2186;
assign x_17566 = v_2735 | ~v_2045;
assign x_17567 = v_2735 | ~v_2048;
assign x_17568 = v_2735 | ~v_897;
assign x_17569 = v_2735 | ~v_898;
assign x_17570 = v_2735 | ~v_1089;
assign x_17571 = v_2735 | ~v_1090;
assign x_17572 = v_2735 | ~v_1091;
assign x_17573 = v_2735 | ~v_1092;
assign x_17574 = v_2735 | ~v_1055;
assign x_17575 = v_2735 | ~v_1056;
assign x_17576 = v_2735 | ~v_182;
assign x_17577 = v_2735 | ~v_163;
assign x_17578 = v_2735 | ~v_162;
assign x_17579 = v_2735 | ~v_137;
assign x_17580 = v_2735 | ~v_136;
assign x_17581 = v_2735 | ~v_18;
assign x_17582 = v_2735 | ~v_17;
assign x_17583 = v_2735 | ~v_16;
assign x_17584 = v_2735 | ~v_15;
assign x_17585 = v_2735 | ~v_11;
assign x_17586 = v_2735 | ~v_10;
assign x_17587 = v_2735 | ~v_8;
assign x_17588 = ~v_2733 | ~v_2732 | ~v_2731 | v_2734;
assign x_17589 = v_2733 | ~v_2681;
assign x_17590 = v_2733 | ~v_2682;
assign x_17591 = v_2733 | ~v_2683;
assign x_17592 = v_2733 | ~v_2684;
assign x_17593 = v_2733 | ~v_1782;
assign x_17594 = v_2733 | ~v_1783;
assign x_17595 = v_2733 | ~v_1784;
assign x_17596 = v_2733 | ~v_1785;
assign x_17597 = v_2733 | ~v_1632;
assign x_17598 = v_2733 | ~v_1633;
assign x_17599 = v_2733 | ~v_1634;
assign x_17600 = v_2733 | ~v_1635;
assign x_17601 = v_2733 | ~v_1636;
assign x_17602 = v_2733 | ~v_1639;
assign x_17603 = v_2733 | ~v_2109;
assign x_17604 = v_2733 | ~v_2110;
assign x_17605 = v_2733 | ~v_2111;
assign x_17606 = v_2733 | ~v_2112;
assign x_17607 = v_2733 | ~v_2193;
assign x_17608 = v_2733 | ~v_2194;
assign x_17609 = v_2733 | ~v_2195;
assign x_17610 = v_2733 | ~v_2196;
assign x_17611 = v_2733 | ~v_2075;
assign x_17612 = v_2733 | ~v_2078;
assign x_17613 = v_2733 | ~v_975;
assign x_17614 = v_2733 | ~v_976;
assign x_17615 = v_2733 | ~v_1115;
assign x_17616 = v_2733 | ~v_1116;
assign x_17617 = v_2733 | ~v_1085;
assign x_17618 = v_2733 | ~v_1086;
assign x_17619 = v_2733 | ~v_1117;
assign x_17620 = v_2733 | ~v_1118;
assign x_17621 = v_2733 | ~v_184;
assign x_17622 = v_2733 | ~v_171;
assign x_17623 = v_2733 | ~v_170;
assign x_17624 = v_2733 | ~v_151;
assign x_17625 = v_2733 | ~v_150;
assign x_17626 = v_2733 | ~v_148;
assign x_17627 = v_2733 | ~v_147;
assign x_17628 = v_2733 | ~v_103;
assign x_17629 = v_2733 | ~v_101;
assign x_17630 = v_2733 | ~v_100;
assign x_17631 = v_2733 | ~v_97;
assign x_17632 = v_2733 | ~v_93;
assign x_17633 = v_2732 | ~v_2676;
assign x_17634 = v_2732 | ~v_2677;
assign x_17635 = v_2732 | ~v_2678;
assign x_17636 = v_2732 | ~v_2679;
assign x_17637 = v_2732 | ~v_1773;
assign x_17638 = v_2732 | ~v_1774;
assign x_17639 = v_2732 | ~v_1775;
assign x_17640 = v_2732 | ~v_1776;
assign x_17641 = v_2732 | ~v_1607;
assign x_17642 = v_2732 | ~v_1608;
assign x_17643 = v_2732 | ~v_1609;
assign x_17644 = v_2732 | ~v_1610;
assign x_17645 = v_2732 | ~v_1611;
assign x_17646 = v_2732 | ~v_1614;
assign x_17647 = v_2732 | ~v_2104;
assign x_17648 = v_2732 | ~v_2105;
assign x_17649 = v_2732 | ~v_2106;
assign x_17650 = v_2732 | ~v_2107;
assign x_17651 = v_2732 | ~v_2188;
assign x_17652 = v_2732 | ~v_2189;
assign x_17653 = v_2732 | ~v_2190;
assign x_17654 = v_2732 | ~v_2191;
assign x_17655 = v_2732 | ~v_2060;
assign x_17656 = v_2732 | ~v_2063;
assign x_17657 = v_2732 | ~v_960;
assign x_17658 = v_2732 | ~v_961;
assign x_17659 = v_2732 | ~v_1110;
assign x_17660 = v_2732 | ~v_1111;
assign x_17661 = v_2732 | ~v_1070;
assign x_17662 = v_2732 | ~v_1071;
assign x_17663 = v_2732 | ~v_1112;
assign x_17664 = v_2732 | ~v_1113;
assign x_17665 = v_2732 | ~v_183;
assign x_17666 = v_2732 | ~v_167;
assign x_17667 = v_2732 | ~v_166;
assign x_17668 = v_2732 | ~v_146;
assign x_17669 = v_2732 | ~v_145;
assign x_17670 = v_2732 | ~v_143;
assign x_17671 = v_2732 | ~v_142;
assign x_17672 = v_2732 | ~v_61;
assign x_17673 = v_2732 | ~v_59;
assign x_17674 = v_2732 | ~v_58;
assign x_17675 = v_2732 | ~v_55;
assign x_17676 = v_2732 | ~v_51;
assign x_17677 = v_2731 | ~v_2671;
assign x_17678 = v_2731 | ~v_2672;
assign x_17679 = v_2731 | ~v_2673;
assign x_17680 = v_2731 | ~v_2674;
assign x_17681 = v_2731 | ~v_1764;
assign x_17682 = v_2731 | ~v_1765;
assign x_17683 = v_2731 | ~v_1766;
assign x_17684 = v_2731 | ~v_1767;
assign x_17685 = v_2731 | ~v_1582;
assign x_17686 = v_2731 | ~v_1583;
assign x_17687 = v_2731 | ~v_1584;
assign x_17688 = v_2731 | ~v_1585;
assign x_17689 = v_2731 | ~v_1586;
assign x_17690 = v_2731 | ~v_1589;
assign x_17691 = v_2731 | ~v_2099;
assign x_17692 = v_2731 | ~v_2100;
assign x_17693 = v_2731 | ~v_2101;
assign x_17694 = v_2731 | ~v_2102;
assign x_17695 = v_2731 | ~v_2183;
assign x_17696 = v_2731 | ~v_2184;
assign x_17697 = v_2731 | ~v_2185;
assign x_17698 = v_2731 | ~v_2186;
assign x_17699 = v_2731 | ~v_2045;
assign x_17700 = v_2731 | ~v_2048;
assign x_17701 = v_2731 | ~v_945;
assign x_17702 = v_2731 | ~v_946;
assign x_17703 = v_2731 | ~v_1105;
assign x_17704 = v_2731 | ~v_1106;
assign x_17705 = v_2731 | ~v_1055;
assign x_17706 = v_2731 | ~v_1056;
assign x_17707 = v_2731 | ~v_1107;
assign x_17708 = v_2731 | ~v_1108;
assign x_17709 = v_2731 | ~v_182;
assign x_17710 = v_2731 | ~v_163;
assign x_17711 = v_2731 | ~v_162;
assign x_17712 = v_2731 | ~v_138;
assign x_17713 = v_2731 | ~v_137;
assign x_17714 = v_2731 | ~v_135;
assign x_17715 = v_2731 | ~v_134;
assign x_17716 = v_2731 | ~v_18;
assign x_17717 = v_2731 | ~v_16;
assign x_17718 = v_2731 | ~v_15;
assign x_17719 = v_2731 | ~v_12;
assign x_17720 = v_2731 | ~v_8;
assign x_17721 = ~v_2729 | ~v_2728 | ~v_2727 | v_2730;
assign x_17722 = v_2729 | ~v_2681;
assign x_17723 = v_2729 | ~v_2682;
assign x_17724 = v_2729 | ~v_2683;
assign x_17725 = v_2729 | ~v_2684;
assign x_17726 = v_2729 | ~v_1782;
assign x_17727 = v_2729 | ~v_1783;
assign x_17728 = v_2729 | ~v_1784;
assign x_17729 = v_2729 | ~v_1785;
assign x_17730 = v_2729 | ~v_1722;
assign x_17731 = v_2729 | ~v_1723;
assign x_17732 = v_2729 | ~v_1724;
assign x_17733 = v_2729 | ~v_1725;
assign x_17734 = v_2729 | ~v_1636;
assign x_17735 = v_2729 | ~v_1639;
assign x_17736 = v_2729 | ~v_2071;
assign x_17737 = v_2729 | ~v_2072;
assign x_17738 = v_2729 | ~v_2073;
assign x_17739 = v_2729 | ~v_2074;
assign x_17740 = v_2729 | ~v_2193;
assign x_17741 = v_2729 | ~v_2194;
assign x_17742 = v_2729 | ~v_2195;
assign x_17743 = v_2729 | ~v_2196;
assign x_17744 = v_2729 | ~v_2075;
assign x_17745 = v_2729 | ~v_2078;
assign x_17746 = v_2729 | ~v_837;
assign x_17747 = v_2729 | ~v_838;
assign x_17748 = v_2729 | ~v_1081;
assign x_17749 = v_2729 | ~v_1082;
assign x_17750 = v_2729 | ~v_1083;
assign x_17751 = v_2729 | ~v_1084;
assign x_17752 = v_2729 | ~v_1085;
assign x_17753 = v_2729 | ~v_1086;
assign x_17754 = v_2729 | ~v_184;
assign x_17755 = v_2729 | ~v_171;
assign x_17756 = v_2729 | ~v_170;
assign x_17757 = v_2729 | ~v_160;
assign x_17758 = v_2729 | ~v_150;
assign x_17759 = v_2729 | ~v_149;
assign x_17760 = v_2729 | ~v_148;
assign x_17761 = v_2729 | ~v_147;
assign x_17762 = v_2729 | ~v_103;
assign x_17763 = v_2729 | ~v_102;
assign x_17764 = v_2729 | ~v_100;
assign x_17765 = v_2729 | ~v_93;
assign x_17766 = v_2728 | ~v_2676;
assign x_17767 = v_2728 | ~v_2677;
assign x_17768 = v_2728 | ~v_2678;
assign x_17769 = v_2728 | ~v_2679;
assign x_17770 = v_2728 | ~v_1773;
assign x_17771 = v_2728 | ~v_1774;
assign x_17772 = v_2728 | ~v_1775;
assign x_17773 = v_2728 | ~v_1776;
assign x_17774 = v_2728 | ~v_1713;
assign x_17775 = v_2728 | ~v_1714;
assign x_17776 = v_2728 | ~v_1715;
assign x_17777 = v_2728 | ~v_1716;
assign x_17778 = v_2728 | ~v_1611;
assign x_17779 = v_2728 | ~v_1614;
assign x_17780 = v_2728 | ~v_2056;
assign x_17781 = v_2728 | ~v_2057;
assign x_17782 = v_2728 | ~v_2058;
assign x_17783 = v_2728 | ~v_2059;
assign x_17784 = v_2728 | ~v_2188;
assign x_17785 = v_2728 | ~v_2189;
assign x_17786 = v_2728 | ~v_2190;
assign x_17787 = v_2728 | ~v_2191;
assign x_17788 = v_2728 | ~v_2060;
assign x_17789 = v_2728 | ~v_2063;
assign x_17790 = v_2728 | ~v_804;
assign x_17791 = v_2728 | ~v_805;
assign x_17792 = v_2728 | ~v_1066;
assign x_17793 = v_2728 | ~v_1067;
assign x_17794 = v_2728 | ~v_1068;
assign x_17795 = v_2728 | ~v_1069;
assign x_17796 = v_2728 | ~v_1070;
assign x_17797 = v_2728 | ~v_1071;
assign x_17798 = v_2728 | ~v_183;
assign x_17799 = v_2728 | ~v_167;
assign x_17800 = v_2728 | ~v_166;
assign x_17801 = v_2728 | ~v_159;
assign x_17802 = v_2728 | ~v_145;
assign x_17803 = v_2728 | ~v_144;
assign x_17804 = v_2728 | ~v_143;
assign x_17805 = v_2728 | ~v_142;
assign x_17806 = v_2728 | ~v_61;
assign x_17807 = v_2728 | ~v_60;
assign x_17808 = v_2728 | ~v_58;
assign x_17809 = v_2728 | ~v_51;
assign x_17810 = v_2727 | ~v_2671;
assign x_17811 = v_2727 | ~v_2672;
assign x_17812 = v_2727 | ~v_2673;
assign x_17813 = v_2727 | ~v_2674;
assign x_17814 = v_2727 | ~v_1764;
assign x_17815 = v_2727 | ~v_1765;
assign x_17816 = v_2727 | ~v_1766;
assign x_17817 = v_2727 | ~v_1767;
assign x_17818 = v_2727 | ~v_1704;
assign x_17819 = v_2727 | ~v_1705;
assign x_17820 = v_2727 | ~v_1706;
assign x_17821 = v_2727 | ~v_1707;
assign x_17822 = v_2727 | ~v_1586;
assign x_17823 = v_2727 | ~v_1589;
assign x_17824 = v_2727 | ~v_2041;
assign x_17825 = v_2727 | ~v_2042;
assign x_17826 = v_2727 | ~v_2043;
assign x_17827 = v_2727 | ~v_2044;
assign x_17828 = v_2727 | ~v_2183;
assign x_17829 = v_2727 | ~v_2184;
assign x_17830 = v_2727 | ~v_2185;
assign x_17831 = v_2727 | ~v_2186;
assign x_17832 = v_2727 | ~v_2045;
assign x_17833 = v_2727 | ~v_2048;
assign x_17834 = v_2727 | ~v_771;
assign x_17835 = v_2727 | ~v_772;
assign x_17836 = v_2727 | ~v_1051;
assign x_17837 = v_2727 | ~v_1052;
assign x_17838 = v_2727 | ~v_1053;
assign x_17839 = v_2727 | ~v_1054;
assign x_17840 = v_2727 | ~v_1055;
assign x_17841 = v_2727 | ~v_1056;
assign x_17842 = v_2727 | ~v_182;
assign x_17843 = v_2727 | ~v_163;
assign x_17844 = v_2727 | ~v_162;
assign x_17845 = v_2727 | ~v_155;
assign x_17846 = v_2727 | ~v_137;
assign x_17847 = v_2727 | ~v_136;
assign x_17848 = v_2727 | ~v_135;
assign x_17849 = v_2727 | ~v_134;
assign x_17850 = v_2727 | ~v_18;
assign x_17851 = v_2727 | ~v_17;
assign x_17852 = v_2727 | ~v_15;
assign x_17853 = v_2727 | ~v_8;
assign x_17854 = ~v_2725 | ~v_2724 | ~v_2723 | v_2726;
assign x_17855 = v_2725 | ~v_2681;
assign x_17856 = v_2725 | ~v_2682;
assign x_17857 = v_2725 | ~v_2683;
assign x_17858 = v_2725 | ~v_2684;
assign x_17859 = v_2725 | ~v_1694;
assign x_17860 = v_2725 | ~v_1695;
assign x_17861 = v_2725 | ~v_1696;
assign x_17862 = v_2725 | ~v_1697;
assign x_17863 = v_2725 | ~v_1636;
assign x_17864 = v_2725 | ~v_1637;
assign x_17865 = v_2725 | ~v_1638;
assign x_17866 = v_2725 | ~v_1639;
assign x_17867 = v_2725 | ~v_1640;
assign x_17868 = v_2725 | ~v_1641;
assign x_17869 = v_2725 | ~v_2125;
assign x_17870 = v_2725 | ~v_2126;
assign x_17871 = v_2725 | ~v_2127;
assign x_17872 = v_2725 | ~v_2128;
assign x_17873 = v_2725 | ~v_2075;
assign x_17874 = v_2725 | ~v_2076;
assign x_17875 = v_2725 | ~v_2077;
assign x_17876 = v_2725 | ~v_2078;
assign x_17877 = v_2725 | ~v_2079;
assign x_17878 = v_2725 | ~v_2080;
assign x_17879 = v_2725 | ~v_1037;
assign x_17880 = v_2725 | ~v_1038;
assign x_17881 = v_2725 | ~v_1039;
assign x_17882 = v_2725 | ~v_1040;
assign x_17883 = v_2725 | ~v_927;
assign x_17884 = v_2725 | ~v_928;
assign x_17885 = v_2725 | ~v_839;
assign x_17886 = v_2725 | ~v_840;
assign x_17887 = v_2725 | ~v_184;
assign x_17888 = v_2725 | ~v_170;
assign x_17889 = v_2725 | ~v_169;
assign x_17890 = v_2725 | ~v_151;
assign x_17891 = v_2725 | ~v_150;
assign x_17892 = v_2725 | ~v_149;
assign x_17893 = v_2725 | ~v_147;
assign x_17894 = v_2725 | ~v_103;
assign x_17895 = v_2725 | ~v_101;
assign x_17896 = v_2725 | ~v_100;
assign x_17897 = v_2725 | ~v_98;
assign x_17898 = v_2725 | ~v_96;
assign x_17899 = v_2724 | ~v_2676;
assign x_17900 = v_2724 | ~v_2677;
assign x_17901 = v_2724 | ~v_2678;
assign x_17902 = v_2724 | ~v_2679;
assign x_17903 = v_2724 | ~v_1685;
assign x_17904 = v_2724 | ~v_1686;
assign x_17905 = v_2724 | ~v_1687;
assign x_17906 = v_2724 | ~v_1688;
assign x_17907 = v_2724 | ~v_1611;
assign x_17908 = v_2724 | ~v_1612;
assign x_17909 = v_2724 | ~v_1613;
assign x_17910 = v_2724 | ~v_1614;
assign x_17911 = v_2724 | ~v_1615;
assign x_17912 = v_2724 | ~v_1616;
assign x_17913 = v_2724 | ~v_2120;
assign x_17914 = v_2724 | ~v_2121;
assign x_17915 = v_2724 | ~v_2122;
assign x_17916 = v_2724 | ~v_2123;
assign x_17917 = v_2724 | ~v_2060;
assign x_17918 = v_2724 | ~v_2061;
assign x_17919 = v_2724 | ~v_2062;
assign x_17920 = v_2724 | ~v_2063;
assign x_17921 = v_2724 | ~v_2064;
assign x_17922 = v_2724 | ~v_2065;
assign x_17923 = v_2724 | ~v_1032;
assign x_17924 = v_2724 | ~v_1033;
assign x_17925 = v_2724 | ~v_1034;
assign x_17926 = v_2724 | ~v_1035;
assign x_17927 = v_2724 | ~v_912;
assign x_17928 = v_2724 | ~v_913;
assign x_17929 = v_2724 | ~v_806;
assign x_17930 = v_2724 | ~v_807;
assign x_17931 = v_2724 | ~v_183;
assign x_17932 = v_2724 | ~v_166;
assign x_17933 = v_2724 | ~v_165;
assign x_17934 = v_2724 | ~v_146;
assign x_17935 = v_2724 | ~v_145;
assign x_17936 = v_2724 | ~v_144;
assign x_17937 = v_2724 | ~v_142;
assign x_17938 = v_2724 | ~v_61;
assign x_17939 = v_2724 | ~v_59;
assign x_17940 = v_2724 | ~v_58;
assign x_17941 = v_2724 | ~v_56;
assign x_17942 = v_2724 | ~v_54;
assign x_17943 = v_2723 | ~v_2671;
assign x_17944 = v_2723 | ~v_2672;
assign x_17945 = v_2723 | ~v_2673;
assign x_17946 = v_2723 | ~v_2674;
assign x_17947 = v_2723 | ~v_1676;
assign x_17948 = v_2723 | ~v_1677;
assign x_17949 = v_2723 | ~v_1678;
assign x_17950 = v_2723 | ~v_1679;
assign x_17951 = v_2723 | ~v_1586;
assign x_17952 = v_2723 | ~v_1587;
assign x_17953 = v_2723 | ~v_1588;
assign x_17954 = v_2723 | ~v_1589;
assign x_17955 = v_2723 | ~v_1590;
assign x_17956 = v_2723 | ~v_1591;
assign x_17957 = v_2723 | ~v_2115;
assign x_17958 = v_2723 | ~v_2116;
assign x_17959 = v_2723 | ~v_2117;
assign x_17960 = v_2723 | ~v_2118;
assign x_17961 = v_2723 | ~v_2045;
assign x_17962 = v_2723 | ~v_2046;
assign x_17963 = v_2723 | ~v_2047;
assign x_17964 = v_2723 | ~v_2048;
assign x_17965 = v_2723 | ~v_2049;
assign x_17966 = v_2723 | ~v_2050;
assign x_17967 = v_2723 | ~v_1027;
assign x_17968 = v_2723 | ~v_1028;
assign x_17969 = v_2723 | ~v_1029;
assign x_17970 = v_2723 | ~v_1030;
assign x_17971 = v_2723 | ~v_897;
assign x_17972 = v_2723 | ~v_898;
assign x_17973 = v_2723 | ~v_773;
assign x_17974 = v_2723 | ~v_774;
assign x_17975 = v_2723 | ~v_182;
assign x_17976 = v_2723 | ~v_162;
assign x_17977 = v_2723 | ~v_161;
assign x_17978 = v_2723 | ~v_138;
assign x_17979 = v_2723 | ~v_137;
assign x_17980 = v_2723 | ~v_136;
assign x_17981 = v_2723 | ~v_134;
assign x_17982 = v_2723 | ~v_18;
assign x_17983 = v_2723 | ~v_16;
assign x_17984 = v_2723 | ~v_15;
assign x_17985 = v_2723 | ~v_13;
assign x_17986 = v_2723 | ~v_11;
assign x_17987 = ~v_2721 | ~v_2720 | ~v_2719 | v_2722;
assign x_17988 = v_2721 | ~v_2681;
assign x_17989 = v_2721 | ~v_2682;
assign x_17990 = v_2721 | ~v_2683;
assign x_17991 = v_2721 | ~v_2684;
assign x_17992 = v_2721 | ~v_1666;
assign x_17993 = v_2721 | ~v_1667;
assign x_17994 = v_2721 | ~v_1668;
assign x_17995 = v_2721 | ~v_1669;
assign x_17996 = v_2721 | ~v_1636;
assign x_17997 = v_2721 | ~v_1750;
assign x_17998 = v_2721 | ~v_1751;
assign x_17999 = v_2721 | ~v_1639;
assign x_18000 = v_2721 | ~v_1752;
assign x_18001 = v_2721 | ~v_1753;
assign x_18002 = v_2721 | ~v_2161;
assign x_18003 = v_2721 | ~v_2162;
assign x_18004 = v_2721 | ~v_2163;
assign x_18005 = v_2721 | ~v_2164;
assign x_18006 = v_2721 | ~v_2075;
assign x_18007 = v_2721 | ~v_2141;
assign x_18008 = v_2721 | ~v_2142;
assign x_18009 = v_2721 | ~v_2078;
assign x_18010 = v_2721 | ~v_2143;
assign x_18011 = v_2721 | ~v_2144;
assign x_18012 = v_2721 | ~v_1193;
assign x_18013 = v_2721 | ~v_1241;
assign x_18014 = v_2721 | ~v_1194;
assign x_18015 = v_2721 | ~v_1242;
assign x_18016 = v_2721 | ~v_1023;
assign x_18017 = v_2721 | ~v_1024;
assign x_18018 = v_2721 | ~v_1243;
assign x_18019 = v_2721 | ~v_1244;
assign x_18020 = v_2721 | ~v_184;
assign x_18021 = v_2721 | ~v_171;
assign x_18022 = v_2721 | ~v_169;
assign x_18023 = v_2721 | ~v_149;
assign x_18024 = v_2721 | ~v_148;
assign x_18025 = v_2721 | ~v_147;
assign x_18026 = v_2721 | ~v_103;
assign x_18027 = v_2721 | ~v_102;
assign x_18028 = v_2721 | ~v_101;
assign x_18029 = v_2721 | ~v_100;
assign x_18030 = v_2721 | ~v_99;
assign x_18031 = v_2721 | ~v_94;
assign x_18032 = v_2720 | ~v_2676;
assign x_18033 = v_2720 | ~v_2677;
assign x_18034 = v_2720 | ~v_2678;
assign x_18035 = v_2720 | ~v_2679;
assign x_18036 = v_2720 | ~v_1657;
assign x_18037 = v_2720 | ~v_1658;
assign x_18038 = v_2720 | ~v_1659;
assign x_18039 = v_2720 | ~v_1660;
assign x_18040 = v_2720 | ~v_1611;
assign x_18041 = v_2720 | ~v_1741;
assign x_18042 = v_2720 | ~v_1742;
assign x_18043 = v_2720 | ~v_1614;
assign x_18044 = v_2720 | ~v_1743;
assign x_18045 = v_2720 | ~v_1744;
assign x_18046 = v_2720 | ~v_2156;
assign x_18047 = v_2720 | ~v_2157;
assign x_18048 = v_2720 | ~v_2158;
assign x_18049 = v_2720 | ~v_2159;
assign x_18050 = v_2720 | ~v_2060;
assign x_18051 = v_2720 | ~v_2136;
assign x_18052 = v_2720 | ~v_2137;
assign x_18053 = v_2720 | ~v_2063;
assign x_18054 = v_2720 | ~v_2138;
assign x_18055 = v_2720 | ~v_2139;
assign x_18056 = v_2720 | ~v_1178;
assign x_18057 = v_2720 | ~v_1236;
assign x_18058 = v_2720 | ~v_1179;
assign x_18059 = v_2720 | ~v_1237;
assign x_18060 = v_2720 | ~v_1008;
assign x_18061 = v_2720 | ~v_1009;
assign x_18062 = v_2720 | ~v_1238;
assign x_18063 = v_2720 | ~v_1239;
assign x_18064 = v_2720 | ~v_183;
assign x_18065 = v_2720 | ~v_167;
assign x_18066 = v_2720 | ~v_165;
assign x_18067 = v_2720 | ~v_144;
assign x_18068 = v_2720 | ~v_143;
assign x_18069 = v_2720 | ~v_142;
assign x_18070 = v_2720 | ~v_61;
assign x_18071 = v_2720 | ~v_60;
assign x_18072 = v_2720 | ~v_59;
assign x_18073 = v_2720 | ~v_58;
assign x_18074 = v_2720 | ~v_57;
assign x_18075 = v_2720 | ~v_52;
assign x_18076 = v_2719 | ~v_2671;
assign x_18077 = v_2719 | ~v_2672;
assign x_18078 = v_2719 | ~v_2673;
assign x_18079 = v_2719 | ~v_2674;
assign x_18080 = v_2719 | ~v_1648;
assign x_18081 = v_2719 | ~v_1649;
assign x_18082 = v_2719 | ~v_1650;
assign x_18083 = v_2719 | ~v_1651;
assign x_18084 = v_2719 | ~v_1586;
assign x_18085 = v_2719 | ~v_1732;
assign x_18086 = v_2719 | ~v_1733;
assign x_18087 = v_2719 | ~v_1589;
assign x_18088 = v_2719 | ~v_1734;
assign x_18089 = v_2719 | ~v_1735;
assign x_18090 = v_2719 | ~v_2151;
assign x_18091 = v_2719 | ~v_2152;
assign x_18092 = v_2719 | ~v_2153;
assign x_18093 = v_2719 | ~v_2154;
assign x_18094 = v_2719 | ~v_2045;
assign x_18095 = v_2719 | ~v_2131;
assign x_18096 = v_2719 | ~v_2132;
assign x_18097 = v_2719 | ~v_2048;
assign x_18098 = v_2719 | ~v_2133;
assign x_18099 = v_2719 | ~v_2134;
assign x_18100 = v_2719 | ~v_1163;
assign x_18101 = v_2719 | ~v_1231;
assign x_18102 = v_2719 | ~v_1164;
assign x_18103 = v_2719 | ~v_1232;
assign x_18104 = v_2719 | ~v_1233;
assign x_18105 = v_2719 | ~v_1234;
assign x_18106 = v_2719 | ~v_182;
assign x_18107 = v_2719 | ~v_163;
assign x_18108 = v_2719 | ~v_161;
assign x_18109 = v_2719 | ~v_136;
assign x_18110 = v_2719 | ~v_135;
assign x_18111 = v_2719 | ~v_134;
assign x_18112 = v_2719 | ~v_993;
assign x_18113 = v_2719 | ~v_994;
assign x_18114 = v_2719 | ~v_18;
assign x_18115 = v_2719 | ~v_17;
assign x_18116 = v_2719 | ~v_16;
assign x_18117 = v_2719 | ~v_15;
assign x_18118 = v_2719 | ~v_14;
assign x_18119 = v_2719 | ~v_9;
assign x_18120 = ~v_2717 | ~v_2716 | ~v_2715 | v_2718;
assign x_18121 = v_2717 | ~v_2681;
assign x_18122 = v_2717 | ~v_2682;
assign x_18123 = v_2717 | ~v_2683;
assign x_18124 = v_2717 | ~v_2684;
assign x_18125 = v_2717 | ~v_1694;
assign x_18126 = v_2717 | ~v_1695;
assign x_18127 = v_2717 | ~v_1696;
assign x_18128 = v_2717 | ~v_1697;
assign x_18129 = v_2717 | ~v_1666;
assign x_18130 = v_2717 | ~v_1667;
assign x_18131 = v_2717 | ~v_1668;
assign x_18132 = v_2717 | ~v_1669;
assign x_18133 = v_2717 | ~v_1636;
assign x_18134 = v_2717 | ~v_1639;
assign x_18135 = v_2717 | ~v_2161;
assign x_18136 = v_2717 | ~v_2162;
assign x_18137 = v_2717 | ~v_2163;
assign x_18138 = v_2717 | ~v_2164;
assign x_18139 = v_2717 | ~v_2125;
assign x_18140 = v_2717 | ~v_2126;
assign x_18141 = v_2717 | ~v_2127;
assign x_18142 = v_2717 | ~v_2128;
assign x_18143 = v_2717 | ~v_2075;
assign x_18144 = v_2717 | ~v_2078;
assign x_18145 = v_2717 | ~v_1209;
assign x_18146 = v_2717 | ~v_1210;
assign x_18147 = v_2717 | ~v_1193;
assign x_18148 = v_2717 | ~v_1194;
assign x_18149 = v_2717 | ~v_927;
assign x_18150 = v_2717 | ~v_928;
assign x_18151 = v_2717 | ~v_1211;
assign x_18152 = v_2717 | ~v_1212;
assign x_18153 = v_2717 | ~v_184;
assign x_18154 = v_2717 | ~v_172;
assign x_18155 = v_2717 | ~v_171;
assign x_18156 = v_2717 | ~v_169;
assign x_18157 = v_2717 | ~v_150;
assign x_18158 = v_2717 | ~v_149;
assign x_18159 = v_2717 | ~v_147;
assign x_18160 = v_2717 | ~v_102;
assign x_18161 = v_2717 | ~v_101;
assign x_18162 = v_2717 | ~v_100;
assign x_18163 = v_2717 | ~v_96;
assign x_18164 = v_2717 | ~v_94;
assign x_18165 = v_2716 | ~v_2676;
assign x_18166 = v_2716 | ~v_2677;
assign x_18167 = v_2716 | ~v_2678;
assign x_18168 = v_2716 | ~v_2679;
assign x_18169 = v_2716 | ~v_1685;
assign x_18170 = v_2716 | ~v_1686;
assign x_18171 = v_2716 | ~v_1687;
assign x_18172 = v_2716 | ~v_1688;
assign x_18173 = v_2716 | ~v_1657;
assign x_18174 = v_2716 | ~v_1658;
assign x_18175 = v_2716 | ~v_1659;
assign x_18176 = v_2716 | ~v_1660;
assign x_18177 = v_2716 | ~v_1611;
assign x_18178 = v_2716 | ~v_1614;
assign x_18179 = v_2716 | ~v_2156;
assign x_18180 = v_2716 | ~v_2157;
assign x_18181 = v_2716 | ~v_2158;
assign x_18182 = v_2716 | ~v_2159;
assign x_18183 = v_2716 | ~v_2120;
assign x_18184 = v_2716 | ~v_2121;
assign x_18185 = v_2716 | ~v_2122;
assign x_18186 = v_2716 | ~v_2123;
assign x_18187 = v_2716 | ~v_2060;
assign x_18188 = v_2716 | ~v_2063;
assign x_18189 = v_2716 | ~v_1204;
assign x_18190 = v_2716 | ~v_1205;
assign x_18191 = v_2716 | ~v_1178;
assign x_18192 = v_2716 | ~v_1179;
assign x_18193 = v_2716 | ~v_912;
assign x_18194 = v_2716 | ~v_913;
assign x_18195 = v_2716 | ~v_1206;
assign x_18196 = v_2716 | ~v_1207;
assign x_18197 = v_2716 | ~v_183;
assign x_18198 = v_2716 | ~v_168;
assign x_18199 = v_2716 | ~v_167;
assign x_18200 = v_2716 | ~v_165;
assign x_18201 = v_2716 | ~v_145;
assign x_18202 = v_2716 | ~v_144;
assign x_18203 = v_2716 | ~v_142;
assign x_18204 = v_2716 | ~v_60;
assign x_18205 = v_2716 | ~v_59;
assign x_18206 = v_2716 | ~v_58;
assign x_18207 = v_2716 | ~v_54;
assign x_18208 = v_2716 | ~v_52;
assign x_18209 = v_2715 | ~v_2671;
assign x_18210 = v_2715 | ~v_2672;
assign x_18211 = v_2715 | ~v_2673;
assign x_18212 = v_2715 | ~v_2674;
assign x_18213 = v_2715 | ~v_1676;
assign x_18214 = v_2715 | ~v_1677;
assign x_18215 = v_2715 | ~v_1678;
assign x_18216 = v_2715 | ~v_1679;
assign x_18217 = v_2715 | ~v_1648;
assign x_18218 = v_2715 | ~v_1649;
assign x_18219 = v_2715 | ~v_1650;
assign x_18220 = v_2715 | ~v_1651;
assign x_18221 = v_2715 | ~v_1586;
assign x_18222 = v_2715 | ~v_1589;
assign x_18223 = v_2715 | ~v_2151;
assign x_18224 = v_2715 | ~v_2152;
assign x_18225 = v_2715 | ~v_2153;
assign x_18226 = v_2715 | ~v_2154;
assign x_18227 = v_2715 | ~v_2115;
assign x_18228 = v_2715 | ~v_2116;
assign x_18229 = v_2715 | ~v_2117;
assign x_18230 = v_2715 | ~v_2118;
assign x_18231 = v_2715 | ~v_2045;
assign x_18232 = v_2715 | ~v_2048;
assign x_18233 = v_2715 | ~v_1199;
assign x_18234 = v_2715 | ~v_1200;
assign x_18235 = v_2715 | ~v_1163;
assign x_18236 = v_2715 | ~v_1164;
assign x_18237 = v_2715 | ~v_897;
assign x_18238 = v_2715 | ~v_898;
assign x_18239 = v_2715 | ~v_1201;
assign x_18240 = v_2715 | ~v_1202;
assign x_18241 = v_2715 | ~v_182;
assign x_18242 = v_2715 | ~v_164;
assign x_18243 = v_2715 | ~v_163;
assign x_18244 = v_2715 | ~v_161;
assign x_18245 = v_2715 | ~v_137;
assign x_18246 = v_2715 | ~v_136;
assign x_18247 = v_2715 | ~v_134;
assign x_18248 = v_2715 | ~v_17;
assign x_18249 = v_2715 | ~v_16;
assign x_18250 = v_2715 | ~v_15;
assign x_18251 = v_2715 | ~v_11;
assign x_18252 = v_2715 | ~v_9;
assign x_18253 = ~v_2713 | ~v_2712 | ~v_2711 | v_2714;
assign x_18254 = v_2713 | ~v_2681;
assign x_18255 = v_2713 | ~v_2682;
assign x_18256 = v_2713 | ~v_2683;
assign x_18257 = v_2713 | ~v_2684;
assign x_18258 = v_2713 | ~v_1632;
assign x_18259 = v_2713 | ~v_1633;
assign x_18260 = v_2713 | ~v_1634;
assign x_18261 = v_2713 | ~v_1635;
assign x_18262 = v_2713 | ~v_1666;
assign x_18263 = v_2713 | ~v_1667;
assign x_18264 = v_2713 | ~v_1668;
assign x_18265 = v_2713 | ~v_1669;
assign x_18266 = v_2713 | ~v_1636;
assign x_18267 = v_2713 | ~v_1639;
assign x_18268 = v_2713 | ~v_2161;
assign x_18269 = v_2713 | ~v_2162;
assign x_18270 = v_2713 | ~v_2163;
assign x_18271 = v_2713 | ~v_2164;
assign x_18272 = v_2713 | ~v_2109;
assign x_18273 = v_2713 | ~v_2110;
assign x_18274 = v_2713 | ~v_2111;
assign x_18275 = v_2713 | ~v_2112;
assign x_18276 = v_2713 | ~v_2075;
assign x_18277 = v_2713 | ~v_2078;
assign x_18278 = v_2713 | ~v_1225;
assign x_18279 = v_2713 | ~v_1226;
assign x_18280 = v_2713 | ~v_1227;
assign x_18281 = v_2713 | ~v_1228;
assign x_18282 = v_2713 | ~v_1193;
assign x_18283 = v_2713 | ~v_1194;
assign x_18284 = v_2713 | ~v_975;
assign x_18285 = v_2713 | ~v_976;
assign x_18286 = v_2713 | ~v_184;
assign x_18287 = v_2713 | ~v_171;
assign x_18288 = v_2713 | ~v_169;
assign x_18289 = v_2713 | ~v_150;
assign x_18290 = v_2713 | ~v_148;
assign x_18291 = v_2713 | ~v_103;
assign x_18292 = v_2713 | ~v_102;
assign x_18293 = v_2713 | ~v_101;
assign x_18294 = v_2713 | ~v_100;
assign x_18295 = v_2713 | ~v_97;
assign x_18296 = v_2713 | ~v_95;
assign x_18297 = v_2713 | ~v_94;
assign x_18298 = v_2712 | ~v_2676;
assign x_18299 = v_2712 | ~v_2677;
assign x_18300 = v_2712 | ~v_2678;
assign x_18301 = v_2712 | ~v_2679;
assign x_18302 = v_2712 | ~v_1607;
assign x_18303 = v_2712 | ~v_1608;
assign x_18304 = v_2712 | ~v_1609;
assign x_18305 = v_2712 | ~v_1610;
assign x_18306 = v_2712 | ~v_1657;
assign x_18307 = v_2712 | ~v_1658;
assign x_18308 = v_2712 | ~v_1659;
assign x_18309 = v_2712 | ~v_1660;
assign x_18310 = v_2712 | ~v_1611;
assign x_18311 = v_2712 | ~v_1614;
assign x_18312 = v_2712 | ~v_2156;
assign x_18313 = v_2712 | ~v_2157;
assign x_18314 = v_2712 | ~v_2158;
assign x_18315 = v_2712 | ~v_2159;
assign x_18316 = v_2712 | ~v_2104;
assign x_18317 = v_2712 | ~v_2105;
assign x_18318 = v_2712 | ~v_2106;
assign x_18319 = v_2712 | ~v_2107;
assign x_18320 = v_2712 | ~v_2060;
assign x_18321 = v_2712 | ~v_2063;
assign x_18322 = v_2712 | ~v_1220;
assign x_18323 = v_2712 | ~v_1221;
assign x_18324 = v_2712 | ~v_1222;
assign x_18325 = v_2712 | ~v_1223;
assign x_18326 = v_2712 | ~v_1178;
assign x_18327 = v_2712 | ~v_1179;
assign x_18328 = v_2712 | ~v_960;
assign x_18329 = v_2712 | ~v_961;
assign x_18330 = v_2712 | ~v_183;
assign x_18331 = v_2712 | ~v_167;
assign x_18332 = v_2712 | ~v_165;
assign x_18333 = v_2712 | ~v_145;
assign x_18334 = v_2712 | ~v_143;
assign x_18335 = v_2712 | ~v_61;
assign x_18336 = v_2712 | ~v_60;
assign x_18337 = v_2712 | ~v_59;
assign x_18338 = v_2712 | ~v_58;
assign x_18339 = v_2712 | ~v_55;
assign x_18340 = v_2712 | ~v_53;
assign x_18341 = v_2712 | ~v_52;
assign x_18342 = v_2711 | ~v_2671;
assign x_18343 = v_2711 | ~v_2672;
assign x_18344 = v_2711 | ~v_2673;
assign x_18345 = v_2711 | ~v_2674;
assign x_18346 = v_2711 | ~v_1582;
assign x_18347 = v_2711 | ~v_1583;
assign x_18348 = v_2711 | ~v_1584;
assign x_18349 = v_2711 | ~v_1585;
assign x_18350 = v_2711 | ~v_1648;
assign x_18351 = v_2711 | ~v_1649;
assign x_18352 = v_2711 | ~v_1650;
assign x_18353 = v_2711 | ~v_1651;
assign x_18354 = v_2711 | ~v_1586;
assign x_18355 = v_2711 | ~v_1589;
assign x_18356 = v_2711 | ~v_2151;
assign x_18357 = v_2711 | ~v_2152;
assign x_18358 = v_2711 | ~v_2153;
assign x_18359 = v_2711 | ~v_2154;
assign x_18360 = v_2711 | ~v_2099;
assign x_18361 = v_2711 | ~v_2100;
assign x_18362 = v_2711 | ~v_2101;
assign x_18363 = v_2711 | ~v_2102;
assign x_18364 = v_2711 | ~v_2045;
assign x_18365 = v_2711 | ~v_2048;
assign x_18366 = v_2711 | ~v_1215;
assign x_18367 = v_2711 | ~v_1216;
assign x_18368 = v_2711 | ~v_1217;
assign x_18369 = v_2711 | ~v_1218;
assign x_18370 = v_2711 | ~v_1163;
assign x_18371 = v_2711 | ~v_1164;
assign x_18372 = v_2711 | ~v_945;
assign x_18373 = v_2711 | ~v_946;
assign x_18374 = v_2711 | ~v_182;
assign x_18375 = v_2711 | ~v_163;
assign x_18376 = v_2711 | ~v_161;
assign x_18377 = v_2711 | ~v_137;
assign x_18378 = v_2711 | ~v_135;
assign x_18379 = v_2711 | ~v_18;
assign x_18380 = v_2711 | ~v_17;
assign x_18381 = v_2711 | ~v_16;
assign x_18382 = v_2711 | ~v_15;
assign x_18383 = v_2711 | ~v_12;
assign x_18384 = v_2711 | ~v_10;
assign x_18385 = v_2711 | ~v_9;
assign x_18386 = ~v_2709 | ~v_2708 | ~v_2707 | v_2710;
assign x_18387 = v_2709 | ~v_2681;
assign x_18388 = v_2709 | ~v_2682;
assign x_18389 = v_2709 | ~v_2683;
assign x_18390 = v_2709 | ~v_2684;
assign x_18391 = v_2709 | ~v_1722;
assign x_18392 = v_2709 | ~v_1723;
assign x_18393 = v_2709 | ~v_1724;
assign x_18394 = v_2709 | ~v_1725;
assign x_18395 = v_2709 | ~v_1666;
assign x_18396 = v_2709 | ~v_1667;
assign x_18397 = v_2709 | ~v_1668;
assign x_18398 = v_2709 | ~v_1669;
assign x_18399 = v_2709 | ~v_1636;
assign x_18400 = v_2709 | ~v_1639;
assign x_18401 = v_2709 | ~v_2161;
assign x_18402 = v_2709 | ~v_2162;
assign x_18403 = v_2709 | ~v_2163;
assign x_18404 = v_2709 | ~v_2164;
assign x_18405 = v_2709 | ~v_2071;
assign x_18406 = v_2709 | ~v_2072;
assign x_18407 = v_2709 | ~v_2073;
assign x_18408 = v_2709 | ~v_2074;
assign x_18409 = v_2709 | ~v_2075;
assign x_18410 = v_2709 | ~v_2078;
assign x_18411 = v_2709 | ~v_1191;
assign x_18412 = v_2709 | ~v_1192;
assign x_18413 = v_2709 | ~v_1193;
assign x_18414 = v_2709 | ~v_1194;
assign x_18415 = v_2709 | ~v_837;
assign x_18416 = v_2709 | ~v_838;
assign x_18417 = v_2709 | ~v_1195;
assign x_18418 = v_2709 | ~v_1196;
assign x_18419 = v_2709 | ~v_184;
assign x_18420 = v_2709 | ~v_171;
assign x_18421 = v_2709 | ~v_169;
assign x_18422 = v_2709 | ~v_160;
assign x_18423 = v_2709 | ~v_151;
assign x_18424 = v_2709 | ~v_150;
assign x_18425 = v_2709 | ~v_149;
assign x_18426 = v_2709 | ~v_148;
assign x_18427 = v_2709 | ~v_147;
assign x_18428 = v_2709 | ~v_103;
assign x_18429 = v_2709 | ~v_100;
assign x_18430 = v_2709 | ~v_94;
assign x_18431 = v_2708 | ~v_2676;
assign x_18432 = v_2708 | ~v_2677;
assign x_18433 = v_2708 | ~v_2678;
assign x_18434 = v_2708 | ~v_2679;
assign x_18435 = v_2708 | ~v_1713;
assign x_18436 = v_2708 | ~v_1714;
assign x_18437 = v_2708 | ~v_1715;
assign x_18438 = v_2708 | ~v_1716;
assign x_18439 = v_2708 | ~v_1657;
assign x_18440 = v_2708 | ~v_1658;
assign x_18441 = v_2708 | ~v_1659;
assign x_18442 = v_2708 | ~v_1660;
assign x_18443 = v_2708 | ~v_1611;
assign x_18444 = v_2708 | ~v_1614;
assign x_18445 = v_2708 | ~v_2156;
assign x_18446 = v_2708 | ~v_2157;
assign x_18447 = v_2708 | ~v_2158;
assign x_18448 = v_2708 | ~v_2159;
assign x_18449 = v_2708 | ~v_2056;
assign x_18450 = v_2708 | ~v_2057;
assign x_18451 = v_2708 | ~v_2058;
assign x_18452 = v_2708 | ~v_2059;
assign x_18453 = v_2708 | ~v_2060;
assign x_18454 = v_2708 | ~v_2063;
assign x_18455 = v_2708 | ~v_1176;
assign x_18456 = v_2708 | ~v_1177;
assign x_18457 = v_2708 | ~v_1178;
assign x_18458 = v_2708 | ~v_1179;
assign x_18459 = v_2708 | ~v_804;
assign x_18460 = v_2708 | ~v_805;
assign x_18461 = v_2708 | ~v_1180;
assign x_18462 = v_2708 | ~v_1181;
assign x_18463 = v_2708 | ~v_183;
assign x_18464 = v_2708 | ~v_167;
assign x_18465 = v_2708 | ~v_165;
assign x_18466 = v_2708 | ~v_159;
assign x_18467 = v_2708 | ~v_146;
assign x_18468 = v_2708 | ~v_145;
assign x_18469 = v_2708 | ~v_144;
assign x_18470 = v_2708 | ~v_143;
assign x_18471 = v_2708 | ~v_142;
assign x_18472 = v_2708 | ~v_61;
assign x_18473 = v_2708 | ~v_58;
assign x_18474 = v_2708 | ~v_52;
assign x_18475 = v_2707 | ~v_2671;
assign x_18476 = v_2707 | ~v_2672;
assign x_18477 = v_2707 | ~v_2673;
assign x_18478 = v_2707 | ~v_2674;
assign x_18479 = v_2707 | ~v_1704;
assign x_18480 = v_2707 | ~v_1705;
assign x_18481 = v_2707 | ~v_1706;
assign x_18482 = v_2707 | ~v_1707;
assign x_18483 = v_2707 | ~v_1648;
assign x_18484 = v_2707 | ~v_1649;
assign x_18485 = v_2707 | ~v_1650;
assign x_18486 = v_2707 | ~v_1651;
assign x_18487 = v_2707 | ~v_1586;
assign x_18488 = v_2707 | ~v_1589;
assign x_18489 = v_2707 | ~v_2151;
assign x_18490 = v_2707 | ~v_2152;
assign x_18491 = v_2707 | ~v_2153;
assign x_18492 = v_2707 | ~v_2154;
assign x_18493 = v_2707 | ~v_2041;
assign x_18494 = v_2707 | ~v_2042;
assign x_18495 = v_2707 | ~v_2043;
assign x_18496 = v_2707 | ~v_2044;
assign x_18497 = v_2707 | ~v_2045;
assign x_18498 = v_2707 | ~v_2048;
assign x_18499 = v_2707 | ~v_1161;
assign x_18500 = v_2707 | ~v_1162;
assign x_18501 = v_2707 | ~v_1163;
assign x_18502 = v_2707 | ~v_1164;
assign x_18503 = v_2707 | ~v_771;
assign x_18504 = v_2707 | ~v_772;
assign x_18505 = v_2707 | ~v_1165;
assign x_18506 = v_2707 | ~v_1166;
assign x_18507 = v_2707 | ~v_182;
assign x_18508 = v_2707 | ~v_163;
assign x_18509 = v_2707 | ~v_161;
assign x_18510 = v_2707 | ~v_155;
assign x_18511 = v_2707 | ~v_138;
assign x_18512 = v_2707 | ~v_137;
assign x_18513 = v_2707 | ~v_136;
assign x_18514 = v_2707 | ~v_135;
assign x_18515 = v_2707 | ~v_134;
assign x_18516 = v_2707 | ~v_18;
assign x_18517 = v_2707 | ~v_15;
assign x_18518 = v_2707 | ~v_9;
assign x_18519 = ~v_2705 | ~v_2704 | ~v_2703 | v_2706;
assign x_18520 = v_2705 | ~v_2681;
assign x_18521 = v_2705 | ~v_2682;
assign x_18522 = v_2705 | ~v_2683;
assign x_18523 = v_2705 | ~v_2684;
assign x_18524 = v_2705 | ~v_1632;
assign x_18525 = v_2705 | ~v_1633;
assign x_18526 = v_2705 | ~v_1634;
assign x_18527 = v_2705 | ~v_1635;
assign x_18528 = v_2705 | ~v_1636;
assign x_18529 = v_2705 | ~v_1637;
assign x_18530 = v_2705 | ~v_1638;
assign x_18531 = v_2705 | ~v_1639;
assign x_18532 = v_2705 | ~v_1640;
assign x_18533 = v_2705 | ~v_1641;
assign x_18534 = v_2705 | ~v_2109;
assign x_18535 = v_2705 | ~v_2110;
assign x_18536 = v_2705 | ~v_2111;
assign x_18537 = v_2705 | ~v_2112;
assign x_18538 = v_2705 | ~v_2075;
assign x_18539 = v_2705 | ~v_2076;
assign x_18540 = v_2705 | ~v_2077;
assign x_18541 = v_2705 | ~v_2078;
assign x_18542 = v_2705 | ~v_2079;
assign x_18543 = v_2705 | ~v_2080;
assign x_18544 = v_2705 | ~v_1147;
assign x_18545 = v_2705 | ~v_1148;
assign x_18546 = v_2705 | ~v_975;
assign x_18547 = v_2705 | ~v_976;
assign x_18548 = v_2705 | ~v_839;
assign x_18549 = v_2705 | ~v_840;
assign x_18550 = v_2705 | ~v_1149;
assign x_18551 = v_2705 | ~v_1150;
assign x_18552 = v_2705 | ~v_184;
assign x_18553 = v_2705 | ~v_170;
assign x_18554 = v_2705 | ~v_169;
assign x_18555 = v_2705 | ~v_150;
assign x_18556 = v_2705 | ~v_148;
assign x_18557 = v_2705 | ~v_147;
assign x_18558 = v_2705 | ~v_103;
assign x_18559 = v_2705 | ~v_102;
assign x_18560 = v_2705 | ~v_101;
assign x_18561 = v_2705 | ~v_100;
assign x_18562 = v_2705 | ~v_98;
assign x_18563 = v_2705 | ~v_97;
assign x_18564 = v_2704 | ~v_2676;
assign x_18565 = v_2704 | ~v_2677;
assign x_18566 = v_2704 | ~v_2678;
assign x_18567 = v_2704 | ~v_2679;
assign x_18568 = v_2704 | ~v_1607;
assign x_18569 = v_2704 | ~v_1608;
assign x_18570 = v_2704 | ~v_1609;
assign x_18571 = v_2704 | ~v_1610;
assign x_18572 = v_2704 | ~v_1611;
assign x_18573 = v_2704 | ~v_1612;
assign x_18574 = v_2704 | ~v_1613;
assign x_18575 = v_2704 | ~v_1614;
assign x_18576 = v_2704 | ~v_1615;
assign x_18577 = v_2704 | ~v_1616;
assign x_18578 = v_2704 | ~v_2104;
assign x_18579 = v_2704 | ~v_2105;
assign x_18580 = v_2704 | ~v_2106;
assign x_18581 = v_2704 | ~v_2107;
assign x_18582 = v_2704 | ~v_2060;
assign x_18583 = v_2704 | ~v_2061;
assign x_18584 = v_2704 | ~v_2062;
assign x_18585 = v_2704 | ~v_2063;
assign x_18586 = v_2704 | ~v_2064;
assign x_18587 = v_2704 | ~v_2065;
assign x_18588 = v_2704 | ~v_1142;
assign x_18589 = v_2704 | ~v_1143;
assign x_18590 = v_2704 | ~v_960;
assign x_18591 = v_2704 | ~v_961;
assign x_18592 = v_2704 | ~v_806;
assign x_18593 = v_2704 | ~v_807;
assign x_18594 = v_2704 | ~v_1144;
assign x_18595 = v_2704 | ~v_1145;
assign x_18596 = v_2704 | ~v_183;
assign x_18597 = v_2704 | ~v_166;
assign x_18598 = v_2704 | ~v_165;
assign x_18599 = v_2704 | ~v_145;
assign x_18600 = v_2704 | ~v_143;
assign x_18601 = v_2704 | ~v_142;
assign x_18602 = v_2704 | ~v_61;
assign x_18603 = v_2704 | ~v_60;
assign x_18604 = v_2704 | ~v_59;
assign x_18605 = v_2704 | ~v_58;
assign x_18606 = v_2704 | ~v_56;
assign x_18607 = v_2704 | ~v_55;
assign x_18608 = v_2703 | ~v_2671;
assign x_18609 = v_2703 | ~v_2672;
assign x_18610 = v_2703 | ~v_2673;
assign x_18611 = v_2703 | ~v_2674;
assign x_18612 = v_2703 | ~v_1582;
assign x_18613 = v_2703 | ~v_1583;
assign x_18614 = v_2703 | ~v_1584;
assign x_18615 = v_2703 | ~v_1585;
assign x_18616 = v_2703 | ~v_1586;
assign x_18617 = v_2703 | ~v_1587;
assign x_18618 = v_2703 | ~v_1588;
assign x_18619 = v_2703 | ~v_1589;
assign x_18620 = v_2703 | ~v_1590;
assign x_18621 = v_2703 | ~v_1591;
assign x_18622 = v_2703 | ~v_2099;
assign x_18623 = v_2703 | ~v_2100;
assign x_18624 = v_2703 | ~v_2101;
assign x_18625 = v_2703 | ~v_2102;
assign x_18626 = v_2703 | ~v_2045;
assign x_18627 = v_2703 | ~v_2046;
assign x_18628 = v_2703 | ~v_2047;
assign x_18629 = v_2703 | ~v_2048;
assign x_18630 = v_2703 | ~v_2049;
assign x_18631 = v_2703 | ~v_2050;
assign x_18632 = v_2703 | ~v_1137;
assign x_18633 = v_2703 | ~v_1138;
assign x_18634 = v_2703 | ~v_945;
assign x_18635 = v_2703 | ~v_946;
assign x_18636 = v_2703 | ~v_773;
assign x_18637 = v_2703 | ~v_774;
assign x_18638 = v_2703 | ~v_1139;
assign x_18639 = v_2703 | ~v_1140;
assign x_18640 = v_2703 | ~v_182;
assign x_18641 = v_2703 | ~v_162;
assign x_18642 = v_2703 | ~v_161;
assign x_18643 = v_2703 | ~v_137;
assign x_18644 = v_2703 | ~v_135;
assign x_18645 = v_2703 | ~v_134;
assign x_18646 = v_2703 | ~v_18;
assign x_18647 = v_2703 | ~v_17;
assign x_18648 = v_2703 | ~v_16;
assign x_18649 = v_2703 | ~v_15;
assign x_18650 = v_2703 | ~v_13;
assign x_18651 = v_2703 | ~v_12;
assign x_18652 = ~v_2701 | ~v_2700 | ~v_2699 | v_2702;
assign x_18653 = v_2701 | ~v_2681;
assign x_18654 = v_2701 | ~v_2682;
assign x_18655 = v_2701 | ~v_2683;
assign x_18656 = v_2701 | ~v_2684;
assign x_18657 = v_2701 | ~v_1826;
assign x_18658 = v_2701 | ~v_1827;
assign x_18659 = v_2701 | ~v_1828;
assign x_18660 = v_2701 | ~v_1829;
assign x_18661 = v_2701 | ~v_1636;
assign x_18662 = v_2701 | ~v_1750;
assign x_18663 = v_2701 | ~v_1751;
assign x_18664 = v_2701 | ~v_1639;
assign x_18665 = v_2701 | ~v_1752;
assign x_18666 = v_2701 | ~v_1753;
assign x_18667 = v_2701 | ~v_2093;
assign x_18668 = v_2701 | ~v_2094;
assign x_18669 = v_2701 | ~v_2095;
assign x_18670 = v_2701 | ~v_2096;
assign x_18671 = v_2701 | ~v_2075;
assign x_18672 = v_2701 | ~v_2141;
assign x_18673 = v_2701 | ~v_2142;
assign x_18674 = v_2701 | ~v_2078;
assign x_18675 = v_2701 | ~v_2143;
assign x_18676 = v_2701 | ~v_2144;
assign x_18677 = v_2701 | ~v_885;
assign x_18678 = v_2701 | ~v_1019;
assign x_18679 = v_2701 | ~v_1020;
assign x_18680 = v_2701 | ~v_886;
assign x_18681 = v_2701 | ~v_1021;
assign x_18682 = v_2701 | ~v_1022;
assign x_18683 = v_2701 | ~v_1023;
assign x_18684 = v_2701 | ~v_1024;
assign x_18685 = v_2701 | ~v_184;
assign x_18686 = v_2701 | ~v_181;
assign x_18687 = v_2701 | ~v_171;
assign x_18688 = v_2701 | ~v_170;
assign x_18689 = v_2701 | ~v_169;
assign x_18690 = v_2701 | ~v_149;
assign x_18691 = v_2701 | ~v_148;
assign x_18692 = v_2701 | ~v_147;
assign x_18693 = v_2701 | ~v_103;
assign x_18694 = v_2701 | ~v_102;
assign x_18695 = v_2701 | ~v_101;
assign x_18696 = v_2701 | ~v_99;
assign x_18697 = v_2700 | ~v_2676;
assign x_18698 = v_2700 | ~v_2677;
assign x_18699 = v_2700 | ~v_2678;
assign x_18700 = v_2700 | ~v_2679;
assign x_18701 = v_2700 | ~v_1817;
assign x_18702 = v_2700 | ~v_1818;
assign x_18703 = v_2700 | ~v_1819;
assign x_18704 = v_2700 | ~v_1820;
assign x_18705 = v_2700 | ~v_1611;
assign x_18706 = v_2700 | ~v_1741;
assign x_18707 = v_2700 | ~v_1742;
assign x_18708 = v_2700 | ~v_1614;
assign x_18709 = v_2700 | ~v_1743;
assign x_18710 = v_2700 | ~v_1744;
assign x_18711 = v_2700 | ~v_2088;
assign x_18712 = v_2700 | ~v_2089;
assign x_18713 = v_2700 | ~v_2090;
assign x_18714 = v_2700 | ~v_2091;
assign x_18715 = v_2700 | ~v_2060;
assign x_18716 = v_2700 | ~v_2136;
assign x_18717 = v_2700 | ~v_2137;
assign x_18718 = v_2700 | ~v_2063;
assign x_18719 = v_2700 | ~v_2138;
assign x_18720 = v_2700 | ~v_2139;
assign x_18721 = v_2700 | ~v_870;
assign x_18722 = v_2700 | ~v_1004;
assign x_18723 = v_2700 | ~v_1005;
assign x_18724 = v_2700 | ~v_871;
assign x_18725 = v_2700 | ~v_1006;
assign x_18726 = v_2700 | ~v_1007;
assign x_18727 = v_2700 | ~v_1008;
assign x_18728 = v_2700 | ~v_1009;
assign x_18729 = v_2700 | ~v_183;
assign x_18730 = v_2700 | ~v_180;
assign x_18731 = v_2700 | ~v_167;
assign x_18732 = v_2700 | ~v_166;
assign x_18733 = v_2700 | ~v_165;
assign x_18734 = v_2700 | ~v_144;
assign x_18735 = v_2700 | ~v_143;
assign x_18736 = v_2700 | ~v_142;
assign x_18737 = v_2700 | ~v_61;
assign x_18738 = v_2700 | ~v_60;
assign x_18739 = v_2700 | ~v_59;
assign x_18740 = v_2700 | ~v_57;
assign x_18741 = v_2699 | ~v_2671;
assign x_18742 = v_2699 | ~v_2672;
assign x_18743 = v_2699 | ~v_2673;
assign x_18744 = v_2699 | ~v_2674;
assign x_18745 = v_2699 | ~v_1808;
assign x_18746 = v_2699 | ~v_1809;
assign x_18747 = v_2699 | ~v_1810;
assign x_18748 = v_2699 | ~v_1811;
assign x_18749 = v_2699 | ~v_1586;
assign x_18750 = v_2699 | ~v_1732;
assign x_18751 = v_2699 | ~v_1733;
assign x_18752 = v_2699 | ~v_1589;
assign x_18753 = v_2699 | ~v_1734;
assign x_18754 = v_2699 | ~v_1735;
assign x_18755 = v_2699 | ~v_2083;
assign x_18756 = v_2699 | ~v_2084;
assign x_18757 = v_2699 | ~v_2085;
assign x_18758 = v_2699 | ~v_2086;
assign x_18759 = v_2699 | ~v_2045;
assign x_18760 = v_2699 | ~v_2131;
assign x_18761 = v_2699 | ~v_2132;
assign x_18762 = v_2699 | ~v_2048;
assign x_18763 = v_2699 | ~v_2133;
assign x_18764 = v_2699 | ~v_2134;
assign x_18765 = v_2699 | ~v_855;
assign x_18766 = v_2699 | ~v_989;
assign x_18767 = v_2699 | ~v_990;
assign x_18768 = v_2699 | ~v_856;
assign x_18769 = v_2699 | ~v_991;
assign x_18770 = v_2699 | ~v_992;
assign x_18771 = v_2699 | ~v_182;
assign x_18772 = v_2699 | ~v_179;
assign x_18773 = v_2699 | ~v_163;
assign x_18774 = v_2699 | ~v_162;
assign x_18775 = v_2699 | ~v_161;
assign x_18776 = v_2699 | ~v_136;
assign x_18777 = v_2699 | ~v_135;
assign x_18778 = v_2699 | ~v_134;
assign x_18779 = v_2699 | ~v_993;
assign x_18780 = v_2699 | ~v_994;
assign x_18781 = v_2699 | ~v_18;
assign x_18782 = v_2699 | ~v_17;
assign x_18783 = v_2699 | ~v_16;
assign x_18784 = v_2699 | ~v_14;
assign x_18785 = ~v_2697 | ~v_2696 | ~v_2695 | v_2698;
assign x_18786 = v_2697 | ~v_2681;
assign x_18787 = v_2697 | ~v_2682;
assign x_18788 = v_2697 | ~v_2683;
assign x_18789 = v_2697 | ~v_2684;
assign x_18790 = v_2697 | ~v_1826;
assign x_18791 = v_2697 | ~v_1827;
assign x_18792 = v_2697 | ~v_1828;
assign x_18793 = v_2697 | ~v_1829;
assign x_18794 = v_2697 | ~v_1694;
assign x_18795 = v_2697 | ~v_1695;
assign x_18796 = v_2697 | ~v_1696;
assign x_18797 = v_2697 | ~v_1697;
assign x_18798 = v_2697 | ~v_1636;
assign x_18799 = v_2697 | ~v_1639;
assign x_18800 = v_2697 | ~v_2093;
assign x_18801 = v_2697 | ~v_2094;
assign x_18802 = v_2697 | ~v_2095;
assign x_18803 = v_2697 | ~v_2096;
assign x_18804 = v_2697 | ~v_2125;
assign x_18805 = v_2697 | ~v_2126;
assign x_18806 = v_2697 | ~v_2127;
assign x_18807 = v_2697 | ~v_2128;
assign x_18808 = v_2697 | ~v_2075;
assign x_18809 = v_2697 | ~v_2078;
assign x_18810 = v_2697 | ~v_925;
assign x_18811 = v_2697 | ~v_926;
assign x_18812 = v_2697 | ~v_885;
assign x_18813 = v_2697 | ~v_886;
assign x_18814 = v_2697 | ~v_927;
assign x_18815 = v_2697 | ~v_928;
assign x_18816 = v_2697 | ~v_929;
assign x_18817 = v_2697 | ~v_930;
assign x_18818 = v_2697 | ~v_184;
assign x_18819 = v_2697 | ~v_181;
assign x_18820 = v_2697 | ~v_171;
assign x_18821 = v_2697 | ~v_170;
assign x_18822 = v_2697 | ~v_169;
assign x_18823 = v_2697 | ~v_150;
assign x_18824 = v_2697 | ~v_149;
assign x_18825 = v_2697 | ~v_147;
assign x_18826 = v_2697 | ~v_103;
assign x_18827 = v_2697 | ~v_102;
assign x_18828 = v_2697 | ~v_101;
assign x_18829 = v_2697 | ~v_96;
assign x_18830 = v_2696 | ~v_2676;
assign x_18831 = v_2696 | ~v_2677;
assign x_18832 = v_2696 | ~v_2678;
assign x_18833 = v_2696 | ~v_2679;
assign x_18834 = v_2696 | ~v_1817;
assign x_18835 = v_2696 | ~v_1818;
assign x_18836 = v_2696 | ~v_1819;
assign x_18837 = v_2696 | ~v_1820;
assign x_18838 = v_2696 | ~v_1685;
assign x_18839 = v_2696 | ~v_1686;
assign x_18840 = v_2696 | ~v_1687;
assign x_18841 = v_2696 | ~v_1688;
assign x_18842 = v_2696 | ~v_1611;
assign x_18843 = v_2696 | ~v_1614;
assign x_18844 = v_2696 | ~v_2088;
assign x_18845 = v_2696 | ~v_2089;
assign x_18846 = v_2696 | ~v_2090;
assign x_18847 = v_2696 | ~v_2091;
assign x_18848 = v_2696 | ~v_2120;
assign x_18849 = v_2696 | ~v_2121;
assign x_18850 = v_2696 | ~v_2122;
assign x_18851 = v_2696 | ~v_2123;
assign x_18852 = v_2696 | ~v_2060;
assign x_18853 = v_2696 | ~v_2063;
assign x_18854 = v_2696 | ~v_910;
assign x_18855 = v_2696 | ~v_911;
assign x_18856 = v_2696 | ~v_870;
assign x_18857 = v_2696 | ~v_871;
assign x_18858 = v_2696 | ~v_912;
assign x_18859 = v_2696 | ~v_913;
assign x_18860 = v_2696 | ~v_914;
assign x_18861 = v_2696 | ~v_915;
assign x_18862 = v_2696 | ~v_183;
assign x_18863 = v_2696 | ~v_180;
assign x_18864 = v_2696 | ~v_167;
assign x_18865 = v_2696 | ~v_166;
assign x_18866 = v_2696 | ~v_165;
assign x_18867 = v_2696 | ~v_145;
assign x_18868 = v_2696 | ~v_144;
assign x_18869 = v_2696 | ~v_142;
assign x_18870 = v_2696 | ~v_61;
assign x_18871 = v_2696 | ~v_60;
assign x_18872 = v_2696 | ~v_59;
assign x_18873 = v_2696 | ~v_54;
assign x_18874 = v_2695 | ~v_2671;
assign x_18875 = v_2695 | ~v_2672;
assign x_18876 = v_2695 | ~v_2673;
assign x_18877 = v_2695 | ~v_2674;
assign x_18878 = v_2695 | ~v_1808;
assign x_18879 = v_2695 | ~v_1809;
assign x_18880 = v_2695 | ~v_1810;
assign x_18881 = v_2695 | ~v_1811;
assign x_18882 = v_2695 | ~v_1676;
assign x_18883 = v_2695 | ~v_1677;
assign x_18884 = v_2695 | ~v_1678;
assign x_18885 = v_2695 | ~v_1679;
assign x_18886 = v_2695 | ~v_1586;
assign x_18887 = v_2695 | ~v_1589;
assign x_18888 = v_2695 | ~v_2083;
assign x_18889 = v_2695 | ~v_2084;
assign x_18890 = v_2695 | ~v_2085;
assign x_18891 = v_2695 | ~v_2086;
assign x_18892 = v_2695 | ~v_2115;
assign x_18893 = v_2695 | ~v_2116;
assign x_18894 = v_2695 | ~v_2117;
assign x_18895 = v_2695 | ~v_2118;
assign x_18896 = v_2695 | ~v_2045;
assign x_18897 = v_2695 | ~v_2048;
assign x_18898 = v_2695 | ~v_895;
assign x_18899 = v_2695 | ~v_896;
assign x_18900 = v_2695 | ~v_855;
assign x_18901 = v_2695 | ~v_856;
assign x_18902 = v_2695 | ~v_897;
assign x_18903 = v_2695 | ~v_898;
assign x_18904 = v_2695 | ~v_899;
assign x_18905 = v_2695 | ~v_900;
assign x_18906 = v_2695 | ~v_182;
assign x_18907 = v_2695 | ~v_179;
assign x_18908 = v_2695 | ~v_163;
assign x_18909 = v_2695 | ~v_162;
assign x_18910 = v_2695 | ~v_161;
assign x_18911 = v_2695 | ~v_137;
assign x_18912 = v_2695 | ~v_136;
assign x_18913 = v_2695 | ~v_134;
assign x_18914 = v_2695 | ~v_18;
assign x_18915 = v_2695 | ~v_17;
assign x_18916 = v_2695 | ~v_16;
assign x_18917 = v_2695 | ~v_11;
assign x_18918 = ~v_2693 | ~v_2692 | ~v_2691 | v_2694;
assign x_18919 = v_2693 | ~v_2681;
assign x_18920 = v_2693 | ~v_2682;
assign x_18921 = v_2693 | ~v_2683;
assign x_18922 = v_2693 | ~v_2684;
assign x_18923 = v_2693 | ~v_1826;
assign x_18924 = v_2693 | ~v_1827;
assign x_18925 = v_2693 | ~v_1828;
assign x_18926 = v_2693 | ~v_1829;
assign x_18927 = v_2693 | ~v_1632;
assign x_18928 = v_2693 | ~v_1633;
assign x_18929 = v_2693 | ~v_1634;
assign x_18930 = v_2693 | ~v_1635;
assign x_18931 = v_2693 | ~v_1636;
assign x_18932 = v_2693 | ~v_1639;
assign x_18933 = v_2693 | ~v_2093;
assign x_18934 = v_2693 | ~v_2094;
assign x_18935 = v_2693 | ~v_2095;
assign x_18936 = v_2693 | ~v_2096;
assign x_18937 = v_2693 | ~v_2109;
assign x_18938 = v_2693 | ~v_2110;
assign x_18939 = v_2693 | ~v_2111;
assign x_18940 = v_2693 | ~v_2112;
assign x_18941 = v_2693 | ~v_2075;
assign x_18942 = v_2693 | ~v_2078;
assign x_18943 = v_2693 | ~v_973;
assign x_18944 = v_2693 | ~v_974;
assign x_18945 = v_2693 | ~v_885;
assign x_18946 = v_2693 | ~v_886;
assign x_18947 = v_2693 | ~v_975;
assign x_18948 = v_2693 | ~v_976;
assign x_18949 = v_2693 | ~v_977;
assign x_18950 = v_2693 | ~v_978;
assign x_18951 = v_2693 | ~v_184;
assign x_18952 = v_2693 | ~v_181;
assign x_18953 = v_2693 | ~v_172;
assign x_18954 = v_2693 | ~v_171;
assign x_18955 = v_2693 | ~v_170;
assign x_18956 = v_2693 | ~v_169;
assign x_18957 = v_2693 | ~v_150;
assign x_18958 = v_2693 | ~v_148;
assign x_18959 = v_2693 | ~v_147;
assign x_18960 = v_2693 | ~v_102;
assign x_18961 = v_2693 | ~v_101;
assign x_18962 = v_2693 | ~v_97;
assign x_18963 = v_2692 | ~v_2676;
assign x_18964 = v_2692 | ~v_2677;
assign x_18965 = v_2692 | ~v_2678;
assign x_18966 = v_2692 | ~v_2679;
assign x_18967 = v_2692 | ~v_1817;
assign x_18968 = v_2692 | ~v_1818;
assign x_18969 = v_2692 | ~v_1819;
assign x_18970 = v_2692 | ~v_1820;
assign x_18971 = v_2692 | ~v_1607;
assign x_18972 = v_2692 | ~v_1608;
assign x_18973 = v_2692 | ~v_1609;
assign x_18974 = v_2692 | ~v_1610;
assign x_18975 = v_2692 | ~v_1611;
assign x_18976 = v_2692 | ~v_1614;
assign x_18977 = v_2692 | ~v_2088;
assign x_18978 = v_2692 | ~v_2089;
assign x_18979 = v_2692 | ~v_2090;
assign x_18980 = v_2692 | ~v_2091;
assign x_18981 = v_2692 | ~v_2104;
assign x_18982 = v_2692 | ~v_2105;
assign x_18983 = v_2692 | ~v_2106;
assign x_18984 = v_2692 | ~v_2107;
assign x_18985 = v_2692 | ~v_2060;
assign x_18986 = v_2692 | ~v_2063;
assign x_18987 = v_2692 | ~v_958;
assign x_18988 = v_2692 | ~v_959;
assign x_18989 = v_2692 | ~v_870;
assign x_18990 = v_2692 | ~v_871;
assign x_18991 = v_2692 | ~v_960;
assign x_18992 = v_2692 | ~v_961;
assign x_18993 = v_2692 | ~v_962;
assign x_18994 = v_2692 | ~v_963;
assign x_18995 = v_2692 | ~v_183;
assign x_18996 = v_2692 | ~v_180;
assign x_18997 = v_2692 | ~v_168;
assign x_18998 = v_2692 | ~v_167;
assign x_18999 = v_2692 | ~v_166;
assign x_19000 = v_2692 | ~v_165;
assign x_19001 = v_2692 | ~v_145;
assign x_19002 = v_2692 | ~v_143;
assign x_19003 = v_2692 | ~v_142;
assign x_19004 = v_2692 | ~v_60;
assign x_19005 = v_2692 | ~v_59;
assign x_19006 = v_2692 | ~v_55;
assign x_19007 = v_2691 | ~v_2671;
assign x_19008 = v_2691 | ~v_2672;
assign x_19009 = v_2691 | ~v_2673;
assign x_19010 = v_2691 | ~v_2674;
assign x_19011 = v_2691 | ~v_1808;
assign x_19012 = v_2691 | ~v_1809;
assign x_19013 = v_2691 | ~v_1810;
assign x_19014 = v_2691 | ~v_1811;
assign x_19015 = v_2691 | ~v_1582;
assign x_19016 = v_2691 | ~v_1583;
assign x_19017 = v_2691 | ~v_1584;
assign x_19018 = v_2691 | ~v_1585;
assign x_19019 = v_2691 | ~v_1586;
assign x_19020 = v_2691 | ~v_1589;
assign x_19021 = v_2691 | ~v_2083;
assign x_19022 = v_2691 | ~v_2084;
assign x_19023 = v_2691 | ~v_2085;
assign x_19024 = v_2691 | ~v_2086;
assign x_19025 = v_2691 | ~v_2099;
assign x_19026 = v_2691 | ~v_2100;
assign x_19027 = v_2691 | ~v_2101;
assign x_19028 = v_2691 | ~v_2102;
assign x_19029 = v_2691 | ~v_2045;
assign x_19030 = v_2691 | ~v_2048;
assign x_19031 = v_2691 | ~v_943;
assign x_19032 = v_2691 | ~v_944;
assign x_19033 = v_2691 | ~v_855;
assign x_19034 = v_2691 | ~v_856;
assign x_19035 = v_2691 | ~v_945;
assign x_19036 = v_2691 | ~v_946;
assign x_19037 = v_2691 | ~v_947;
assign x_19038 = v_2691 | ~v_948;
assign x_19039 = v_2691 | ~v_182;
assign x_19040 = v_2691 | ~v_179;
assign x_19041 = v_2691 | ~v_164;
assign x_19042 = v_2691 | ~v_163;
assign x_19043 = v_2691 | ~v_162;
assign x_19044 = v_2691 | ~v_161;
assign x_19045 = v_2691 | ~v_137;
assign x_19046 = v_2691 | ~v_135;
assign x_19047 = v_2691 | ~v_134;
assign x_19048 = v_2691 | ~v_17;
assign x_19049 = v_2691 | ~v_16;
assign x_19050 = v_2691 | ~v_12;
assign x_19051 = ~v_2689 | ~v_2688 | ~v_2687 | v_2690;
assign x_19052 = v_2689 | ~v_2681;
assign x_19053 = v_2689 | ~v_2682;
assign x_19054 = v_2689 | ~v_2683;
assign x_19055 = v_2689 | ~v_2684;
assign x_19056 = v_2689 | ~v_1826;
assign x_19057 = v_2689 | ~v_1827;
assign x_19058 = v_2689 | ~v_1828;
assign x_19059 = v_2689 | ~v_1829;
assign x_19060 = v_2689 | ~v_1722;
assign x_19061 = v_2689 | ~v_1723;
assign x_19062 = v_2689 | ~v_1724;
assign x_19063 = v_2689 | ~v_1725;
assign x_19064 = v_2689 | ~v_1636;
assign x_19065 = v_2689 | ~v_1639;
assign x_19066 = v_2689 | ~v_2093;
assign x_19067 = v_2689 | ~v_2094;
assign x_19068 = v_2689 | ~v_2095;
assign x_19069 = v_2689 | ~v_2096;
assign x_19070 = v_2689 | ~v_2071;
assign x_19071 = v_2689 | ~v_2072;
assign x_19072 = v_2689 | ~v_2073;
assign x_19073 = v_2689 | ~v_2074;
assign x_19074 = v_2689 | ~v_2075;
assign x_19075 = v_2689 | ~v_2078;
assign x_19076 = v_2689 | ~v_881;
assign x_19077 = v_2689 | ~v_882;
assign x_19078 = v_2689 | ~v_883;
assign x_19079 = v_2689 | ~v_884;
assign x_19080 = v_2689 | ~v_885;
assign x_19081 = v_2689 | ~v_886;
assign x_19082 = v_2689 | ~v_837;
assign x_19083 = v_2689 | ~v_838;
assign x_19084 = v_2689 | ~v_184;
assign x_19085 = v_2689 | ~v_181;
assign x_19086 = v_2689 | ~v_171;
assign x_19087 = v_2689 | ~v_170;
assign x_19088 = v_2689 | ~v_169;
assign x_19089 = v_2689 | ~v_160;
assign x_19090 = v_2689 | ~v_150;
assign x_19091 = v_2689 | ~v_149;
assign x_19092 = v_2689 | ~v_148;
assign x_19093 = v_2689 | ~v_103;
assign x_19094 = v_2689 | ~v_102;
assign x_19095 = v_2689 | ~v_95;
assign x_19096 = v_2688 | ~v_2676;
assign x_19097 = v_2688 | ~v_2677;
assign x_19098 = v_2688 | ~v_2678;
assign x_19099 = v_2688 | ~v_2679;
assign x_19100 = v_2688 | ~v_1817;
assign x_19101 = v_2688 | ~v_1818;
assign x_19102 = v_2688 | ~v_1819;
assign x_19103 = v_2688 | ~v_1820;
assign x_19104 = v_2688 | ~v_1713;
assign x_19105 = v_2688 | ~v_1714;
assign x_19106 = v_2688 | ~v_1715;
assign x_19107 = v_2688 | ~v_1716;
assign x_19108 = v_2688 | ~v_1611;
assign x_19109 = v_2688 | ~v_1614;
assign x_19110 = v_2688 | ~v_2088;
assign x_19111 = v_2688 | ~v_2089;
assign x_19112 = v_2688 | ~v_2090;
assign x_19113 = v_2688 | ~v_2091;
assign x_19114 = v_2688 | ~v_2056;
assign x_19115 = v_2688 | ~v_2057;
assign x_19116 = v_2688 | ~v_2058;
assign x_19117 = v_2688 | ~v_2059;
assign x_19118 = v_2688 | ~v_2060;
assign x_19119 = v_2688 | ~v_2063;
assign x_19120 = v_2688 | ~v_866;
assign x_19121 = v_2688 | ~v_867;
assign x_19122 = v_2688 | ~v_868;
assign x_19123 = v_2688 | ~v_869;
assign x_19124 = v_2688 | ~v_870;
assign x_19125 = v_2688 | ~v_871;
assign x_19126 = v_2688 | ~v_804;
assign x_19127 = v_2688 | ~v_805;
assign x_19128 = v_2688 | ~v_183;
assign x_19129 = v_2688 | ~v_180;
assign x_19130 = v_2688 | ~v_167;
assign x_19131 = v_2688 | ~v_166;
assign x_19132 = v_2688 | ~v_165;
assign x_19133 = v_2688 | ~v_159;
assign x_19134 = v_2688 | ~v_145;
assign x_19135 = v_2688 | ~v_144;
assign x_19136 = v_2688 | ~v_143;
assign x_19137 = v_2688 | ~v_61;
assign x_19138 = v_2688 | ~v_60;
assign x_19139 = v_2688 | ~v_53;
assign x_19140 = v_2687 | ~v_2671;
assign x_19141 = v_2687 | ~v_2672;
assign x_19142 = v_2687 | ~v_2673;
assign x_19143 = v_2687 | ~v_2674;
assign x_19144 = v_2687 | ~v_1808;
assign x_19145 = v_2687 | ~v_1809;
assign x_19146 = v_2687 | ~v_1810;
assign x_19147 = v_2687 | ~v_1811;
assign x_19148 = v_2687 | ~v_1704;
assign x_19149 = v_2687 | ~v_1705;
assign x_19150 = v_2687 | ~v_1706;
assign x_19151 = v_2687 | ~v_1707;
assign x_19152 = v_2687 | ~v_1586;
assign x_19153 = v_2687 | ~v_1589;
assign x_19154 = v_2687 | ~v_2083;
assign x_19155 = v_2687 | ~v_2084;
assign x_19156 = v_2687 | ~v_2085;
assign x_19157 = v_2687 | ~v_2086;
assign x_19158 = v_2687 | ~v_2041;
assign x_19159 = v_2687 | ~v_2042;
assign x_19160 = v_2687 | ~v_2043;
assign x_19161 = v_2687 | ~v_2044;
assign x_19162 = v_2687 | ~v_2045;
assign x_19163 = v_2687 | ~v_2048;
assign x_19164 = v_2687 | ~v_851;
assign x_19165 = v_2687 | ~v_852;
assign x_19166 = v_2687 | ~v_853;
assign x_19167 = v_2687 | ~v_854;
assign x_19168 = v_2687 | ~v_855;
assign x_19169 = v_2687 | ~v_856;
assign x_19170 = v_2687 | ~v_771;
assign x_19171 = v_2687 | ~v_772;
assign x_19172 = v_2687 | ~v_182;
assign x_19173 = v_2687 | ~v_179;
assign x_19174 = v_2687 | ~v_163;
assign x_19175 = v_2687 | ~v_162;
assign x_19176 = v_2687 | ~v_161;
assign x_19177 = v_2687 | ~v_155;
assign x_19178 = v_2687 | ~v_137;
assign x_19179 = v_2687 | ~v_136;
assign x_19180 = v_2687 | ~v_135;
assign x_19181 = v_2687 | ~v_18;
assign x_19182 = v_2687 | ~v_17;
assign x_19183 = v_2687 | ~v_10;
assign x_19184 = ~v_2685 | ~v_2680 | ~v_2675 | v_2686;
assign x_19185 = v_2685 | ~v_2681;
assign x_19186 = v_2685 | ~v_2682;
assign x_19187 = v_2685 | ~v_2683;
assign x_19188 = v_2685 | ~v_2684;
assign x_19189 = v_2685 | ~v_1722;
assign x_19190 = v_2685 | ~v_1723;
assign x_19191 = v_2685 | ~v_1724;
assign x_19192 = v_2685 | ~v_1725;
assign x_19193 = v_2685 | ~v_1636;
assign x_19194 = v_2685 | ~v_1637;
assign x_19195 = v_2685 | ~v_1638;
assign x_19196 = v_2685 | ~v_1639;
assign x_19197 = v_2685 | ~v_1640;
assign x_19198 = v_2685 | ~v_1641;
assign x_19199 = v_2685 | ~v_2071;
assign x_19200 = v_2685 | ~v_2072;
assign x_19201 = v_2685 | ~v_2073;
assign x_19202 = v_2685 | ~v_2074;
assign x_19203 = v_2685 | ~v_2075;
assign x_19204 = v_2685 | ~v_2076;
assign x_19205 = v_2685 | ~v_2077;
assign x_19206 = v_2685 | ~v_2078;
assign x_19207 = v_2685 | ~v_2079;
assign x_19208 = v_2685 | ~v_2080;
assign x_19209 = v_2685 | ~v_833;
assign x_19210 = v_2685 | ~v_834;
assign x_19211 = v_2685 | ~v_835;
assign x_19212 = v_2685 | ~v_836;
assign x_19213 = v_2685 | ~v_837;
assign x_19214 = v_2685 | ~v_838;
assign x_19215 = v_2685 | ~v_839;
assign x_19216 = v_2685 | ~v_840;
assign x_19217 = v_2685 | ~v_184;
assign x_19218 = v_2685 | ~v_170;
assign x_19219 = v_2685 | ~v_169;
assign x_19220 = v_2685 | ~v_160;
assign x_19221 = v_2685 | ~v_150;
assign x_19222 = v_2685 | ~v_149;
assign x_19223 = v_2685 | ~v_148;
assign x_19224 = v_2685 | ~v_147;
assign x_19225 = v_2685 | ~v_103;
assign x_19226 = v_2685 | ~v_102;
assign x_19227 = v_2685 | ~v_100;
assign x_19228 = v_2685 | ~v_98;
assign x_19229 = ~v_123 | ~v_174 | v_2684;
assign x_19230 = ~v_120 | ~v_173 | v_2683;
assign x_19231 = ~v_108 | v_174 | v_2682;
assign x_19232 = ~v_105 | v_173 | v_2681;
assign x_19233 = v_2680 | ~v_2676;
assign x_19234 = v_2680 | ~v_2677;
assign x_19235 = v_2680 | ~v_2678;
assign x_19236 = v_2680 | ~v_2679;
assign x_19237 = v_2680 | ~v_1713;
assign x_19238 = v_2680 | ~v_1714;
assign x_19239 = v_2680 | ~v_1715;
assign x_19240 = v_2680 | ~v_1716;
assign x_19241 = v_2680 | ~v_1611;
assign x_19242 = v_2680 | ~v_1612;
assign x_19243 = v_2680 | ~v_1613;
assign x_19244 = v_2680 | ~v_1614;
assign x_19245 = v_2680 | ~v_1615;
assign x_19246 = v_2680 | ~v_1616;
assign x_19247 = v_2680 | ~v_2056;
assign x_19248 = v_2680 | ~v_2057;
assign x_19249 = v_2680 | ~v_2058;
assign x_19250 = v_2680 | ~v_2059;
assign x_19251 = v_2680 | ~v_2060;
assign x_19252 = v_2680 | ~v_2061;
assign x_19253 = v_2680 | ~v_2062;
assign x_19254 = v_2680 | ~v_2063;
assign x_19255 = v_2680 | ~v_2064;
assign x_19256 = v_2680 | ~v_2065;
assign x_19257 = v_2680 | ~v_800;
assign x_19258 = v_2680 | ~v_801;
assign x_19259 = v_2680 | ~v_802;
assign x_19260 = v_2680 | ~v_803;
assign x_19261 = v_2680 | ~v_804;
assign x_19262 = v_2680 | ~v_805;
assign x_19263 = v_2680 | ~v_806;
assign x_19264 = v_2680 | ~v_807;
assign x_19265 = v_2680 | ~v_183;
assign x_19266 = v_2680 | ~v_166;
assign x_19267 = v_2680 | ~v_165;
assign x_19268 = v_2680 | ~v_159;
assign x_19269 = v_2680 | ~v_145;
assign x_19270 = v_2680 | ~v_144;
assign x_19271 = v_2680 | ~v_143;
assign x_19272 = v_2680 | ~v_142;
assign x_19273 = v_2680 | ~v_61;
assign x_19274 = v_2680 | ~v_60;
assign x_19275 = v_2680 | ~v_58;
assign x_19276 = v_2680 | ~v_56;
assign x_19277 = ~v_81 | ~v_174 | v_2679;
assign x_19278 = ~v_78 | ~v_173 | v_2678;
assign x_19279 = ~v_66 | v_174 | v_2677;
assign x_19280 = ~v_63 | v_173 | v_2676;
assign x_19281 = v_2675 | ~v_2671;
assign x_19282 = v_2675 | ~v_2672;
assign x_19283 = v_2675 | ~v_2673;
assign x_19284 = v_2675 | ~v_2674;
assign x_19285 = v_2675 | ~v_1704;
assign x_19286 = v_2675 | ~v_1705;
assign x_19287 = v_2675 | ~v_1706;
assign x_19288 = v_2675 | ~v_1707;
assign x_19289 = v_2675 | ~v_1586;
assign x_19290 = v_2675 | ~v_1587;
assign x_19291 = v_2675 | ~v_1588;
assign x_19292 = v_2675 | ~v_1589;
assign x_19293 = v_2675 | ~v_1590;
assign x_19294 = v_2675 | ~v_1591;
assign x_19295 = v_2675 | ~v_2041;
assign x_19296 = v_2675 | ~v_2042;
assign x_19297 = v_2675 | ~v_2043;
assign x_19298 = v_2675 | ~v_2044;
assign x_19299 = v_2675 | ~v_2045;
assign x_19300 = v_2675 | ~v_2046;
assign x_19301 = v_2675 | ~v_2047;
assign x_19302 = v_2675 | ~v_2048;
assign x_19303 = v_2675 | ~v_2049;
assign x_19304 = v_2675 | ~v_2050;
assign x_19305 = v_2675 | ~v_767;
assign x_19306 = v_2675 | ~v_768;
assign x_19307 = v_2675 | ~v_769;
assign x_19308 = v_2675 | ~v_770;
assign x_19309 = v_2675 | ~v_771;
assign x_19310 = v_2675 | ~v_772;
assign x_19311 = v_2675 | ~v_773;
assign x_19312 = v_2675 | ~v_774;
assign x_19313 = v_2675 | ~v_182;
assign x_19314 = v_2675 | ~v_162;
assign x_19315 = v_2675 | ~v_161;
assign x_19316 = v_2675 | ~v_155;
assign x_19317 = v_2675 | ~v_137;
assign x_19318 = v_2675 | ~v_136;
assign x_19319 = v_2675 | ~v_135;
assign x_19320 = v_2675 | ~v_134;
assign x_19321 = v_2675 | ~v_18;
assign x_19322 = v_2675 | ~v_17;
assign x_19323 = v_2675 | ~v_15;
assign x_19324 = v_2675 | ~v_13;
assign x_19325 = ~v_39 | ~v_174 | v_2674;
assign x_19326 = ~v_36 | ~v_173 | v_2673;
assign x_19327 = ~v_24 | v_174 | v_2672;
assign x_19328 = ~v_21 | v_173 | v_2671;
assign x_19329 = v_2670 | ~v_1566;
assign x_19330 = v_2670 | ~v_728;
assign x_19331 = v_2669 | ~v_2034;
assign x_19332 = v_2669 | ~v_735;
assign x_19333 = ~v_725 | ~v_724 | ~v_723 | ~v_722 | ~v_2667 | ~v_2663 | ~v_2659 | ~v_2655 | ~v_2651 | ~v_2647 | ~v_2643 | ~v_2639 | ~v_2635 | ~v_2631 | ~v_2627 | ~v_2623 | ~v_2619 | ~v_2615 | ~v_2611 | ~v_2607 | ~v_2591 | v_2668;
assign x_19334 = v_2667 | ~v_2664;
assign x_19335 = v_2667 | ~v_2665;
assign x_19336 = v_2667 | ~v_2666;
assign x_19337 = v_98 | v_103 | v_101 | v_100 | v_95 | v_99 | v_102 | ~v_719 | ~v_718 | v_170 | v_169 | v_149 | v_148 | v_184 | ~v_483 | ~v_717 | ~v_299 | ~v_482 | ~v_716 | ~v_298 | ~v_1962 | ~v_1898 | ~v_1961 | ~v_1897 | ~v_1896 | ~v_1960 | ~v_1895 | ~v_1959 | ~v_1894 | ~v_1893 | ~v_1464 | ~v_1352 | ~v_1463 | ~v_1351 | ~v_1350 | ~v_1462 | ~v_1349 | ~v_1461 | ~v_1348 | ~v_1347 | ~v_2605 | ~v_2604 | ~v_2603 | ~v_2602 | v_2666;
assign x_19338 = v_53 | v_56 | v_61 | v_60 | v_59 | v_58 | v_57 | ~v_714 | ~v_713 | v_144 | v_143 | v_166 | v_165 | v_183 | ~v_266 | ~v_468 | ~v_712 | ~v_467 | ~v_711 | ~v_265 | ~v_1957 | ~v_1883 | ~v_1956 | ~v_1882 | ~v_1881 | ~v_1955 | ~v_1880 | ~v_1954 | ~v_1879 | ~v_1878 | ~v_1455 | ~v_1327 | ~v_1454 | ~v_1326 | ~v_1325 | ~v_1453 | ~v_1324 | ~v_1452 | ~v_1323 | ~v_1322 | ~v_2600 | ~v_2599 | ~v_2598 | ~v_2597 | v_2665;
assign x_19339 = v_13 | v_18 | v_17 | v_16 | v_15 | v_14 | v_10 | ~v_453 | ~v_709 | ~v_452 | ~v_708 | v_136 | v_135 | ~v_707 | ~v_706 | v_162 | v_161 | v_182 | ~v_233 | ~v_232 | ~v_1952 | ~v_1868 | ~v_1951 | ~v_1867 | ~v_1866 | ~v_1950 | ~v_1865 | ~v_1949 | ~v_1864 | ~v_1863 | ~v_1446 | ~v_1302 | ~v_1445 | ~v_1301 | ~v_1300 | ~v_1444 | ~v_1299 | ~v_1443 | ~v_1298 | ~v_1297 | ~v_2595 | ~v_2594 | ~v_2593 | ~v_2592 | v_2664;
assign x_19340 = v_2663 | ~v_2660;
assign x_19341 = v_2663 | ~v_2661;
assign x_19342 = v_2663 | ~v_2662;
assign x_19343 = v_101 | v_100 | v_99 | v_93 | v_102 | v_172 | v_171 | v_170 | v_149 | v_148 | v_147 | v_184 | ~v_483 | ~v_482 | ~v_593 | ~v_592 | ~v_545 | ~v_591 | ~v_590 | ~v_544 | ~v_1962 | ~v_1961 | ~v_1896 | ~v_1960 | ~v_1959 | ~v_1893 | ~v_2014 | ~v_2013 | ~v_2012 | ~v_2011 | ~v_1464 | ~v_1463 | ~v_1350 | ~v_1462 | ~v_1461 | ~v_1347 | ~v_1496 | ~v_1495 | ~v_1494 | ~v_1493 | ~v_2605 | ~v_2604 | ~v_2603 | ~v_2602 | v_2662;
assign x_19344 = v_51 | v_60 | v_59 | v_58 | v_57 | v_144 | v_143 | v_142 | v_168 | v_167 | v_166 | v_183 | ~v_468 | ~v_467 | ~v_588 | ~v_587 | ~v_530 | ~v_586 | ~v_585 | ~v_529 | ~v_1957 | ~v_1956 | ~v_1881 | ~v_1955 | ~v_1954 | ~v_1878 | ~v_2009 | ~v_2008 | ~v_2007 | ~v_2006 | ~v_1455 | ~v_1454 | ~v_1325 | ~v_1453 | ~v_1452 | ~v_1322 | ~v_1487 | ~v_1486 | ~v_1485 | ~v_1484 | ~v_2600 | ~v_2599 | ~v_2598 | ~v_2597 | v_2661;
assign x_19345 = v_17 | v_16 | v_8 | v_15 | v_14 | ~v_453 | ~v_452 | v_136 | v_135 | v_134 | v_164 | v_163 | v_162 | v_182 | ~v_583 | ~v_582 | ~v_515 | ~v_581 | ~v_580 | ~v_514 | ~v_1952 | ~v_1951 | ~v_1866 | ~v_1950 | ~v_1949 | ~v_1863 | ~v_2004 | ~v_2003 | ~v_2002 | ~v_2001 | ~v_1446 | ~v_1445 | ~v_1300 | ~v_1444 | ~v_1443 | ~v_1297 | ~v_1478 | ~v_1477 | ~v_1476 | ~v_1475 | ~v_2595 | ~v_2594 | ~v_2593 | ~v_2592 | v_2660;
assign x_19346 = v_2659 | ~v_2656;
assign x_19347 = v_2659 | ~v_2657;
assign x_19348 = v_2659 | ~v_2658;
assign x_19349 = v_103 | v_101 | v_96 | v_100 | v_95 | v_93 | v_102 | v_171 | v_170 | v_150 | v_149 | v_184 | ~v_545 | ~v_544 | ~v_561 | ~v_560 | ~v_559 | ~v_558 | ~v_387 | ~v_386 | ~v_1896 | ~v_1893 | ~v_2014 | ~v_2013 | ~v_2012 | ~v_2011 | ~v_1946 | ~v_1945 | ~v_1944 | ~v_1943 | ~v_1350 | ~v_1347 | ~v_1408 | ~v_1407 | ~v_1406 | ~v_1405 | ~v_1496 | ~v_1495 | ~v_1494 | ~v_1493 | ~v_2605 | ~v_2604 | ~v_2603 | ~v_2602 | v_2658;
assign x_19350 = v_54 | v_53 | v_61 | v_51 | v_60 | v_59 | v_58 | v_144 | v_145 | v_167 | v_166 | v_183 | ~v_530 | ~v_529 | ~v_556 | ~v_555 | ~v_554 | ~v_553 | ~v_372 | ~v_371 | ~v_1881 | ~v_1878 | ~v_2009 | ~v_2008 | ~v_2007 | ~v_2006 | ~v_1941 | ~v_1940 | ~v_1939 | ~v_1938 | ~v_1325 | ~v_1322 | ~v_1399 | ~v_1398 | ~v_1397 | ~v_1396 | ~v_1487 | ~v_1486 | ~v_1485 | ~v_1484 | ~v_2600 | ~v_2599 | ~v_2598 | ~v_2597 | v_2657;
assign x_19351 = v_18 | v_17 | v_16 | v_8 | v_15 | v_11 | v_10 | v_136 | v_137 | v_163 | v_162 | v_182 | ~v_515 | ~v_514 | ~v_551 | ~v_550 | ~v_549 | ~v_548 | ~v_357 | ~v_356 | ~v_1866 | ~v_1863 | ~v_2004 | ~v_2003 | ~v_2002 | ~v_2001 | ~v_1936 | ~v_1935 | ~v_1934 | ~v_1933 | ~v_1300 | ~v_1297 | ~v_1390 | ~v_1389 | ~v_1388 | ~v_1387 | ~v_1478 | ~v_1477 | ~v_1476 | ~v_1475 | ~v_2595 | ~v_2594 | ~v_2593 | ~v_2592 | v_2656;
assign x_19352 = v_2655 | ~v_2652;
assign x_19353 = v_2655 | ~v_2653;
assign x_19354 = v_2655 | ~v_2654;
assign x_19355 = v_103 | v_101 | v_97 | v_100 | v_93 | v_151 | v_171 | v_170 | v_150 | v_148 | v_147 | v_184 | ~v_577 | ~v_576 | ~v_545 | ~v_544 | ~v_575 | ~v_574 | ~v_435 | ~v_434 | ~v_1896 | ~v_1893 | ~v_2014 | ~v_2013 | ~v_2012 | ~v_2011 | ~v_1930 | ~v_1929 | ~v_1928 | ~v_1927 | ~v_1350 | ~v_1347 | ~v_1346 | ~v_1345 | ~v_1344 | ~v_1343 | ~v_1496 | ~v_1495 | ~v_1494 | ~v_1493 | ~v_2605 | ~v_2604 | ~v_2603 | ~v_2602 | v_2654;
assign x_19356 = v_55 | v_61 | v_51 | v_59 | v_58 | v_145 | v_143 | v_142 | v_167 | v_166 | v_146 | v_183 | ~v_572 | ~v_571 | ~v_530 | ~v_529 | ~v_570 | ~v_569 | ~v_420 | ~v_419 | ~v_1881 | ~v_1878 | ~v_2009 | ~v_2008 | ~v_2007 | ~v_2006 | ~v_1925 | ~v_1924 | ~v_1923 | ~v_1922 | ~v_1325 | ~v_1322 | ~v_1321 | ~v_1320 | ~v_1319 | ~v_1318 | ~v_1487 | ~v_1486 | ~v_1485 | ~v_1484 | ~v_2600 | ~v_2599 | ~v_2598 | ~v_2597 | v_2653;
assign x_19357 = v_18 | v_16 | v_8 | v_15 | v_12 | v_135 | v_134 | v_137 | v_138 | v_163 | v_162 | v_182 | ~v_567 | ~v_566 | ~v_515 | ~v_514 | ~v_565 | ~v_564 | ~v_405 | ~v_404 | ~v_1866 | ~v_1863 | ~v_2004 | ~v_2003 | ~v_2002 | ~v_2001 | ~v_1920 | ~v_1919 | ~v_1918 | ~v_1917 | ~v_1300 | ~v_1297 | ~v_1296 | ~v_1295 | ~v_1294 | ~v_1293 | ~v_1478 | ~v_1477 | ~v_1476 | ~v_1475 | ~v_2595 | ~v_2594 | ~v_2593 | ~v_2592 | v_2652;
assign x_19358 = v_2651 | ~v_2648;
assign x_19359 = v_2651 | ~v_2649;
assign x_19360 = v_2651 | ~v_2650;
assign x_19361 = v_103 | v_100 | v_93 | v_102 | v_171 | v_170 | v_160 | v_150 | v_149 | v_148 | v_147 | v_184 | ~v_545 | ~v_544 | ~v_543 | ~v_542 | ~v_541 | ~v_540 | ~v_297 | ~v_296 | ~v_1896 | ~v_1893 | ~v_2014 | ~v_2013 | ~v_2012 | ~v_2011 | ~v_1892 | ~v_1891 | ~v_1890 | ~v_1889 | ~v_1350 | ~v_1347 | ~v_1436 | ~v_1435 | ~v_1434 | ~v_1433 | ~v_1496 | ~v_1495 | ~v_1494 | ~v_1493 | ~v_2605 | ~v_2604 | ~v_2603 | ~v_2602 | v_2650;
assign x_19362 = v_61 | v_51 | v_60 | v_58 | v_144 | v_159 | v_145 | v_143 | v_142 | v_167 | v_166 | v_183 | ~v_530 | ~v_529 | ~v_528 | ~v_527 | ~v_526 | ~v_525 | ~v_264 | ~v_263 | ~v_1881 | ~v_1878 | ~v_2009 | ~v_2008 | ~v_2007 | ~v_2006 | ~v_1877 | ~v_1876 | ~v_1875 | ~v_1874 | ~v_1325 | ~v_1322 | ~v_1427 | ~v_1426 | ~v_1425 | ~v_1424 | ~v_1487 | ~v_1486 | ~v_1485 | ~v_1484 | ~v_2600 | ~v_2599 | ~v_2598 | ~v_2597 | v_2649;
assign x_19363 = v_18 | v_17 | v_8 | v_15 | v_136 | v_135 | v_134 | v_137 | v_163 | v_162 | v_155 | v_182 | ~v_515 | ~v_514 | ~v_513 | ~v_512 | ~v_511 | ~v_510 | ~v_231 | ~v_230 | ~v_1866 | ~v_1863 | ~v_2004 | ~v_2003 | ~v_2002 | ~v_2001 | ~v_1862 | ~v_1861 | ~v_1860 | ~v_1859 | ~v_1300 | ~v_1297 | ~v_1418 | ~v_1417 | ~v_1416 | ~v_1415 | ~v_1478 | ~v_1477 | ~v_1476 | ~v_1475 | ~v_2595 | ~v_2594 | ~v_2593 | ~v_2592 | v_2648;
assign x_19364 = v_2647 | ~v_2644;
assign x_19365 = v_2647 | ~v_2645;
assign x_19366 = v_2647 | ~v_2646;
assign x_19367 = v_98 | v_103 | v_101 | v_96 | v_100 | v_151 | v_170 | v_169 | v_150 | v_149 | v_147 | v_184 | ~v_299 | ~v_298 | ~v_387 | ~v_386 | ~v_499 | ~v_498 | ~v_497 | ~v_496 | ~v_1898 | ~v_1897 | ~v_1896 | ~v_1895 | ~v_1894 | ~v_1893 | ~v_1946 | ~v_1945 | ~v_1944 | ~v_1943 | ~v_1352 | ~v_1351 | ~v_1350 | ~v_1349 | ~v_1348 | ~v_1347 | ~v_1408 | ~v_1407 | ~v_1406 | ~v_1405 | ~v_2605 | ~v_2604 | ~v_2603 | ~v_2602 | v_2646;
assign x_19368 = v_54 | v_56 | v_61 | v_59 | v_58 | v_144 | v_145 | v_142 | v_166 | v_165 | v_146 | v_183 | ~v_266 | ~v_265 | ~v_372 | ~v_371 | ~v_494 | ~v_493 | ~v_492 | ~v_491 | ~v_1883 | ~v_1882 | ~v_1881 | ~v_1880 | ~v_1879 | ~v_1878 | ~v_1941 | ~v_1940 | ~v_1939 | ~v_1938 | ~v_1327 | ~v_1326 | ~v_1325 | ~v_1324 | ~v_1323 | ~v_1322 | ~v_1399 | ~v_1398 | ~v_1397 | ~v_1396 | ~v_2600 | ~v_2599 | ~v_2598 | ~v_2597 | v_2645;
assign x_19369 = v_13 | v_18 | v_16 | v_15 | v_11 | v_136 | v_134 | v_137 | v_138 | v_162 | v_161 | v_182 | ~v_233 | ~v_232 | ~v_357 | ~v_356 | ~v_489 | ~v_488 | ~v_487 | ~v_486 | ~v_1868 | ~v_1867 | ~v_1866 | ~v_1865 | ~v_1864 | ~v_1863 | ~v_1936 | ~v_1935 | ~v_1934 | ~v_1933 | ~v_1302 | ~v_1301 | ~v_1300 | ~v_1299 | ~v_1298 | ~v_1297 | ~v_1390 | ~v_1389 | ~v_1388 | ~v_1387 | ~v_2595 | ~v_2594 | ~v_2593 | ~v_2592 | v_2644;
assign x_19370 = v_2643 | ~v_2640;
assign x_19371 = v_2643 | ~v_2641;
assign x_19372 = v_2643 | ~v_2642;
assign x_19373 = v_103 | v_101 | v_100 | v_94 | v_99 | v_102 | v_171 | v_169 | v_149 | v_148 | v_147 | v_184 | ~v_703 | ~v_702 | ~v_483 | ~v_482 | ~v_701 | ~v_653 | ~v_700 | ~v_652 | ~v_1962 | ~v_1961 | ~v_1896 | ~v_1960 | ~v_1959 | ~v_1893 | ~v_1982 | ~v_1981 | ~v_1980 | ~v_1979 | ~v_1464 | ~v_1463 | ~v_1350 | ~v_1462 | ~v_1461 | ~v_1347 | ~v_1380 | ~v_1379 | ~v_1378 | ~v_1377 | ~v_2605 | ~v_2604 | ~v_2603 | ~v_2602 | v_2642;
assign x_19374 = v_61 | v_52 | v_60 | v_59 | v_58 | v_57 | v_144 | v_143 | v_142 | v_167 | v_165 | v_183 | ~v_698 | ~v_697 | ~v_468 | ~v_467 | ~v_696 | ~v_638 | ~v_695 | ~v_637 | ~v_1957 | ~v_1956 | ~v_1881 | ~v_1955 | ~v_1954 | ~v_1878 | ~v_1977 | ~v_1976 | ~v_1975 | ~v_1974 | ~v_1455 | ~v_1454 | ~v_1325 | ~v_1453 | ~v_1452 | ~v_1322 | ~v_1371 | ~v_1370 | ~v_1369 | ~v_1368 | ~v_2600 | ~v_2599 | ~v_2598 | ~v_2597 | v_2641;
assign x_19375 = v_9 | v_18 | v_17 | v_16 | v_15 | v_14 | ~v_453 | ~v_452 | v_136 | v_135 | v_134 | v_163 | v_161 | v_182 | ~v_693 | ~v_692 | ~v_691 | ~v_623 | ~v_690 | ~v_622 | ~v_1952 | ~v_1951 | ~v_1866 | ~v_1950 | ~v_1949 | ~v_1863 | ~v_1972 | ~v_1971 | ~v_1970 | ~v_1969 | ~v_1446 | ~v_1445 | ~v_1300 | ~v_1444 | ~v_1443 | ~v_1297 | ~v_1362 | ~v_1361 | ~v_1360 | ~v_1359 | ~v_2595 | ~v_2594 | ~v_2593 | ~v_2592 | v_2640;
assign x_19376 = v_2639 | ~v_2636;
assign x_19377 = v_2639 | ~v_2637;
assign x_19378 = v_2639 | ~v_2638;
assign x_19379 = v_101 | v_96 | v_100 | v_94 | v_102 | v_172 | v_171 | v_169 | v_150 | v_149 | v_147 | v_184 | ~v_671 | ~v_670 | ~v_387 | ~v_386 | ~v_653 | ~v_652 | ~v_669 | ~v_668 | ~v_1896 | ~v_1893 | ~v_1946 | ~v_1945 | ~v_1944 | ~v_1943 | ~v_1982 | ~v_1981 | ~v_1980 | ~v_1979 | ~v_1350 | ~v_1347 | ~v_1380 | ~v_1379 | ~v_1378 | ~v_1377 | ~v_1408 | ~v_1407 | ~v_1406 | ~v_1405 | ~v_2605 | ~v_2604 | ~v_2603 | ~v_2602 | v_2638;
assign x_19380 = v_54 | v_52 | v_60 | v_59 | v_58 | v_144 | v_145 | v_142 | v_168 | v_167 | v_165 | v_183 | ~v_666 | ~v_665 | ~v_372 | ~v_371 | ~v_638 | ~v_637 | ~v_664 | ~v_663 | ~v_1881 | ~v_1878 | ~v_1941 | ~v_1940 | ~v_1939 | ~v_1938 | ~v_1977 | ~v_1976 | ~v_1975 | ~v_1974 | ~v_1325 | ~v_1322 | ~v_1371 | ~v_1370 | ~v_1369 | ~v_1368 | ~v_1399 | ~v_1398 | ~v_1397 | ~v_1396 | ~v_2600 | ~v_2599 | ~v_2598 | ~v_2597 | v_2637;
assign x_19381 = v_9 | v_17 | v_16 | v_15 | v_11 | v_136 | v_134 | v_137 | v_164 | v_163 | v_161 | v_182 | ~v_661 | ~v_660 | ~v_357 | ~v_356 | ~v_623 | ~v_622 | ~v_659 | ~v_658 | ~v_1866 | ~v_1863 | ~v_1936 | ~v_1935 | ~v_1934 | ~v_1933 | ~v_1972 | ~v_1971 | ~v_1970 | ~v_1969 | ~v_1300 | ~v_1297 | ~v_1362 | ~v_1361 | ~v_1360 | ~v_1359 | ~v_1390 | ~v_1389 | ~v_1388 | ~v_1387 | ~v_2595 | ~v_2594 | ~v_2593 | ~v_2592 | v_2636;
assign x_19382 = v_2635 | ~v_2632;
assign x_19383 = v_2635 | ~v_2633;
assign x_19384 = v_2635 | ~v_2634;
assign x_19385 = v_103 | v_101 | v_97 | v_100 | v_95 | v_94 | v_102 | v_171 | v_169 | v_150 | v_148 | v_184 | ~v_435 | ~v_434 | ~v_653 | ~v_652 | ~v_687 | ~v_686 | ~v_685 | ~v_684 | ~v_1896 | ~v_1893 | ~v_1930 | ~v_1929 | ~v_1928 | ~v_1927 | ~v_1982 | ~v_1981 | ~v_1980 | ~v_1979 | ~v_1350 | ~v_1347 | ~v_1380 | ~v_1379 | ~v_1378 | ~v_1377 | ~v_1346 | ~v_1345 | ~v_1344 | ~v_1343 | ~v_2605 | ~v_2604 | ~v_2603 | ~v_2602 | v_2634;
assign x_19386 = v_53 | v_55 | v_61 | v_52 | v_60 | v_59 | v_58 | v_145 | v_143 | v_167 | v_165 | v_183 | ~v_420 | ~v_419 | ~v_638 | ~v_637 | ~v_682 | ~v_681 | ~v_680 | ~v_679 | ~v_1881 | ~v_1878 | ~v_1925 | ~v_1924 | ~v_1923 | ~v_1922 | ~v_1977 | ~v_1976 | ~v_1975 | ~v_1974 | ~v_1325 | ~v_1322 | ~v_1371 | ~v_1370 | ~v_1369 | ~v_1368 | ~v_1321 | ~v_1320 | ~v_1319 | ~v_1318 | ~v_2600 | ~v_2599 | ~v_2598 | ~v_2597 | v_2633;
assign x_19387 = v_9 | v_18 | v_17 | v_16 | v_15 | v_12 | v_10 | v_135 | v_137 | v_163 | v_161 | v_182 | ~v_405 | ~v_404 | ~v_623 | ~v_622 | ~v_677 | ~v_676 | ~v_675 | ~v_674 | ~v_1866 | ~v_1863 | ~v_1920 | ~v_1919 | ~v_1918 | ~v_1917 | ~v_1972 | ~v_1971 | ~v_1970 | ~v_1969 | ~v_1300 | ~v_1297 | ~v_1362 | ~v_1361 | ~v_1360 | ~v_1359 | ~v_1296 | ~v_1295 | ~v_1294 | ~v_1293 | ~v_2595 | ~v_2594 | ~v_2593 | ~v_2592 | v_2632;
assign x_19388 = v_2631 | ~v_2628;
assign x_19389 = v_2631 | ~v_2629;
assign x_19390 = v_2631 | ~v_2630;
assign x_19391 = v_103 | v_100 | v_94 | v_151 | v_171 | v_169 | v_160 | v_150 | v_149 | v_148 | v_147 | v_184 | ~v_655 | ~v_654 | ~v_297 | ~v_296 | ~v_653 | ~v_652 | ~v_651 | ~v_650 | ~v_1896 | ~v_1893 | ~v_1892 | ~v_1891 | ~v_1890 | ~v_1889 | ~v_1982 | ~v_1981 | ~v_1980 | ~v_1979 | ~v_1350 | ~v_1347 | ~v_1380 | ~v_1379 | ~v_1378 | ~v_1377 | ~v_1436 | ~v_1435 | ~v_1434 | ~v_1433 | ~v_2605 | ~v_2604 | ~v_2603 | ~v_2602 | v_2630;
assign x_19392 = v_61 | v_52 | v_58 | v_144 | v_159 | v_145 | v_143 | v_142 | v_167 | v_165 | v_146 | v_183 | ~v_640 | ~v_639 | ~v_264 | ~v_263 | ~v_638 | ~v_637 | ~v_636 | ~v_635 | ~v_1881 | ~v_1878 | ~v_1877 | ~v_1876 | ~v_1875 | ~v_1874 | ~v_1977 | ~v_1976 | ~v_1975 | ~v_1974 | ~v_1325 | ~v_1322 | ~v_1371 | ~v_1370 | ~v_1369 | ~v_1368 | ~v_1427 | ~v_1426 | ~v_1425 | ~v_1424 | ~v_2600 | ~v_2599 | ~v_2598 | ~v_2597 | v_2629;
assign x_19393 = v_9 | v_18 | v_15 | v_136 | v_135 | v_134 | v_137 | v_138 | v_163 | v_161 | v_155 | v_182 | ~v_625 | ~v_624 | ~v_231 | ~v_230 | ~v_623 | ~v_622 | ~v_621 | ~v_620 | ~v_1866 | ~v_1863 | ~v_1862 | ~v_1861 | ~v_1860 | ~v_1859 | ~v_1972 | ~v_1971 | ~v_1970 | ~v_1969 | ~v_1300 | ~v_1297 | ~v_1362 | ~v_1361 | ~v_1360 | ~v_1359 | ~v_1418 | ~v_1417 | ~v_1416 | ~v_1415 | ~v_2595 | ~v_2594 | ~v_2593 | ~v_2592 | v_2628;
assign x_19394 = v_2627 | ~v_2624;
assign x_19395 = v_2627 | ~v_2625;
assign x_19396 = v_2627 | ~v_2626;
assign x_19397 = v_98 | v_103 | v_101 | v_97 | v_100 | v_102 | v_170 | v_169 | v_150 | v_148 | v_147 | v_184 | ~v_609 | ~v_608 | ~v_299 | ~v_298 | ~v_435 | ~v_434 | ~v_607 | ~v_606 | ~v_1898 | ~v_1897 | ~v_1896 | ~v_1895 | ~v_1894 | ~v_1893 | ~v_1930 | ~v_1929 | ~v_1928 | ~v_1927 | ~v_1352 | ~v_1351 | ~v_1350 | ~v_1349 | ~v_1348 | ~v_1347 | ~v_1346 | ~v_1345 | ~v_1344 | ~v_1343 | ~v_2605 | ~v_2604 | ~v_2603 | ~v_2602 | v_2626;
assign x_19398 = v_56 | v_55 | v_61 | v_60 | v_59 | v_58 | v_145 | v_143 | v_142 | v_166 | v_165 | v_183 | ~v_604 | ~v_603 | ~v_266 | ~v_265 | ~v_420 | ~v_419 | ~v_602 | ~v_601 | ~v_1883 | ~v_1882 | ~v_1881 | ~v_1880 | ~v_1879 | ~v_1878 | ~v_1925 | ~v_1924 | ~v_1923 | ~v_1922 | ~v_1327 | ~v_1326 | ~v_1325 | ~v_1324 | ~v_1323 | ~v_1322 | ~v_1321 | ~v_1320 | ~v_1319 | ~v_1318 | ~v_2600 | ~v_2599 | ~v_2598 | ~v_2597 | v_2625;
assign x_19399 = v_13 | v_18 | v_17 | v_16 | v_15 | v_12 | v_135 | v_134 | v_137 | v_162 | v_161 | v_182 | ~v_599 | ~v_598 | ~v_233 | ~v_232 | ~v_405 | ~v_404 | ~v_597 | ~v_596 | ~v_1868 | ~v_1867 | ~v_1866 | ~v_1865 | ~v_1864 | ~v_1863 | ~v_1920 | ~v_1919 | ~v_1918 | ~v_1917 | ~v_1302 | ~v_1301 | ~v_1300 | ~v_1299 | ~v_1298 | ~v_1297 | ~v_1296 | ~v_1295 | ~v_1294 | ~v_1293 | ~v_2595 | ~v_2594 | ~v_2593 | ~v_2592 | v_2624;
assign x_19400 = v_2623 | ~v_2620;
assign x_19401 = v_2623 | ~v_2621;
assign x_19402 = v_2623 | ~v_2622;
assign x_19403 = v_103 | v_101 | v_99 | v_102 | v_171 | v_170 | v_169 | v_149 | v_148 | v_147 | v_184 | v_181 | ~v_483 | ~v_482 | ~v_481 | ~v_480 | ~v_345 | ~v_479 | ~v_478 | ~v_344 | ~v_1962 | ~v_1961 | ~v_1896 | ~v_1960 | ~v_1959 | ~v_1893 | ~v_1914 | ~v_1913 | ~v_1912 | ~v_1911 | ~v_1464 | ~v_1463 | ~v_1350 | ~v_1462 | ~v_1461 | ~v_1347 | ~v_1540 | ~v_1539 | ~v_1538 | ~v_1537 | ~v_2605 | ~v_2604 | ~v_2603 | ~v_2602 | v_2622;
assign x_19404 = v_61 | v_60 | v_59 | v_57 | v_144 | v_180 | v_143 | v_142 | v_167 | v_166 | v_165 | v_183 | ~v_468 | ~v_467 | ~v_466 | ~v_465 | ~v_330 | ~v_464 | ~v_463 | ~v_329 | ~v_1957 | ~v_1956 | ~v_1881 | ~v_1955 | ~v_1954 | ~v_1878 | ~v_1909 | ~v_1908 | ~v_1907 | ~v_1906 | ~v_1455 | ~v_1454 | ~v_1325 | ~v_1453 | ~v_1452 | ~v_1322 | ~v_1531 | ~v_1530 | ~v_1529 | ~v_1528 | ~v_2600 | ~v_2599 | ~v_2598 | ~v_2597 | v_2621;
assign x_19405 = v_18 | v_17 | v_16 | v_14 | ~v_453 | ~v_452 | v_136 | v_135 | v_134 | v_179 | v_163 | v_162 | v_161 | v_182 | ~v_451 | ~v_450 | ~v_315 | ~v_449 | ~v_448 | ~v_314 | ~v_1952 | ~v_1951 | ~v_1866 | ~v_1950 | ~v_1949 | ~v_1863 | ~v_1904 | ~v_1903 | ~v_1902 | ~v_1901 | ~v_1446 | ~v_1445 | ~v_1300 | ~v_1444 | ~v_1443 | ~v_1297 | ~v_1522 | ~v_1521 | ~v_1520 | ~v_1519 | ~v_2595 | ~v_2594 | ~v_2593 | ~v_2592 | v_2620;
assign x_19406 = v_2619 | ~v_2616;
assign x_19407 = v_2619 | ~v_2617;
assign x_19408 = v_2619 | ~v_2618;
assign x_19409 = v_103 | v_101 | v_96 | v_102 | v_171 | v_170 | v_169 | v_150 | v_149 | v_147 | v_184 | v_181 | ~v_391 | ~v_390 | ~v_387 | ~v_386 | ~v_345 | ~v_344 | ~v_385 | ~v_384 | ~v_1896 | ~v_1893 | ~v_1946 | ~v_1945 | ~v_1944 | ~v_1943 | ~v_1914 | ~v_1913 | ~v_1912 | ~v_1911 | ~v_1350 | ~v_1347 | ~v_1408 | ~v_1407 | ~v_1406 | ~v_1405 | ~v_1540 | ~v_1539 | ~v_1538 | ~v_1537 | ~v_2605 | ~v_2604 | ~v_2603 | ~v_2602 | v_2618;
assign x_19410 = v_54 | v_61 | v_60 | v_59 | v_144 | v_180 | v_145 | v_142 | v_167 | v_166 | v_165 | v_183 | ~v_376 | ~v_375 | ~v_372 | ~v_371 | ~v_330 | ~v_329 | ~v_370 | ~v_369 | ~v_1881 | ~v_1878 | ~v_1941 | ~v_1940 | ~v_1939 | ~v_1938 | ~v_1909 | ~v_1908 | ~v_1907 | ~v_1906 | ~v_1325 | ~v_1322 | ~v_1399 | ~v_1398 | ~v_1397 | ~v_1396 | ~v_1531 | ~v_1530 | ~v_1529 | ~v_1528 | ~v_2600 | ~v_2599 | ~v_2598 | ~v_2597 | v_2617;
assign x_19411 = v_18 | v_17 | v_16 | v_11 | v_136 | v_134 | v_137 | v_179 | v_163 | v_162 | v_161 | v_182 | ~v_361 | ~v_360 | ~v_357 | ~v_356 | ~v_315 | ~v_314 | ~v_355 | ~v_354 | ~v_1866 | ~v_1863 | ~v_1936 | ~v_1935 | ~v_1934 | ~v_1933 | ~v_1904 | ~v_1903 | ~v_1902 | ~v_1901 | ~v_1300 | ~v_1297 | ~v_1390 | ~v_1389 | ~v_1388 | ~v_1387 | ~v_1522 | ~v_1521 | ~v_1520 | ~v_1519 | ~v_2595 | ~v_2594 | ~v_2593 | ~v_2592 | v_2616;
assign x_19412 = v_2615 | ~v_2612;
assign x_19413 = v_2615 | ~v_2613;
assign x_19414 = v_2615 | ~v_2614;
assign x_19415 = v_101 | v_97 | v_102 | v_172 | v_171 | v_170 | v_169 | v_150 | v_148 | v_147 | v_184 | v_181 | ~v_437 | ~v_436 | ~v_435 | ~v_434 | ~v_345 | ~v_344 | ~v_433 | ~v_432 | ~v_1896 | ~v_1893 | ~v_1930 | ~v_1929 | ~v_1928 | ~v_1927 | ~v_1914 | ~v_1913 | ~v_1912 | ~v_1911 | ~v_1350 | ~v_1347 | ~v_1346 | ~v_1345 | ~v_1344 | ~v_1343 | ~v_1540 | ~v_1539 | ~v_1538 | ~v_1537 | ~v_2605 | ~v_2604 | ~v_2603 | ~v_2602 | v_2614;
assign x_19416 = v_55 | v_60 | v_59 | v_180 | v_145 | v_143 | v_142 | v_168 | v_167 | v_166 | v_165 | v_183 | ~v_422 | ~v_421 | ~v_420 | ~v_419 | ~v_330 | ~v_329 | ~v_418 | ~v_417 | ~v_1881 | ~v_1878 | ~v_1925 | ~v_1924 | ~v_1923 | ~v_1922 | ~v_1909 | ~v_1908 | ~v_1907 | ~v_1906 | ~v_1325 | ~v_1322 | ~v_1321 | ~v_1320 | ~v_1319 | ~v_1318 | ~v_1531 | ~v_1530 | ~v_1529 | ~v_1528 | ~v_2600 | ~v_2599 | ~v_2598 | ~v_2597 | v_2613;
assign x_19417 = v_17 | v_16 | v_12 | v_135 | v_134 | v_137 | v_179 | v_164 | v_163 | v_162 | v_161 | v_182 | ~v_407 | ~v_406 | ~v_405 | ~v_404 | ~v_315 | ~v_314 | ~v_403 | ~v_402 | ~v_1866 | ~v_1863 | ~v_1920 | ~v_1919 | ~v_1918 | ~v_1917 | ~v_1904 | ~v_1903 | ~v_1902 | ~v_1901 | ~v_1300 | ~v_1297 | ~v_1296 | ~v_1295 | ~v_1294 | ~v_1293 | ~v_1522 | ~v_1521 | ~v_1520 | ~v_1519 | ~v_2595 | ~v_2594 | ~v_2593 | ~v_2592 | v_2612;
assign x_19418 = v_2611 | ~v_2608;
assign x_19419 = v_2611 | ~v_2609;
assign x_19420 = v_2611 | ~v_2610;
assign x_19421 = v_103 | v_95 | v_102 | v_171 | v_170 | v_169 | v_160 | v_150 | v_149 | v_148 | v_184 | v_181 | ~v_297 | ~v_296 | ~v_345 | ~v_344 | ~v_343 | ~v_342 | ~v_341 | ~v_340 | ~v_1896 | ~v_1893 | ~v_1892 | ~v_1891 | ~v_1890 | ~v_1889 | ~v_1914 | ~v_1913 | ~v_1912 | ~v_1911 | ~v_1350 | ~v_1347 | ~v_1436 | ~v_1435 | ~v_1434 | ~v_1433 | ~v_1540 | ~v_1539 | ~v_1538 | ~v_1537 | ~v_2605 | ~v_2604 | ~v_2603 | ~v_2602 | v_2610;
assign x_19422 = v_53 | v_61 | v_60 | v_144 | v_180 | v_159 | v_145 | v_143 | v_167 | v_166 | v_165 | v_183 | ~v_264 | ~v_263 | ~v_330 | ~v_329 | ~v_328 | ~v_327 | ~v_326 | ~v_325 | ~v_1881 | ~v_1878 | ~v_1877 | ~v_1876 | ~v_1875 | ~v_1874 | ~v_1909 | ~v_1908 | ~v_1907 | ~v_1906 | ~v_1325 | ~v_1322 | ~v_1427 | ~v_1426 | ~v_1425 | ~v_1424 | ~v_1531 | ~v_1530 | ~v_1529 | ~v_1528 | ~v_2600 | ~v_2599 | ~v_2598 | ~v_2597 | v_2609;
assign x_19423 = v_18 | v_17 | v_10 | v_136 | v_135 | v_137 | v_179 | v_163 | v_162 | v_161 | v_155 | v_182 | ~v_231 | ~v_230 | ~v_315 | ~v_314 | ~v_313 | ~v_312 | ~v_311 | ~v_310 | ~v_1866 | ~v_1863 | ~v_1862 | ~v_1861 | ~v_1860 | ~v_1859 | ~v_1904 | ~v_1903 | ~v_1902 | ~v_1901 | ~v_1300 | ~v_1297 | ~v_1418 | ~v_1417 | ~v_1416 | ~v_1415 | ~v_1522 | ~v_1521 | ~v_1520 | ~v_1519 | ~v_2595 | ~v_2594 | ~v_2593 | ~v_2592 | v_2608;
assign x_19424 = v_2607 | ~v_2596;
assign x_19425 = v_2607 | ~v_2601;
assign x_19426 = v_2607 | ~v_2606;
assign x_19427 = v_98 | v_103 | v_100 | v_102 | v_170 | v_169 | v_160 | v_150 | v_149 | v_148 | v_147 | v_184 | ~v_299 | ~v_298 | ~v_297 | ~v_296 | ~v_295 | ~v_294 | ~v_293 | ~v_292 | ~v_1898 | ~v_1897 | ~v_1896 | ~v_1895 | ~v_1894 | ~v_1893 | ~v_1892 | ~v_1891 | ~v_1890 | ~v_1889 | ~v_1352 | ~v_1351 | ~v_1350 | ~v_1349 | ~v_1348 | ~v_1347 | ~v_1436 | ~v_1435 | ~v_1434 | ~v_1433 | ~v_2605 | ~v_2604 | ~v_2603 | ~v_2602 | v_2606;
assign x_19428 = v_2605 | v_174;
assign x_19429 = v_2605 | v_123;
assign x_19430 = v_2604 | v_173;
assign x_19431 = v_2604 | v_120;
assign x_19432 = v_2603 | ~v_174;
assign x_19433 = v_2603 | v_108;
assign x_19434 = v_2602 | ~v_173;
assign x_19435 = v_2602 | v_105;
assign x_19436 = v_56 | v_61 | v_60 | v_58 | v_144 | v_159 | v_145 | v_143 | v_142 | v_166 | v_165 | v_183 | ~v_266 | ~v_265 | ~v_264 | ~v_263 | ~v_262 | ~v_261 | ~v_260 | ~v_259 | ~v_1883 | ~v_1882 | ~v_1881 | ~v_1880 | ~v_1879 | ~v_1878 | ~v_1877 | ~v_1876 | ~v_1875 | ~v_1874 | ~v_1327 | ~v_1326 | ~v_1325 | ~v_1324 | ~v_1323 | ~v_1322 | ~v_1427 | ~v_1426 | ~v_1425 | ~v_1424 | ~v_2600 | ~v_2599 | ~v_2598 | ~v_2597 | v_2601;
assign x_19437 = v_2600 | v_174;
assign x_19438 = v_2600 | v_81;
assign x_19439 = v_2599 | v_173;
assign x_19440 = v_2599 | v_78;
assign x_19441 = v_2598 | ~v_174;
assign x_19442 = v_2598 | v_66;
assign x_19443 = v_2597 | ~v_173;
assign x_19444 = v_2597 | v_63;
assign x_19445 = v_13 | v_18 | v_17 | v_15 | v_136 | v_135 | v_134 | v_137 | v_162 | v_161 | v_155 | v_182 | ~v_233 | ~v_232 | ~v_231 | ~v_230 | ~v_229 | ~v_228 | ~v_227 | ~v_226 | ~v_1868 | ~v_1867 | ~v_1866 | ~v_1865 | ~v_1864 | ~v_1863 | ~v_1862 | ~v_1861 | ~v_1860 | ~v_1859 | ~v_1302 | ~v_1301 | ~v_1300 | ~v_1299 | ~v_1298 | ~v_1297 | ~v_1418 | ~v_1417 | ~v_1416 | ~v_1415 | ~v_2595 | ~v_2594 | ~v_2593 | ~v_2592 | v_2596;
assign x_19446 = v_2595 | v_174;
assign x_19447 = v_2595 | v_39;
assign x_19448 = v_2594 | v_173;
assign x_19449 = v_2594 | v_36;
assign x_19450 = v_2593 | ~v_174;
assign x_19451 = v_2593 | v_24;
assign x_19452 = v_2592 | ~v_173;
assign x_19453 = v_2592 | v_21;
assign x_19454 = v_2591 | ~v_2589;
assign x_19455 = v_2591 | ~v_2590;
assign x_19456 = v_2591 | ~v_1270;
assign x_19457 = v_2591 | ~v_1271;
assign x_19458 = v_2591 | ~v_174;
assign x_19459 = v_2591 | ~v_173;
assign x_19460 = ~v_186 | ~v_1276 | v_2590;
assign x_19461 = ~v_195 | ~v_1851 | v_2589;
assign x_19462 = v_2588 | ~v_2402;
assign x_19463 = v_2588 | ~v_2587;
assign x_19464 = v_176 | v_175 | ~v_2586 | ~v_732 | ~v_729 | ~v_2407 | ~v_2403 | v_2587;
assign x_19465 = v_2586 | ~v_2453;
assign x_19466 = v_2586 | ~v_2469;
assign x_19467 = v_2586 | ~v_2485;
assign x_19468 = v_2586 | ~v_2501;
assign x_19469 = v_2586 | ~v_2517;
assign x_19470 = v_2586 | ~v_2521;
assign x_19471 = v_2586 | ~v_2537;
assign x_19472 = v_2586 | ~v_2541;
assign x_19473 = v_2586 | ~v_2545;
assign x_19474 = v_2586 | ~v_2549;
assign x_19475 = v_2586 | ~v_2553;
assign x_19476 = v_2586 | ~v_2569;
assign x_19477 = v_2586 | ~v_2573;
assign x_19478 = v_2586 | ~v_2577;
assign x_19479 = v_2586 | ~v_2581;
assign x_19480 = v_2586 | ~v_2585;
assign x_19481 = v_2586 | ~v_1263;
assign x_19482 = v_2586 | ~v_1264;
assign x_19483 = v_2586 | ~v_1265;
assign x_19484 = v_2586 | ~v_1266;
assign x_19485 = ~v_2584 | ~v_2583 | ~v_2582 | v_2585;
assign x_19486 = v_2584 | ~v_2438;
assign x_19487 = v_2584 | ~v_2439;
assign x_19488 = v_2584 | ~v_2440;
assign x_19489 = v_2584 | ~v_2441;
assign x_19490 = v_2584 | ~v_1626;
assign x_19491 = v_2584 | ~v_1627;
assign x_19492 = v_2584 | ~v_1746;
assign x_19493 = v_2584 | ~v_1628;
assign x_19494 = v_2584 | ~v_1747;
assign x_19495 = v_2584 | ~v_1629;
assign x_19496 = v_2584 | ~v_1630;
assign x_19497 = v_2584 | ~v_1748;
assign x_19498 = v_2584 | ~v_1631;
assign x_19499 = v_2584 | ~v_1749;
assign x_19500 = v_2584 | ~v_839;
assign x_19501 = v_2584 | ~v_1257;
assign x_19502 = v_2584 | ~v_1023;
assign x_19503 = v_2584 | ~v_840;
assign x_19504 = v_2584 | ~v_1258;
assign x_19505 = v_2584 | ~v_1024;
assign x_19506 = v_2584 | ~v_2446;
assign x_19507 = v_2584 | ~v_2447;
assign x_19508 = v_2584 | ~v_2512;
assign x_19509 = v_2584 | ~v_2448;
assign x_19510 = v_2584 | ~v_2513;
assign x_19511 = v_2584 | ~v_2449;
assign x_19512 = v_2584 | ~v_2450;
assign x_19513 = v_2584 | ~v_2514;
assign x_19514 = v_2584 | ~v_2451;
assign x_19515 = v_2584 | ~v_2515;
assign x_19516 = v_2584 | ~v_184;
assign x_19517 = v_2584 | ~v_170;
assign x_19518 = v_2584 | ~v_169;
assign x_19519 = v_2584 | ~v_149;
assign x_19520 = v_2584 | ~v_148;
assign x_19521 = v_2584 | ~v_1259;
assign x_19522 = v_2584 | ~v_1260;
assign x_19523 = v_2584 | ~v_103;
assign x_19524 = v_2584 | ~v_102;
assign x_19525 = v_2584 | ~v_101;
assign x_19526 = v_2584 | ~v_100;
assign x_19527 = v_2584 | ~v_99;
assign x_19528 = v_2584 | ~v_98;
assign x_19529 = v_2584 | ~v_95;
assign x_19530 = v_2583 | ~v_2423;
assign x_19531 = v_2583 | ~v_2424;
assign x_19532 = v_2583 | ~v_2425;
assign x_19533 = v_2583 | ~v_2426;
assign x_19534 = v_2583 | ~v_1601;
assign x_19535 = v_2583 | ~v_1602;
assign x_19536 = v_2583 | ~v_1737;
assign x_19537 = v_2583 | ~v_1603;
assign x_19538 = v_2583 | ~v_1738;
assign x_19539 = v_2583 | ~v_1604;
assign x_19540 = v_2583 | ~v_1605;
assign x_19541 = v_2583 | ~v_1739;
assign x_19542 = v_2583 | ~v_1606;
assign x_19543 = v_2583 | ~v_1740;
assign x_19544 = v_2583 | ~v_806;
assign x_19545 = v_2583 | ~v_1252;
assign x_19546 = v_2583 | ~v_1008;
assign x_19547 = v_2583 | ~v_1253;
assign x_19548 = v_2583 | ~v_1009;
assign x_19549 = v_2583 | ~v_2431;
assign x_19550 = v_2583 | ~v_2432;
assign x_19551 = v_2583 | ~v_2507;
assign x_19552 = v_2583 | ~v_2433;
assign x_19553 = v_2583 | ~v_2508;
assign x_19554 = v_2583 | ~v_2434;
assign x_19555 = v_2583 | ~v_2435;
assign x_19556 = v_2583 | ~v_2509;
assign x_19557 = v_2583 | ~v_2436;
assign x_19558 = v_2583 | ~v_2510;
assign x_19559 = v_2583 | ~v_807;
assign x_19560 = v_2583 | ~v_183;
assign x_19561 = v_2583 | ~v_166;
assign x_19562 = v_2583 | ~v_165;
assign x_19563 = v_2583 | ~v_144;
assign x_19564 = v_2583 | ~v_143;
assign x_19565 = v_2583 | ~v_1254;
assign x_19566 = v_2583 | ~v_1255;
assign x_19567 = v_2583 | ~v_61;
assign x_19568 = v_2583 | ~v_60;
assign x_19569 = v_2583 | ~v_59;
assign x_19570 = v_2583 | ~v_58;
assign x_19571 = v_2583 | ~v_57;
assign x_19572 = v_2583 | ~v_56;
assign x_19573 = v_2583 | ~v_53;
assign x_19574 = v_2582 | ~v_2408;
assign x_19575 = v_2582 | ~v_2409;
assign x_19576 = v_2582 | ~v_2410;
assign x_19577 = v_2582 | ~v_2411;
assign x_19578 = v_2582 | ~v_1576;
assign x_19579 = v_2582 | ~v_1577;
assign x_19580 = v_2582 | ~v_1728;
assign x_19581 = v_2582 | ~v_1578;
assign x_19582 = v_2582 | ~v_1729;
assign x_19583 = v_2582 | ~v_1579;
assign x_19584 = v_2582 | ~v_1580;
assign x_19585 = v_2582 | ~v_1730;
assign x_19586 = v_2582 | ~v_1581;
assign x_19587 = v_2582 | ~v_1731;
assign x_19588 = v_2582 | ~v_773;
assign x_19589 = v_2582 | ~v_774;
assign x_19590 = v_2582 | ~v_2416;
assign x_19591 = v_2582 | ~v_2417;
assign x_19592 = v_2582 | ~v_2502;
assign x_19593 = v_2582 | ~v_2418;
assign x_19594 = v_2582 | ~v_2503;
assign x_19595 = v_2582 | ~v_2419;
assign x_19596 = v_2582 | ~v_2420;
assign x_19597 = v_2582 | ~v_2504;
assign x_19598 = v_2582 | ~v_2421;
assign x_19599 = v_2582 | ~v_2505;
assign x_19600 = v_2582 | ~v_182;
assign x_19601 = v_2582 | ~v_162;
assign x_19602 = v_2582 | ~v_161;
assign x_19603 = v_2582 | ~v_1247;
assign x_19604 = v_2582 | ~v_1248;
assign x_19605 = v_2582 | ~v_136;
assign x_19606 = v_2582 | ~v_135;
assign x_19607 = v_2582 | ~v_1249;
assign x_19608 = v_2582 | ~v_993;
assign x_19609 = v_2582 | ~v_1250;
assign x_19610 = v_2582 | ~v_994;
assign x_19611 = v_2582 | ~v_18;
assign x_19612 = v_2582 | ~v_17;
assign x_19613 = v_2582 | ~v_16;
assign x_19614 = v_2582 | ~v_15;
assign x_19615 = v_2582 | ~v_14;
assign x_19616 = v_2582 | ~v_13;
assign x_19617 = v_2582 | ~v_10;
assign x_19618 = ~v_2580 | ~v_2579 | ~v_2578 | v_2581;
assign x_19619 = v_2580 | ~v_2438;
assign x_19620 = v_2580 | ~v_2439;
assign x_19621 = v_2580 | ~v_2440;
assign x_19622 = v_2580 | ~v_2441;
assign x_19623 = v_2580 | ~v_1822;
assign x_19624 = v_2580 | ~v_1823;
assign x_19625 = v_2580 | ~v_1824;
assign x_19626 = v_2580 | ~v_1825;
assign x_19627 = v_2580 | ~v_1626;
assign x_19628 = v_2580 | ~v_1746;
assign x_19629 = v_2580 | ~v_1747;
assign x_19630 = v_2580 | ~v_1629;
assign x_19631 = v_2580 | ~v_1748;
assign x_19632 = v_2580 | ~v_1749;
assign x_19633 = v_2580 | ~v_885;
assign x_19634 = v_2580 | ~v_1019;
assign x_19635 = v_2580 | ~v_1020;
assign x_19636 = v_2580 | ~v_886;
assign x_19637 = v_2580 | ~v_1021;
assign x_19638 = v_2580 | ~v_1022;
assign x_19639 = v_2580 | ~v_2564;
assign x_19640 = v_2580 | ~v_2565;
assign x_19641 = v_2580 | ~v_2566;
assign x_19642 = v_2580 | ~v_2567;
assign x_19643 = v_2580 | ~v_1023;
assign x_19644 = v_2580 | ~v_1024;
assign x_19645 = v_2580 | ~v_2446;
assign x_19646 = v_2580 | ~v_2512;
assign x_19647 = v_2580 | ~v_2513;
assign x_19648 = v_2580 | ~v_2449;
assign x_19649 = v_2580 | ~v_2514;
assign x_19650 = v_2580 | ~v_2515;
assign x_19651 = v_2580 | ~v_184;
assign x_19652 = v_2580 | ~v_181;
assign x_19653 = v_2580 | ~v_171;
assign x_19654 = v_2580 | ~v_170;
assign x_19655 = v_2580 | ~v_149;
assign x_19656 = v_2580 | ~v_148;
assign x_19657 = v_2580 | ~v_147;
assign x_19658 = v_2580 | ~v_103;
assign x_19659 = v_2580 | ~v_102;
assign x_19660 = v_2580 | ~v_101;
assign x_19661 = v_2580 | ~v_99;
assign x_19662 = v_2580 | ~v_93;
assign x_19663 = v_2579 | ~v_2423;
assign x_19664 = v_2579 | ~v_2424;
assign x_19665 = v_2579 | ~v_2425;
assign x_19666 = v_2579 | ~v_2426;
assign x_19667 = v_2579 | ~v_1813;
assign x_19668 = v_2579 | ~v_1814;
assign x_19669 = v_2579 | ~v_1815;
assign x_19670 = v_2579 | ~v_1816;
assign x_19671 = v_2579 | ~v_1601;
assign x_19672 = v_2579 | ~v_1737;
assign x_19673 = v_2579 | ~v_1738;
assign x_19674 = v_2579 | ~v_1604;
assign x_19675 = v_2579 | ~v_1739;
assign x_19676 = v_2579 | ~v_1740;
assign x_19677 = v_2579 | ~v_870;
assign x_19678 = v_2579 | ~v_1004;
assign x_19679 = v_2579 | ~v_1005;
assign x_19680 = v_2579 | ~v_871;
assign x_19681 = v_2579 | ~v_1006;
assign x_19682 = v_2579 | ~v_1007;
assign x_19683 = v_2579 | ~v_2559;
assign x_19684 = v_2579 | ~v_2560;
assign x_19685 = v_2579 | ~v_2561;
assign x_19686 = v_2579 | ~v_2562;
assign x_19687 = v_2579 | ~v_1008;
assign x_19688 = v_2579 | ~v_1009;
assign x_19689 = v_2579 | ~v_2431;
assign x_19690 = v_2579 | ~v_2507;
assign x_19691 = v_2579 | ~v_2508;
assign x_19692 = v_2579 | ~v_2434;
assign x_19693 = v_2579 | ~v_2509;
assign x_19694 = v_2579 | ~v_2510;
assign x_19695 = v_2579 | ~v_183;
assign x_19696 = v_2579 | ~v_180;
assign x_19697 = v_2579 | ~v_167;
assign x_19698 = v_2579 | ~v_166;
assign x_19699 = v_2579 | ~v_144;
assign x_19700 = v_2579 | ~v_143;
assign x_19701 = v_2579 | ~v_142;
assign x_19702 = v_2579 | ~v_61;
assign x_19703 = v_2579 | ~v_60;
assign x_19704 = v_2579 | ~v_59;
assign x_19705 = v_2579 | ~v_57;
assign x_19706 = v_2579 | ~v_51;
assign x_19707 = v_2578 | ~v_2408;
assign x_19708 = v_2578 | ~v_2409;
assign x_19709 = v_2578 | ~v_2410;
assign x_19710 = v_2578 | ~v_2411;
assign x_19711 = v_2578 | ~v_1804;
assign x_19712 = v_2578 | ~v_1805;
assign x_19713 = v_2578 | ~v_1806;
assign x_19714 = v_2578 | ~v_1807;
assign x_19715 = v_2578 | ~v_1576;
assign x_19716 = v_2578 | ~v_1728;
assign x_19717 = v_2578 | ~v_1729;
assign x_19718 = v_2578 | ~v_1579;
assign x_19719 = v_2578 | ~v_1730;
assign x_19720 = v_2578 | ~v_1731;
assign x_19721 = v_2578 | ~v_855;
assign x_19722 = v_2578 | ~v_989;
assign x_19723 = v_2578 | ~v_990;
assign x_19724 = v_2578 | ~v_856;
assign x_19725 = v_2578 | ~v_991;
assign x_19726 = v_2578 | ~v_992;
assign x_19727 = v_2578 | ~v_2554;
assign x_19728 = v_2578 | ~v_2555;
assign x_19729 = v_2578 | ~v_2556;
assign x_19730 = v_2578 | ~v_2557;
assign x_19731 = v_2578 | ~v_2416;
assign x_19732 = v_2578 | ~v_2502;
assign x_19733 = v_2578 | ~v_2503;
assign x_19734 = v_2578 | ~v_2419;
assign x_19735 = v_2578 | ~v_2504;
assign x_19736 = v_2578 | ~v_2505;
assign x_19737 = v_2578 | ~v_182;
assign x_19738 = v_2578 | ~v_179;
assign x_19739 = v_2578 | ~v_163;
assign x_19740 = v_2578 | ~v_162;
assign x_19741 = v_2578 | ~v_136;
assign x_19742 = v_2578 | ~v_135;
assign x_19743 = v_2578 | ~v_134;
assign x_19744 = v_2578 | ~v_993;
assign x_19745 = v_2578 | ~v_994;
assign x_19746 = v_2578 | ~v_18;
assign x_19747 = v_2578 | ~v_17;
assign x_19748 = v_2578 | ~v_16;
assign x_19749 = v_2578 | ~v_14;
assign x_19750 = v_2578 | ~v_8;
assign x_19751 = ~v_2576 | ~v_2575 | ~v_2574 | v_2577;
assign x_19752 = v_2576 | ~v_2438;
assign x_19753 = v_2576 | ~v_2439;
assign x_19754 = v_2576 | ~v_2440;
assign x_19755 = v_2576 | ~v_2441;
assign x_19756 = v_2576 | ~v_1718;
assign x_19757 = v_2576 | ~v_1719;
assign x_19758 = v_2576 | ~v_1720;
assign x_19759 = v_2576 | ~v_1721;
assign x_19760 = v_2576 | ~v_1822;
assign x_19761 = v_2576 | ~v_1823;
assign x_19762 = v_2576 | ~v_1824;
assign x_19763 = v_2576 | ~v_1825;
assign x_19764 = v_2576 | ~v_1626;
assign x_19765 = v_2576 | ~v_1629;
assign x_19766 = v_2576 | ~v_881;
assign x_19767 = v_2576 | ~v_882;
assign x_19768 = v_2576 | ~v_883;
assign x_19769 = v_2576 | ~v_884;
assign x_19770 = v_2576 | ~v_885;
assign x_19771 = v_2576 | ~v_886;
assign x_19772 = v_2576 | ~v_2564;
assign x_19773 = v_2576 | ~v_2565;
assign x_19774 = v_2576 | ~v_2566;
assign x_19775 = v_2576 | ~v_2567;
assign x_19776 = v_2576 | ~v_837;
assign x_19777 = v_2576 | ~v_838;
assign x_19778 = v_2576 | ~v_2496;
assign x_19779 = v_2576 | ~v_2497;
assign x_19780 = v_2576 | ~v_2498;
assign x_19781 = v_2576 | ~v_2499;
assign x_19782 = v_2576 | ~v_2446;
assign x_19783 = v_2576 | ~v_2449;
assign x_19784 = v_2576 | ~v_184;
assign x_19785 = v_2576 | ~v_181;
assign x_19786 = v_2576 | ~v_171;
assign x_19787 = v_2576 | ~v_170;
assign x_19788 = v_2576 | ~v_160;
assign x_19789 = v_2576 | ~v_150;
assign x_19790 = v_2576 | ~v_149;
assign x_19791 = v_2576 | ~v_103;
assign x_19792 = v_2576 | ~v_102;
assign x_19793 = v_2576 | ~v_96;
assign x_19794 = v_2576 | ~v_95;
assign x_19795 = v_2576 | ~v_93;
assign x_19796 = v_2575 | ~v_2423;
assign x_19797 = v_2575 | ~v_2424;
assign x_19798 = v_2575 | ~v_2425;
assign x_19799 = v_2575 | ~v_2426;
assign x_19800 = v_2575 | ~v_1709;
assign x_19801 = v_2575 | ~v_1710;
assign x_19802 = v_2575 | ~v_1711;
assign x_19803 = v_2575 | ~v_1712;
assign x_19804 = v_2575 | ~v_1813;
assign x_19805 = v_2575 | ~v_1814;
assign x_19806 = v_2575 | ~v_1815;
assign x_19807 = v_2575 | ~v_1816;
assign x_19808 = v_2575 | ~v_1601;
assign x_19809 = v_2575 | ~v_1604;
assign x_19810 = v_2575 | ~v_866;
assign x_19811 = v_2575 | ~v_867;
assign x_19812 = v_2575 | ~v_868;
assign x_19813 = v_2575 | ~v_869;
assign x_19814 = v_2575 | ~v_870;
assign x_19815 = v_2575 | ~v_871;
assign x_19816 = v_2575 | ~v_2559;
assign x_19817 = v_2575 | ~v_2560;
assign x_19818 = v_2575 | ~v_2561;
assign x_19819 = v_2575 | ~v_2562;
assign x_19820 = v_2575 | ~v_804;
assign x_19821 = v_2575 | ~v_805;
assign x_19822 = v_2575 | ~v_2491;
assign x_19823 = v_2575 | ~v_2492;
assign x_19824 = v_2575 | ~v_2493;
assign x_19825 = v_2575 | ~v_2494;
assign x_19826 = v_2575 | ~v_2431;
assign x_19827 = v_2575 | ~v_2434;
assign x_19828 = v_2575 | ~v_183;
assign x_19829 = v_2575 | ~v_180;
assign x_19830 = v_2575 | ~v_167;
assign x_19831 = v_2575 | ~v_166;
assign x_19832 = v_2575 | ~v_159;
assign x_19833 = v_2575 | ~v_145;
assign x_19834 = v_2575 | ~v_144;
assign x_19835 = v_2575 | ~v_61;
assign x_19836 = v_2575 | ~v_60;
assign x_19837 = v_2575 | ~v_54;
assign x_19838 = v_2575 | ~v_53;
assign x_19839 = v_2575 | ~v_51;
assign x_19840 = v_2574 | ~v_2408;
assign x_19841 = v_2574 | ~v_2409;
assign x_19842 = v_2574 | ~v_2410;
assign x_19843 = v_2574 | ~v_2411;
assign x_19844 = v_2574 | ~v_1700;
assign x_19845 = v_2574 | ~v_1701;
assign x_19846 = v_2574 | ~v_1702;
assign x_19847 = v_2574 | ~v_1703;
assign x_19848 = v_2574 | ~v_1804;
assign x_19849 = v_2574 | ~v_1805;
assign x_19850 = v_2574 | ~v_1806;
assign x_19851 = v_2574 | ~v_1807;
assign x_19852 = v_2574 | ~v_1576;
assign x_19853 = v_2574 | ~v_1579;
assign x_19854 = v_2574 | ~v_851;
assign x_19855 = v_2574 | ~v_852;
assign x_19856 = v_2574 | ~v_853;
assign x_19857 = v_2574 | ~v_854;
assign x_19858 = v_2574 | ~v_855;
assign x_19859 = v_2574 | ~v_856;
assign x_19860 = v_2574 | ~v_2554;
assign x_19861 = v_2574 | ~v_2555;
assign x_19862 = v_2574 | ~v_2556;
assign x_19863 = v_2574 | ~v_2557;
assign x_19864 = v_2574 | ~v_771;
assign x_19865 = v_2574 | ~v_772;
assign x_19866 = v_2574 | ~v_2486;
assign x_19867 = v_2574 | ~v_2487;
assign x_19868 = v_2574 | ~v_2488;
assign x_19869 = v_2574 | ~v_2489;
assign x_19870 = v_2574 | ~v_2416;
assign x_19871 = v_2574 | ~v_2419;
assign x_19872 = v_2574 | ~v_182;
assign x_19873 = v_2574 | ~v_179;
assign x_19874 = v_2574 | ~v_163;
assign x_19875 = v_2574 | ~v_162;
assign x_19876 = v_2574 | ~v_155;
assign x_19877 = v_2574 | ~v_137;
assign x_19878 = v_2574 | ~v_136;
assign x_19879 = v_2574 | ~v_18;
assign x_19880 = v_2574 | ~v_17;
assign x_19881 = v_2574 | ~v_11;
assign x_19882 = v_2574 | ~v_10;
assign x_19883 = v_2574 | ~v_8;
assign x_19884 = ~v_2572 | ~v_2571 | ~v_2570 | v_2573;
assign x_19885 = v_2572 | ~v_2438;
assign x_19886 = v_2572 | ~v_2439;
assign x_19887 = v_2572 | ~v_2440;
assign x_19888 = v_2572 | ~v_2441;
assign x_19889 = v_2572 | ~v_1690;
assign x_19890 = v_2572 | ~v_1691;
assign x_19891 = v_2572 | ~v_1692;
assign x_19892 = v_2572 | ~v_1693;
assign x_19893 = v_2572 | ~v_1822;
assign x_19894 = v_2572 | ~v_1823;
assign x_19895 = v_2572 | ~v_1824;
assign x_19896 = v_2572 | ~v_1825;
assign x_19897 = v_2572 | ~v_1626;
assign x_19898 = v_2572 | ~v_1629;
assign x_19899 = v_2572 | ~v_925;
assign x_19900 = v_2572 | ~v_926;
assign x_19901 = v_2572 | ~v_885;
assign x_19902 = v_2572 | ~v_886;
assign x_19903 = v_2572 | ~v_2564;
assign x_19904 = v_2572 | ~v_2565;
assign x_19905 = v_2572 | ~v_2566;
assign x_19906 = v_2572 | ~v_2567;
assign x_19907 = v_2572 | ~v_927;
assign x_19908 = v_2572 | ~v_928;
assign x_19909 = v_2572 | ~v_2480;
assign x_19910 = v_2572 | ~v_2481;
assign x_19911 = v_2572 | ~v_2482;
assign x_19912 = v_2572 | ~v_2483;
assign x_19913 = v_2572 | ~v_2446;
assign x_19914 = v_2572 | ~v_2449;
assign x_19915 = v_2572 | ~v_929;
assign x_19916 = v_2572 | ~v_930;
assign x_19917 = v_2572 | ~v_184;
assign x_19918 = v_2572 | ~v_181;
assign x_19919 = v_2572 | ~v_171;
assign x_19920 = v_2572 | ~v_170;
assign x_19921 = v_2572 | ~v_150;
assign x_19922 = v_2572 | ~v_148;
assign x_19923 = v_2572 | ~v_147;
assign x_19924 = v_2572 | ~v_103;
assign x_19925 = v_2572 | ~v_102;
assign x_19926 = v_2572 | ~v_101;
assign x_19927 = v_2572 | ~v_97;
assign x_19928 = v_2572 | ~v_93;
assign x_19929 = v_2571 | ~v_2423;
assign x_19930 = v_2571 | ~v_2424;
assign x_19931 = v_2571 | ~v_2425;
assign x_19932 = v_2571 | ~v_2426;
assign x_19933 = v_2571 | ~v_1681;
assign x_19934 = v_2571 | ~v_1682;
assign x_19935 = v_2571 | ~v_1683;
assign x_19936 = v_2571 | ~v_1684;
assign x_19937 = v_2571 | ~v_1813;
assign x_19938 = v_2571 | ~v_1814;
assign x_19939 = v_2571 | ~v_1815;
assign x_19940 = v_2571 | ~v_1816;
assign x_19941 = v_2571 | ~v_1601;
assign x_19942 = v_2571 | ~v_1604;
assign x_19943 = v_2571 | ~v_910;
assign x_19944 = v_2571 | ~v_911;
assign x_19945 = v_2571 | ~v_870;
assign x_19946 = v_2571 | ~v_871;
assign x_19947 = v_2571 | ~v_2559;
assign x_19948 = v_2571 | ~v_2560;
assign x_19949 = v_2571 | ~v_2561;
assign x_19950 = v_2571 | ~v_2562;
assign x_19951 = v_2571 | ~v_912;
assign x_19952 = v_2571 | ~v_913;
assign x_19953 = v_2571 | ~v_2475;
assign x_19954 = v_2571 | ~v_2476;
assign x_19955 = v_2571 | ~v_2477;
assign x_19956 = v_2571 | ~v_2478;
assign x_19957 = v_2571 | ~v_2431;
assign x_19958 = v_2571 | ~v_2434;
assign x_19959 = v_2571 | ~v_914;
assign x_19960 = v_2571 | ~v_915;
assign x_19961 = v_2571 | ~v_183;
assign x_19962 = v_2571 | ~v_180;
assign x_19963 = v_2571 | ~v_167;
assign x_19964 = v_2571 | ~v_166;
assign x_19965 = v_2571 | ~v_145;
assign x_19966 = v_2571 | ~v_143;
assign x_19967 = v_2571 | ~v_142;
assign x_19968 = v_2571 | ~v_61;
assign x_19969 = v_2571 | ~v_60;
assign x_19970 = v_2571 | ~v_59;
assign x_19971 = v_2571 | ~v_55;
assign x_19972 = v_2571 | ~v_51;
assign x_19973 = v_2570 | ~v_2408;
assign x_19974 = v_2570 | ~v_2409;
assign x_19975 = v_2570 | ~v_2410;
assign x_19976 = v_2570 | ~v_2411;
assign x_19977 = v_2570 | ~v_1672;
assign x_19978 = v_2570 | ~v_1673;
assign x_19979 = v_2570 | ~v_1674;
assign x_19980 = v_2570 | ~v_1675;
assign x_19981 = v_2570 | ~v_1804;
assign x_19982 = v_2570 | ~v_1805;
assign x_19983 = v_2570 | ~v_1806;
assign x_19984 = v_2570 | ~v_1807;
assign x_19985 = v_2570 | ~v_1576;
assign x_19986 = v_2570 | ~v_1579;
assign x_19987 = v_2570 | ~v_895;
assign x_19988 = v_2570 | ~v_896;
assign x_19989 = v_2570 | ~v_855;
assign x_19990 = v_2570 | ~v_856;
assign x_19991 = v_2570 | ~v_2554;
assign x_19992 = v_2570 | ~v_2555;
assign x_19993 = v_2570 | ~v_2556;
assign x_19994 = v_2570 | ~v_2557;
assign x_19995 = v_2570 | ~v_897;
assign x_19996 = v_2570 | ~v_898;
assign x_19997 = v_2570 | ~v_2470;
assign x_19998 = v_2570 | ~v_2471;
assign x_19999 = v_2570 | ~v_2472;
assign x_20000 = v_2570 | ~v_2473;
assign x_20001 = v_2570 | ~v_2416;
assign x_20002 = v_2570 | ~v_2419;
assign x_20003 = v_2570 | ~v_899;
assign x_20004 = v_2570 | ~v_900;
assign x_20005 = v_2570 | ~v_182;
assign x_20006 = v_2570 | ~v_179;
assign x_20007 = v_2570 | ~v_163;
assign x_20008 = v_2570 | ~v_162;
assign x_20009 = v_2570 | ~v_137;
assign x_20010 = v_2570 | ~v_135;
assign x_20011 = v_2570 | ~v_134;
assign x_20012 = v_2570 | ~v_18;
assign x_20013 = v_2570 | ~v_17;
assign x_20014 = v_2570 | ~v_16;
assign x_20015 = v_2570 | ~v_12;
assign x_20016 = v_2570 | ~v_8;
assign x_20017 = ~v_2568 | ~v_2563 | ~v_2558 | v_2569;
assign x_20018 = v_2568 | ~v_2438;
assign x_20019 = v_2568 | ~v_2439;
assign x_20020 = v_2568 | ~v_2440;
assign x_20021 = v_2568 | ~v_2441;
assign x_20022 = v_2568 | ~v_1622;
assign x_20023 = v_2568 | ~v_1623;
assign x_20024 = v_2568 | ~v_1624;
assign x_20025 = v_2568 | ~v_1625;
assign x_20026 = v_2568 | ~v_1822;
assign x_20027 = v_2568 | ~v_1823;
assign x_20028 = v_2568 | ~v_1824;
assign x_20029 = v_2568 | ~v_1825;
assign x_20030 = v_2568 | ~v_1626;
assign x_20031 = v_2568 | ~v_1629;
assign x_20032 = v_2568 | ~v_973;
assign x_20033 = v_2568 | ~v_974;
assign x_20034 = v_2568 | ~v_885;
assign x_20035 = v_2568 | ~v_886;
assign x_20036 = v_2568 | ~v_2564;
assign x_20037 = v_2568 | ~v_2565;
assign x_20038 = v_2568 | ~v_2566;
assign x_20039 = v_2568 | ~v_2567;
assign x_20040 = v_2568 | ~v_975;
assign x_20041 = v_2568 | ~v_976;
assign x_20042 = v_2568 | ~v_2442;
assign x_20043 = v_2568 | ~v_2443;
assign x_20044 = v_2568 | ~v_2444;
assign x_20045 = v_2568 | ~v_2445;
assign x_20046 = v_2568 | ~v_2446;
assign x_20047 = v_2568 | ~v_2449;
assign x_20048 = v_2568 | ~v_977;
assign x_20049 = v_2568 | ~v_978;
assign x_20050 = v_2568 | ~v_184;
assign x_20051 = v_2568 | ~v_181;
assign x_20052 = v_2568 | ~v_172;
assign x_20053 = v_2568 | ~v_171;
assign x_20054 = v_2568 | ~v_170;
assign x_20055 = v_2568 | ~v_150;
assign x_20056 = v_2568 | ~v_149;
assign x_20057 = v_2568 | ~v_148;
assign x_20058 = v_2568 | ~v_147;
assign x_20059 = v_2568 | ~v_102;
assign x_20060 = v_2568 | ~v_101;
assign x_20061 = v_2568 | ~v_93;
assign x_20062 = ~v_128 | ~v_176 | v_2567;
assign x_20063 = ~v_125 | ~v_175 | v_2566;
assign x_20064 = ~v_113 | v_176 | v_2565;
assign x_20065 = ~v_110 | v_175 | v_2564;
assign x_20066 = v_2563 | ~v_2423;
assign x_20067 = v_2563 | ~v_2424;
assign x_20068 = v_2563 | ~v_2425;
assign x_20069 = v_2563 | ~v_2426;
assign x_20070 = v_2563 | ~v_1597;
assign x_20071 = v_2563 | ~v_1598;
assign x_20072 = v_2563 | ~v_1599;
assign x_20073 = v_2563 | ~v_1600;
assign x_20074 = v_2563 | ~v_1813;
assign x_20075 = v_2563 | ~v_1814;
assign x_20076 = v_2563 | ~v_1815;
assign x_20077 = v_2563 | ~v_1816;
assign x_20078 = v_2563 | ~v_1601;
assign x_20079 = v_2563 | ~v_1604;
assign x_20080 = v_2563 | ~v_958;
assign x_20081 = v_2563 | ~v_959;
assign x_20082 = v_2563 | ~v_870;
assign x_20083 = v_2563 | ~v_871;
assign x_20084 = v_2563 | ~v_2559;
assign x_20085 = v_2563 | ~v_2560;
assign x_20086 = v_2563 | ~v_2561;
assign x_20087 = v_2563 | ~v_2562;
assign x_20088 = v_2563 | ~v_960;
assign x_20089 = v_2563 | ~v_961;
assign x_20090 = v_2563 | ~v_2427;
assign x_20091 = v_2563 | ~v_2428;
assign x_20092 = v_2563 | ~v_2429;
assign x_20093 = v_2563 | ~v_2430;
assign x_20094 = v_2563 | ~v_2431;
assign x_20095 = v_2563 | ~v_2434;
assign x_20096 = v_2563 | ~v_962;
assign x_20097 = v_2563 | ~v_963;
assign x_20098 = v_2563 | ~v_183;
assign x_20099 = v_2563 | ~v_180;
assign x_20100 = v_2563 | ~v_168;
assign x_20101 = v_2563 | ~v_167;
assign x_20102 = v_2563 | ~v_166;
assign x_20103 = v_2563 | ~v_145;
assign x_20104 = v_2563 | ~v_144;
assign x_20105 = v_2563 | ~v_143;
assign x_20106 = v_2563 | ~v_142;
assign x_20107 = v_2563 | ~v_60;
assign x_20108 = v_2563 | ~v_59;
assign x_20109 = v_2563 | ~v_51;
assign x_20110 = ~v_86 | ~v_176 | v_2562;
assign x_20111 = ~v_83 | ~v_175 | v_2561;
assign x_20112 = ~v_71 | v_176 | v_2560;
assign x_20113 = ~v_68 | v_175 | v_2559;
assign x_20114 = v_2558 | ~v_2408;
assign x_20115 = v_2558 | ~v_2409;
assign x_20116 = v_2558 | ~v_2410;
assign x_20117 = v_2558 | ~v_2411;
assign x_20118 = v_2558 | ~v_1572;
assign x_20119 = v_2558 | ~v_1573;
assign x_20120 = v_2558 | ~v_1574;
assign x_20121 = v_2558 | ~v_1575;
assign x_20122 = v_2558 | ~v_1804;
assign x_20123 = v_2558 | ~v_1805;
assign x_20124 = v_2558 | ~v_1806;
assign x_20125 = v_2558 | ~v_1807;
assign x_20126 = v_2558 | ~v_1576;
assign x_20127 = v_2558 | ~v_1579;
assign x_20128 = v_2558 | ~v_943;
assign x_20129 = v_2558 | ~v_944;
assign x_20130 = v_2558 | ~v_855;
assign x_20131 = v_2558 | ~v_856;
assign x_20132 = v_2558 | ~v_2554;
assign x_20133 = v_2558 | ~v_2555;
assign x_20134 = v_2558 | ~v_2556;
assign x_20135 = v_2558 | ~v_2557;
assign x_20136 = v_2558 | ~v_945;
assign x_20137 = v_2558 | ~v_946;
assign x_20138 = v_2558 | ~v_2412;
assign x_20139 = v_2558 | ~v_2413;
assign x_20140 = v_2558 | ~v_2414;
assign x_20141 = v_2558 | ~v_2415;
assign x_20142 = v_2558 | ~v_2416;
assign x_20143 = v_2558 | ~v_2419;
assign x_20144 = v_2558 | ~v_947;
assign x_20145 = v_2558 | ~v_948;
assign x_20146 = v_2558 | ~v_182;
assign x_20147 = v_2558 | ~v_179;
assign x_20148 = v_2558 | ~v_164;
assign x_20149 = v_2558 | ~v_163;
assign x_20150 = v_2558 | ~v_162;
assign x_20151 = v_2558 | ~v_137;
assign x_20152 = v_2558 | ~v_136;
assign x_20153 = v_2558 | ~v_135;
assign x_20154 = v_2558 | ~v_134;
assign x_20155 = v_2558 | ~v_17;
assign x_20156 = v_2558 | ~v_16;
assign x_20157 = v_2558 | ~v_8;
assign x_20158 = ~v_44 | ~v_176 | v_2557;
assign x_20159 = ~v_41 | ~v_175 | v_2556;
assign x_20160 = ~v_29 | v_176 | v_2555;
assign x_20161 = ~v_26 | v_175 | v_2554;
assign x_20162 = ~v_2552 | ~v_2551 | ~v_2550 | v_2553;
assign x_20163 = v_2552 | ~v_2438;
assign x_20164 = v_2552 | ~v_2439;
assign x_20165 = v_2552 | ~v_2440;
assign x_20166 = v_2552 | ~v_2441;
assign x_20167 = v_2552 | ~v_1718;
assign x_20168 = v_2552 | ~v_1719;
assign x_20169 = v_2552 | ~v_1720;
assign x_20170 = v_2552 | ~v_1721;
assign x_20171 = v_2552 | ~v_1626;
assign x_20172 = v_2552 | ~v_1627;
assign x_20173 = v_2552 | ~v_1628;
assign x_20174 = v_2552 | ~v_1629;
assign x_20175 = v_2552 | ~v_1630;
assign x_20176 = v_2552 | ~v_1631;
assign x_20177 = v_2552 | ~v_833;
assign x_20178 = v_2552 | ~v_834;
assign x_20179 = v_2552 | ~v_835;
assign x_20180 = v_2552 | ~v_836;
assign x_20181 = v_2552 | ~v_837;
assign x_20182 = v_2552 | ~v_838;
assign x_20183 = v_2552 | ~v_2496;
assign x_20184 = v_2552 | ~v_2497;
assign x_20185 = v_2552 | ~v_2498;
assign x_20186 = v_2552 | ~v_2499;
assign x_20187 = v_2552 | ~v_839;
assign x_20188 = v_2552 | ~v_840;
assign x_20189 = v_2552 | ~v_2446;
assign x_20190 = v_2552 | ~v_2447;
assign x_20191 = v_2552 | ~v_2448;
assign x_20192 = v_2552 | ~v_2449;
assign x_20193 = v_2552 | ~v_2450;
assign x_20194 = v_2552 | ~v_2451;
assign x_20195 = v_2552 | ~v_184;
assign x_20196 = v_2552 | ~v_170;
assign x_20197 = v_2552 | ~v_169;
assign x_20198 = v_2552 | ~v_160;
assign x_20199 = v_2552 | ~v_150;
assign x_20200 = v_2552 | ~v_149;
assign x_20201 = v_2552 | ~v_147;
assign x_20202 = v_2552 | ~v_103;
assign x_20203 = v_2552 | ~v_102;
assign x_20204 = v_2552 | ~v_100;
assign x_20205 = v_2552 | ~v_98;
assign x_20206 = v_2552 | ~v_96;
assign x_20207 = v_2551 | ~v_2423;
assign x_20208 = v_2551 | ~v_2424;
assign x_20209 = v_2551 | ~v_2425;
assign x_20210 = v_2551 | ~v_2426;
assign x_20211 = v_2551 | ~v_1709;
assign x_20212 = v_2551 | ~v_1710;
assign x_20213 = v_2551 | ~v_1711;
assign x_20214 = v_2551 | ~v_1712;
assign x_20215 = v_2551 | ~v_1601;
assign x_20216 = v_2551 | ~v_1602;
assign x_20217 = v_2551 | ~v_1603;
assign x_20218 = v_2551 | ~v_1604;
assign x_20219 = v_2551 | ~v_1605;
assign x_20220 = v_2551 | ~v_1606;
assign x_20221 = v_2551 | ~v_800;
assign x_20222 = v_2551 | ~v_801;
assign x_20223 = v_2551 | ~v_802;
assign x_20224 = v_2551 | ~v_803;
assign x_20225 = v_2551 | ~v_804;
assign x_20226 = v_2551 | ~v_805;
assign x_20227 = v_2551 | ~v_2491;
assign x_20228 = v_2551 | ~v_2492;
assign x_20229 = v_2551 | ~v_2493;
assign x_20230 = v_2551 | ~v_2494;
assign x_20231 = v_2551 | ~v_806;
assign x_20232 = v_2551 | ~v_2431;
assign x_20233 = v_2551 | ~v_2432;
assign x_20234 = v_2551 | ~v_2433;
assign x_20235 = v_2551 | ~v_2434;
assign x_20236 = v_2551 | ~v_2435;
assign x_20237 = v_2551 | ~v_2436;
assign x_20238 = v_2551 | ~v_807;
assign x_20239 = v_2551 | ~v_183;
assign x_20240 = v_2551 | ~v_166;
assign x_20241 = v_2551 | ~v_165;
assign x_20242 = v_2551 | ~v_159;
assign x_20243 = v_2551 | ~v_145;
assign x_20244 = v_2551 | ~v_144;
assign x_20245 = v_2551 | ~v_142;
assign x_20246 = v_2551 | ~v_61;
assign x_20247 = v_2551 | ~v_60;
assign x_20248 = v_2551 | ~v_58;
assign x_20249 = v_2551 | ~v_56;
assign x_20250 = v_2551 | ~v_54;
assign x_20251 = v_2550 | ~v_2408;
assign x_20252 = v_2550 | ~v_2409;
assign x_20253 = v_2550 | ~v_2410;
assign x_20254 = v_2550 | ~v_2411;
assign x_20255 = v_2550 | ~v_1700;
assign x_20256 = v_2550 | ~v_1701;
assign x_20257 = v_2550 | ~v_1702;
assign x_20258 = v_2550 | ~v_1703;
assign x_20259 = v_2550 | ~v_1576;
assign x_20260 = v_2550 | ~v_1577;
assign x_20261 = v_2550 | ~v_1578;
assign x_20262 = v_2550 | ~v_1579;
assign x_20263 = v_2550 | ~v_1580;
assign x_20264 = v_2550 | ~v_1581;
assign x_20265 = v_2550 | ~v_767;
assign x_20266 = v_2550 | ~v_768;
assign x_20267 = v_2550 | ~v_769;
assign x_20268 = v_2550 | ~v_770;
assign x_20269 = v_2550 | ~v_771;
assign x_20270 = v_2550 | ~v_772;
assign x_20271 = v_2550 | ~v_2486;
assign x_20272 = v_2550 | ~v_2487;
assign x_20273 = v_2550 | ~v_2488;
assign x_20274 = v_2550 | ~v_2489;
assign x_20275 = v_2550 | ~v_773;
assign x_20276 = v_2550 | ~v_774;
assign x_20277 = v_2550 | ~v_2416;
assign x_20278 = v_2550 | ~v_2417;
assign x_20279 = v_2550 | ~v_2418;
assign x_20280 = v_2550 | ~v_2419;
assign x_20281 = v_2550 | ~v_2420;
assign x_20282 = v_2550 | ~v_2421;
assign x_20283 = v_2550 | ~v_182;
assign x_20284 = v_2550 | ~v_162;
assign x_20285 = v_2550 | ~v_161;
assign x_20286 = v_2550 | ~v_155;
assign x_20287 = v_2550 | ~v_137;
assign x_20288 = v_2550 | ~v_136;
assign x_20289 = v_2550 | ~v_134;
assign x_20290 = v_2550 | ~v_18;
assign x_20291 = v_2550 | ~v_17;
assign x_20292 = v_2550 | ~v_15;
assign x_20293 = v_2550 | ~v_13;
assign x_20294 = v_2550 | ~v_11;
assign x_20295 = ~v_2548 | ~v_2547 | ~v_2546 | v_2549;
assign x_20296 = v_2548 | ~v_2438;
assign x_20297 = v_2548 | ~v_2439;
assign x_20298 = v_2548 | ~v_2440;
assign x_20299 = v_2548 | ~v_2441;
assign x_20300 = v_2548 | ~v_1778;
assign x_20301 = v_2548 | ~v_1779;
assign x_20302 = v_2548 | ~v_1780;
assign x_20303 = v_2548 | ~v_1781;
assign x_20304 = v_2548 | ~v_1626;
assign x_20305 = v_2548 | ~v_1746;
assign x_20306 = v_2548 | ~v_1747;
assign x_20307 = v_2548 | ~v_1629;
assign x_20308 = v_2548 | ~v_1748;
assign x_20309 = v_2548 | ~v_1749;
assign x_20310 = v_2548 | ~v_1085;
assign x_20311 = v_2548 | ~v_1131;
assign x_20312 = v_2548 | ~v_1132;
assign x_20313 = v_2548 | ~v_1086;
assign x_20314 = v_2548 | ~v_1133;
assign x_20315 = v_2548 | ~v_1134;
assign x_20316 = v_2548 | ~v_2532;
assign x_20317 = v_2548 | ~v_2533;
assign x_20318 = v_2548 | ~v_2534;
assign x_20319 = v_2548 | ~v_2535;
assign x_20320 = v_2548 | ~v_1023;
assign x_20321 = v_2548 | ~v_1024;
assign x_20322 = v_2548 | ~v_2446;
assign x_20323 = v_2548 | ~v_2512;
assign x_20324 = v_2548 | ~v_2513;
assign x_20325 = v_2548 | ~v_2449;
assign x_20326 = v_2548 | ~v_2514;
assign x_20327 = v_2548 | ~v_2515;
assign x_20328 = v_2548 | ~v_184;
assign x_20329 = v_2548 | ~v_172;
assign x_20330 = v_2548 | ~v_171;
assign x_20331 = v_2548 | ~v_169;
assign x_20332 = v_2548 | ~v_149;
assign x_20333 = v_2548 | ~v_148;
assign x_20334 = v_2548 | ~v_147;
assign x_20335 = v_2548 | ~v_102;
assign x_20336 = v_2548 | ~v_101;
assign x_20337 = v_2548 | ~v_100;
assign x_20338 = v_2548 | ~v_99;
assign x_20339 = v_2548 | ~v_94;
assign x_20340 = v_2547 | ~v_2423;
assign x_20341 = v_2547 | ~v_2424;
assign x_20342 = v_2547 | ~v_2425;
assign x_20343 = v_2547 | ~v_2426;
assign x_20344 = v_2547 | ~v_1769;
assign x_20345 = v_2547 | ~v_1770;
assign x_20346 = v_2547 | ~v_1771;
assign x_20347 = v_2547 | ~v_1772;
assign x_20348 = v_2547 | ~v_1601;
assign x_20349 = v_2547 | ~v_1737;
assign x_20350 = v_2547 | ~v_1738;
assign x_20351 = v_2547 | ~v_1604;
assign x_20352 = v_2547 | ~v_1739;
assign x_20353 = v_2547 | ~v_1740;
assign x_20354 = v_2547 | ~v_1070;
assign x_20355 = v_2547 | ~v_1126;
assign x_20356 = v_2547 | ~v_1127;
assign x_20357 = v_2547 | ~v_1071;
assign x_20358 = v_2547 | ~v_1128;
assign x_20359 = v_2547 | ~v_1129;
assign x_20360 = v_2547 | ~v_2527;
assign x_20361 = v_2547 | ~v_2528;
assign x_20362 = v_2547 | ~v_2529;
assign x_20363 = v_2547 | ~v_2530;
assign x_20364 = v_2547 | ~v_1008;
assign x_20365 = v_2547 | ~v_1009;
assign x_20366 = v_2547 | ~v_2431;
assign x_20367 = v_2547 | ~v_2507;
assign x_20368 = v_2547 | ~v_2508;
assign x_20369 = v_2547 | ~v_2434;
assign x_20370 = v_2547 | ~v_2509;
assign x_20371 = v_2547 | ~v_2510;
assign x_20372 = v_2547 | ~v_183;
assign x_20373 = v_2547 | ~v_168;
assign x_20374 = v_2547 | ~v_167;
assign x_20375 = v_2547 | ~v_165;
assign x_20376 = v_2547 | ~v_144;
assign x_20377 = v_2547 | ~v_143;
assign x_20378 = v_2547 | ~v_142;
assign x_20379 = v_2547 | ~v_60;
assign x_20380 = v_2547 | ~v_59;
assign x_20381 = v_2547 | ~v_58;
assign x_20382 = v_2547 | ~v_57;
assign x_20383 = v_2547 | ~v_52;
assign x_20384 = v_2546 | ~v_2408;
assign x_20385 = v_2546 | ~v_2409;
assign x_20386 = v_2546 | ~v_2410;
assign x_20387 = v_2546 | ~v_2411;
assign x_20388 = v_2546 | ~v_1760;
assign x_20389 = v_2546 | ~v_1761;
assign x_20390 = v_2546 | ~v_1762;
assign x_20391 = v_2546 | ~v_1763;
assign x_20392 = v_2546 | ~v_1576;
assign x_20393 = v_2546 | ~v_1728;
assign x_20394 = v_2546 | ~v_1729;
assign x_20395 = v_2546 | ~v_1579;
assign x_20396 = v_2546 | ~v_1730;
assign x_20397 = v_2546 | ~v_1731;
assign x_20398 = v_2546 | ~v_1055;
assign x_20399 = v_2546 | ~v_1121;
assign x_20400 = v_2546 | ~v_1122;
assign x_20401 = v_2546 | ~v_1056;
assign x_20402 = v_2546 | ~v_1123;
assign x_20403 = v_2546 | ~v_1124;
assign x_20404 = v_2546 | ~v_2522;
assign x_20405 = v_2546 | ~v_2523;
assign x_20406 = v_2546 | ~v_2524;
assign x_20407 = v_2546 | ~v_2525;
assign x_20408 = v_2546 | ~v_2416;
assign x_20409 = v_2546 | ~v_2502;
assign x_20410 = v_2546 | ~v_2503;
assign x_20411 = v_2546 | ~v_2419;
assign x_20412 = v_2546 | ~v_2504;
assign x_20413 = v_2546 | ~v_2505;
assign x_20414 = v_2546 | ~v_182;
assign x_20415 = v_2546 | ~v_164;
assign x_20416 = v_2546 | ~v_163;
assign x_20417 = v_2546 | ~v_161;
assign x_20418 = v_2546 | ~v_136;
assign x_20419 = v_2546 | ~v_135;
assign x_20420 = v_2546 | ~v_134;
assign x_20421 = v_2546 | ~v_993;
assign x_20422 = v_2546 | ~v_994;
assign x_20423 = v_2546 | ~v_17;
assign x_20424 = v_2546 | ~v_16;
assign x_20425 = v_2546 | ~v_15;
assign x_20426 = v_2546 | ~v_14;
assign x_20427 = v_2546 | ~v_9;
assign x_20428 = ~v_2544 | ~v_2543 | ~v_2542 | v_2545;
assign x_20429 = v_2544 | ~v_2438;
assign x_20430 = v_2544 | ~v_2439;
assign x_20431 = v_2544 | ~v_2440;
assign x_20432 = v_2544 | ~v_2441;
assign x_20433 = v_2544 | ~v_1778;
assign x_20434 = v_2544 | ~v_1779;
assign x_20435 = v_2544 | ~v_1780;
assign x_20436 = v_2544 | ~v_1781;
assign x_20437 = v_2544 | ~v_1718;
assign x_20438 = v_2544 | ~v_1719;
assign x_20439 = v_2544 | ~v_1720;
assign x_20440 = v_2544 | ~v_1721;
assign x_20441 = v_2544 | ~v_1626;
assign x_20442 = v_2544 | ~v_1629;
assign x_20443 = v_2544 | ~v_837;
assign x_20444 = v_2544 | ~v_838;
assign x_20445 = v_2544 | ~v_1081;
assign x_20446 = v_2544 | ~v_1082;
assign x_20447 = v_2544 | ~v_1083;
assign x_20448 = v_2544 | ~v_1084;
assign x_20449 = v_2544 | ~v_2496;
assign x_20450 = v_2544 | ~v_2497;
assign x_20451 = v_2544 | ~v_2498;
assign x_20452 = v_2544 | ~v_2499;
assign x_20453 = v_2544 | ~v_1085;
assign x_20454 = v_2544 | ~v_1086;
assign x_20455 = v_2544 | ~v_2532;
assign x_20456 = v_2544 | ~v_2533;
assign x_20457 = v_2544 | ~v_2534;
assign x_20458 = v_2544 | ~v_2535;
assign x_20459 = v_2544 | ~v_2446;
assign x_20460 = v_2544 | ~v_2449;
assign x_20461 = v_2544 | ~v_184;
assign x_20462 = v_2544 | ~v_171;
assign x_20463 = v_2544 | ~v_169;
assign x_20464 = v_2544 | ~v_160;
assign x_20465 = v_2544 | ~v_150;
assign x_20466 = v_2544 | ~v_149;
assign x_20467 = v_2544 | ~v_147;
assign x_20468 = v_2544 | ~v_103;
assign x_20469 = v_2544 | ~v_102;
assign x_20470 = v_2544 | ~v_100;
assign x_20471 = v_2544 | ~v_96;
assign x_20472 = v_2544 | ~v_94;
assign x_20473 = v_2543 | ~v_2423;
assign x_20474 = v_2543 | ~v_2424;
assign x_20475 = v_2543 | ~v_2425;
assign x_20476 = v_2543 | ~v_2426;
assign x_20477 = v_2543 | ~v_1769;
assign x_20478 = v_2543 | ~v_1770;
assign x_20479 = v_2543 | ~v_1771;
assign x_20480 = v_2543 | ~v_1772;
assign x_20481 = v_2543 | ~v_1709;
assign x_20482 = v_2543 | ~v_1710;
assign x_20483 = v_2543 | ~v_1711;
assign x_20484 = v_2543 | ~v_1712;
assign x_20485 = v_2543 | ~v_1601;
assign x_20486 = v_2543 | ~v_1604;
assign x_20487 = v_2543 | ~v_804;
assign x_20488 = v_2543 | ~v_805;
assign x_20489 = v_2543 | ~v_1066;
assign x_20490 = v_2543 | ~v_1067;
assign x_20491 = v_2543 | ~v_1068;
assign x_20492 = v_2543 | ~v_1069;
assign x_20493 = v_2543 | ~v_2491;
assign x_20494 = v_2543 | ~v_2492;
assign x_20495 = v_2543 | ~v_2493;
assign x_20496 = v_2543 | ~v_2494;
assign x_20497 = v_2543 | ~v_1070;
assign x_20498 = v_2543 | ~v_1071;
assign x_20499 = v_2543 | ~v_2527;
assign x_20500 = v_2543 | ~v_2528;
assign x_20501 = v_2543 | ~v_2529;
assign x_20502 = v_2543 | ~v_2530;
assign x_20503 = v_2543 | ~v_2431;
assign x_20504 = v_2543 | ~v_2434;
assign x_20505 = v_2543 | ~v_183;
assign x_20506 = v_2543 | ~v_167;
assign x_20507 = v_2543 | ~v_165;
assign x_20508 = v_2543 | ~v_159;
assign x_20509 = v_2543 | ~v_145;
assign x_20510 = v_2543 | ~v_144;
assign x_20511 = v_2543 | ~v_142;
assign x_20512 = v_2543 | ~v_61;
assign x_20513 = v_2543 | ~v_60;
assign x_20514 = v_2543 | ~v_58;
assign x_20515 = v_2543 | ~v_54;
assign x_20516 = v_2543 | ~v_52;
assign x_20517 = v_2542 | ~v_2408;
assign x_20518 = v_2542 | ~v_2409;
assign x_20519 = v_2542 | ~v_2410;
assign x_20520 = v_2542 | ~v_2411;
assign x_20521 = v_2542 | ~v_1760;
assign x_20522 = v_2542 | ~v_1761;
assign x_20523 = v_2542 | ~v_1762;
assign x_20524 = v_2542 | ~v_1763;
assign x_20525 = v_2542 | ~v_1700;
assign x_20526 = v_2542 | ~v_1701;
assign x_20527 = v_2542 | ~v_1702;
assign x_20528 = v_2542 | ~v_1703;
assign x_20529 = v_2542 | ~v_1576;
assign x_20530 = v_2542 | ~v_1579;
assign x_20531 = v_2542 | ~v_771;
assign x_20532 = v_2542 | ~v_772;
assign x_20533 = v_2542 | ~v_1051;
assign x_20534 = v_2542 | ~v_1052;
assign x_20535 = v_2542 | ~v_1053;
assign x_20536 = v_2542 | ~v_1054;
assign x_20537 = v_2542 | ~v_2486;
assign x_20538 = v_2542 | ~v_2487;
assign x_20539 = v_2542 | ~v_2488;
assign x_20540 = v_2542 | ~v_2489;
assign x_20541 = v_2542 | ~v_1055;
assign x_20542 = v_2542 | ~v_1056;
assign x_20543 = v_2542 | ~v_2522;
assign x_20544 = v_2542 | ~v_2523;
assign x_20545 = v_2542 | ~v_2524;
assign x_20546 = v_2542 | ~v_2525;
assign x_20547 = v_2542 | ~v_2416;
assign x_20548 = v_2542 | ~v_2419;
assign x_20549 = v_2542 | ~v_182;
assign x_20550 = v_2542 | ~v_163;
assign x_20551 = v_2542 | ~v_161;
assign x_20552 = v_2542 | ~v_155;
assign x_20553 = v_2542 | ~v_137;
assign x_20554 = v_2542 | ~v_136;
assign x_20555 = v_2542 | ~v_134;
assign x_20556 = v_2542 | ~v_18;
assign x_20557 = v_2542 | ~v_17;
assign x_20558 = v_2542 | ~v_15;
assign x_20559 = v_2542 | ~v_11;
assign x_20560 = v_2542 | ~v_9;
assign x_20561 = ~v_2540 | ~v_2539 | ~v_2538 | v_2541;
assign x_20562 = v_2540 | ~v_2438;
assign x_20563 = v_2540 | ~v_2439;
assign x_20564 = v_2540 | ~v_2440;
assign x_20565 = v_2540 | ~v_2441;
assign x_20566 = v_2540 | ~v_1778;
assign x_20567 = v_2540 | ~v_1779;
assign x_20568 = v_2540 | ~v_1780;
assign x_20569 = v_2540 | ~v_1781;
assign x_20570 = v_2540 | ~v_1690;
assign x_20571 = v_2540 | ~v_1691;
assign x_20572 = v_2540 | ~v_1692;
assign x_20573 = v_2540 | ~v_1693;
assign x_20574 = v_2540 | ~v_1626;
assign x_20575 = v_2540 | ~v_1629;
assign x_20576 = v_2540 | ~v_927;
assign x_20577 = v_2540 | ~v_928;
assign x_20578 = v_2540 | ~v_1099;
assign x_20579 = v_2540 | ~v_1100;
assign x_20580 = v_2540 | ~v_1101;
assign x_20581 = v_2540 | ~v_1102;
assign x_20582 = v_2540 | ~v_2480;
assign x_20583 = v_2540 | ~v_2481;
assign x_20584 = v_2540 | ~v_2482;
assign x_20585 = v_2540 | ~v_2483;
assign x_20586 = v_2540 | ~v_1085;
assign x_20587 = v_2540 | ~v_1086;
assign x_20588 = v_2540 | ~v_2532;
assign x_20589 = v_2540 | ~v_2533;
assign x_20590 = v_2540 | ~v_2534;
assign x_20591 = v_2540 | ~v_2535;
assign x_20592 = v_2540 | ~v_2446;
assign x_20593 = v_2540 | ~v_2449;
assign x_20594 = v_2540 | ~v_184;
assign x_20595 = v_2540 | ~v_171;
assign x_20596 = v_2540 | ~v_169;
assign x_20597 = v_2540 | ~v_150;
assign x_20598 = v_2540 | ~v_148;
assign x_20599 = v_2540 | ~v_103;
assign x_20600 = v_2540 | ~v_102;
assign x_20601 = v_2540 | ~v_101;
assign x_20602 = v_2540 | ~v_100;
assign x_20603 = v_2540 | ~v_97;
assign x_20604 = v_2540 | ~v_95;
assign x_20605 = v_2540 | ~v_94;
assign x_20606 = v_2539 | ~v_2423;
assign x_20607 = v_2539 | ~v_2424;
assign x_20608 = v_2539 | ~v_2425;
assign x_20609 = v_2539 | ~v_2426;
assign x_20610 = v_2539 | ~v_1769;
assign x_20611 = v_2539 | ~v_1770;
assign x_20612 = v_2539 | ~v_1771;
assign x_20613 = v_2539 | ~v_1772;
assign x_20614 = v_2539 | ~v_1681;
assign x_20615 = v_2539 | ~v_1682;
assign x_20616 = v_2539 | ~v_1683;
assign x_20617 = v_2539 | ~v_1684;
assign x_20618 = v_2539 | ~v_1601;
assign x_20619 = v_2539 | ~v_1604;
assign x_20620 = v_2539 | ~v_912;
assign x_20621 = v_2539 | ~v_913;
assign x_20622 = v_2539 | ~v_1094;
assign x_20623 = v_2539 | ~v_1095;
assign x_20624 = v_2539 | ~v_1096;
assign x_20625 = v_2539 | ~v_1097;
assign x_20626 = v_2539 | ~v_2475;
assign x_20627 = v_2539 | ~v_2476;
assign x_20628 = v_2539 | ~v_2477;
assign x_20629 = v_2539 | ~v_2478;
assign x_20630 = v_2539 | ~v_1070;
assign x_20631 = v_2539 | ~v_1071;
assign x_20632 = v_2539 | ~v_2527;
assign x_20633 = v_2539 | ~v_2528;
assign x_20634 = v_2539 | ~v_2529;
assign x_20635 = v_2539 | ~v_2530;
assign x_20636 = v_2539 | ~v_2431;
assign x_20637 = v_2539 | ~v_2434;
assign x_20638 = v_2539 | ~v_183;
assign x_20639 = v_2539 | ~v_167;
assign x_20640 = v_2539 | ~v_165;
assign x_20641 = v_2539 | ~v_145;
assign x_20642 = v_2539 | ~v_143;
assign x_20643 = v_2539 | ~v_61;
assign x_20644 = v_2539 | ~v_60;
assign x_20645 = v_2539 | ~v_59;
assign x_20646 = v_2539 | ~v_58;
assign x_20647 = v_2539 | ~v_55;
assign x_20648 = v_2539 | ~v_53;
assign x_20649 = v_2539 | ~v_52;
assign x_20650 = v_2538 | ~v_2408;
assign x_20651 = v_2538 | ~v_2409;
assign x_20652 = v_2538 | ~v_2410;
assign x_20653 = v_2538 | ~v_2411;
assign x_20654 = v_2538 | ~v_1760;
assign x_20655 = v_2538 | ~v_1761;
assign x_20656 = v_2538 | ~v_1762;
assign x_20657 = v_2538 | ~v_1763;
assign x_20658 = v_2538 | ~v_1672;
assign x_20659 = v_2538 | ~v_1673;
assign x_20660 = v_2538 | ~v_1674;
assign x_20661 = v_2538 | ~v_1675;
assign x_20662 = v_2538 | ~v_1576;
assign x_20663 = v_2538 | ~v_1579;
assign x_20664 = v_2538 | ~v_897;
assign x_20665 = v_2538 | ~v_898;
assign x_20666 = v_2538 | ~v_1089;
assign x_20667 = v_2538 | ~v_1090;
assign x_20668 = v_2538 | ~v_1091;
assign x_20669 = v_2538 | ~v_1092;
assign x_20670 = v_2538 | ~v_2470;
assign x_20671 = v_2538 | ~v_2471;
assign x_20672 = v_2538 | ~v_2472;
assign x_20673 = v_2538 | ~v_2473;
assign x_20674 = v_2538 | ~v_1055;
assign x_20675 = v_2538 | ~v_1056;
assign x_20676 = v_2538 | ~v_2522;
assign x_20677 = v_2538 | ~v_2523;
assign x_20678 = v_2538 | ~v_2524;
assign x_20679 = v_2538 | ~v_2525;
assign x_20680 = v_2538 | ~v_2416;
assign x_20681 = v_2538 | ~v_2419;
assign x_20682 = v_2538 | ~v_182;
assign x_20683 = v_2538 | ~v_163;
assign x_20684 = v_2538 | ~v_161;
assign x_20685 = v_2538 | ~v_137;
assign x_20686 = v_2538 | ~v_135;
assign x_20687 = v_2538 | ~v_18;
assign x_20688 = v_2538 | ~v_17;
assign x_20689 = v_2538 | ~v_16;
assign x_20690 = v_2538 | ~v_15;
assign x_20691 = v_2538 | ~v_12;
assign x_20692 = v_2538 | ~v_10;
assign x_20693 = v_2538 | ~v_9;
assign x_20694 = ~v_2536 | ~v_2531 | ~v_2526 | v_2537;
assign x_20695 = v_2536 | ~v_2438;
assign x_20696 = v_2536 | ~v_2439;
assign x_20697 = v_2536 | ~v_2440;
assign x_20698 = v_2536 | ~v_2441;
assign x_20699 = v_2536 | ~v_1778;
assign x_20700 = v_2536 | ~v_1779;
assign x_20701 = v_2536 | ~v_1780;
assign x_20702 = v_2536 | ~v_1781;
assign x_20703 = v_2536 | ~v_1622;
assign x_20704 = v_2536 | ~v_1623;
assign x_20705 = v_2536 | ~v_1624;
assign x_20706 = v_2536 | ~v_1625;
assign x_20707 = v_2536 | ~v_1626;
assign x_20708 = v_2536 | ~v_1629;
assign x_20709 = v_2536 | ~v_975;
assign x_20710 = v_2536 | ~v_976;
assign x_20711 = v_2536 | ~v_1115;
assign x_20712 = v_2536 | ~v_1116;
assign x_20713 = v_2536 | ~v_2442;
assign x_20714 = v_2536 | ~v_2443;
assign x_20715 = v_2536 | ~v_2444;
assign x_20716 = v_2536 | ~v_2445;
assign x_20717 = v_2536 | ~v_1085;
assign x_20718 = v_2536 | ~v_1086;
assign x_20719 = v_2536 | ~v_2532;
assign x_20720 = v_2536 | ~v_2533;
assign x_20721 = v_2536 | ~v_2534;
assign x_20722 = v_2536 | ~v_2535;
assign x_20723 = v_2536 | ~v_2446;
assign x_20724 = v_2536 | ~v_2449;
assign x_20725 = v_2536 | ~v_1117;
assign x_20726 = v_2536 | ~v_1118;
assign x_20727 = v_2536 | ~v_184;
assign x_20728 = v_2536 | ~v_171;
assign x_20729 = v_2536 | ~v_169;
assign x_20730 = v_2536 | ~v_151;
assign x_20731 = v_2536 | ~v_150;
assign x_20732 = v_2536 | ~v_149;
assign x_20733 = v_2536 | ~v_148;
assign x_20734 = v_2536 | ~v_147;
assign x_20735 = v_2536 | ~v_103;
assign x_20736 = v_2536 | ~v_101;
assign x_20737 = v_2536 | ~v_100;
assign x_20738 = v_2536 | ~v_94;
assign x_20739 = ~v_128 | ~v_141 | v_2535;
assign x_20740 = ~v_125 | ~v_141 | v_2534;
assign x_20741 = ~v_113 | v_141 | v_2533;
assign x_20742 = ~v_110 | v_141 | v_2532;
assign x_20743 = v_2531 | ~v_2423;
assign x_20744 = v_2531 | ~v_2424;
assign x_20745 = v_2531 | ~v_2425;
assign x_20746 = v_2531 | ~v_2426;
assign x_20747 = v_2531 | ~v_1769;
assign x_20748 = v_2531 | ~v_1770;
assign x_20749 = v_2531 | ~v_1771;
assign x_20750 = v_2531 | ~v_1772;
assign x_20751 = v_2531 | ~v_1597;
assign x_20752 = v_2531 | ~v_1598;
assign x_20753 = v_2531 | ~v_1599;
assign x_20754 = v_2531 | ~v_1600;
assign x_20755 = v_2531 | ~v_1601;
assign x_20756 = v_2531 | ~v_1604;
assign x_20757 = v_2531 | ~v_960;
assign x_20758 = v_2531 | ~v_961;
assign x_20759 = v_2531 | ~v_1110;
assign x_20760 = v_2531 | ~v_1111;
assign x_20761 = v_2531 | ~v_2427;
assign x_20762 = v_2531 | ~v_2428;
assign x_20763 = v_2531 | ~v_2429;
assign x_20764 = v_2531 | ~v_2430;
assign x_20765 = v_2531 | ~v_1070;
assign x_20766 = v_2531 | ~v_1071;
assign x_20767 = v_2531 | ~v_2527;
assign x_20768 = v_2531 | ~v_2528;
assign x_20769 = v_2531 | ~v_2529;
assign x_20770 = v_2531 | ~v_2530;
assign x_20771 = v_2531 | ~v_2431;
assign x_20772 = v_2531 | ~v_2434;
assign x_20773 = v_2531 | ~v_1112;
assign x_20774 = v_2531 | ~v_1113;
assign x_20775 = v_2531 | ~v_183;
assign x_20776 = v_2531 | ~v_167;
assign x_20777 = v_2531 | ~v_165;
assign x_20778 = v_2531 | ~v_146;
assign x_20779 = v_2531 | ~v_145;
assign x_20780 = v_2531 | ~v_144;
assign x_20781 = v_2531 | ~v_143;
assign x_20782 = v_2531 | ~v_142;
assign x_20783 = v_2531 | ~v_61;
assign x_20784 = v_2531 | ~v_59;
assign x_20785 = v_2531 | ~v_58;
assign x_20786 = v_2531 | ~v_52;
assign x_20787 = ~v_86 | ~v_141 | v_2530;
assign x_20788 = ~v_83 | ~v_141 | v_2529;
assign x_20789 = ~v_71 | v_141 | v_2528;
assign x_20790 = ~v_68 | v_141 | v_2527;
assign x_20791 = v_2526 | ~v_2408;
assign x_20792 = v_2526 | ~v_2409;
assign x_20793 = v_2526 | ~v_2410;
assign x_20794 = v_2526 | ~v_2411;
assign x_20795 = v_2526 | ~v_1760;
assign x_20796 = v_2526 | ~v_1761;
assign x_20797 = v_2526 | ~v_1762;
assign x_20798 = v_2526 | ~v_1763;
assign x_20799 = v_2526 | ~v_1572;
assign x_20800 = v_2526 | ~v_1573;
assign x_20801 = v_2526 | ~v_1574;
assign x_20802 = v_2526 | ~v_1575;
assign x_20803 = v_2526 | ~v_1576;
assign x_20804 = v_2526 | ~v_1579;
assign x_20805 = v_2526 | ~v_945;
assign x_20806 = v_2526 | ~v_946;
assign x_20807 = v_2526 | ~v_1105;
assign x_20808 = v_2526 | ~v_1106;
assign x_20809 = v_2526 | ~v_2412;
assign x_20810 = v_2526 | ~v_2413;
assign x_20811 = v_2526 | ~v_2414;
assign x_20812 = v_2526 | ~v_2415;
assign x_20813 = v_2526 | ~v_1055;
assign x_20814 = v_2526 | ~v_1056;
assign x_20815 = v_2526 | ~v_2522;
assign x_20816 = v_2526 | ~v_2523;
assign x_20817 = v_2526 | ~v_2524;
assign x_20818 = v_2526 | ~v_2525;
assign x_20819 = v_2526 | ~v_2416;
assign x_20820 = v_2526 | ~v_2419;
assign x_20821 = v_2526 | ~v_1107;
assign x_20822 = v_2526 | ~v_1108;
assign x_20823 = v_2526 | ~v_182;
assign x_20824 = v_2526 | ~v_163;
assign x_20825 = v_2526 | ~v_161;
assign x_20826 = v_2526 | ~v_138;
assign x_20827 = v_2526 | ~v_137;
assign x_20828 = v_2526 | ~v_136;
assign x_20829 = v_2526 | ~v_135;
assign x_20830 = v_2526 | ~v_134;
assign x_20831 = v_2526 | ~v_18;
assign x_20832 = v_2526 | ~v_16;
assign x_20833 = v_2526 | ~v_15;
assign x_20834 = v_2526 | ~v_9;
assign x_20835 = ~v_44 | ~v_141 | v_2525;
assign x_20836 = ~v_41 | ~v_141 | v_2524;
assign x_20837 = ~v_29 | v_141 | v_2523;
assign x_20838 = ~v_26 | v_141 | v_2522;
assign x_20839 = ~v_2520 | ~v_2519 | ~v_2518 | v_2521;
assign x_20840 = v_2520 | ~v_2438;
assign x_20841 = v_2520 | ~v_2439;
assign x_20842 = v_2520 | ~v_2440;
assign x_20843 = v_2520 | ~v_2441;
assign x_20844 = v_2520 | ~v_1690;
assign x_20845 = v_2520 | ~v_1691;
assign x_20846 = v_2520 | ~v_1692;
assign x_20847 = v_2520 | ~v_1693;
assign x_20848 = v_2520 | ~v_1626;
assign x_20849 = v_2520 | ~v_1627;
assign x_20850 = v_2520 | ~v_1628;
assign x_20851 = v_2520 | ~v_1629;
assign x_20852 = v_2520 | ~v_1630;
assign x_20853 = v_2520 | ~v_1631;
assign x_20854 = v_2520 | ~v_1037;
assign x_20855 = v_2520 | ~v_1038;
assign x_20856 = v_2520 | ~v_1039;
assign x_20857 = v_2520 | ~v_1040;
assign x_20858 = v_2520 | ~v_927;
assign x_20859 = v_2520 | ~v_928;
assign x_20860 = v_2520 | ~v_2480;
assign x_20861 = v_2520 | ~v_2481;
assign x_20862 = v_2520 | ~v_2482;
assign x_20863 = v_2520 | ~v_2483;
assign x_20864 = v_2520 | ~v_839;
assign x_20865 = v_2520 | ~v_840;
assign x_20866 = v_2520 | ~v_2446;
assign x_20867 = v_2520 | ~v_2447;
assign x_20868 = v_2520 | ~v_2448;
assign x_20869 = v_2520 | ~v_2449;
assign x_20870 = v_2520 | ~v_2450;
assign x_20871 = v_2520 | ~v_2451;
assign x_20872 = v_2520 | ~v_184;
assign x_20873 = v_2520 | ~v_170;
assign x_20874 = v_2520 | ~v_169;
assign x_20875 = v_2520 | ~v_151;
assign x_20876 = v_2520 | ~v_150;
assign x_20877 = v_2520 | ~v_148;
assign x_20878 = v_2520 | ~v_147;
assign x_20879 = v_2520 | ~v_103;
assign x_20880 = v_2520 | ~v_101;
assign x_20881 = v_2520 | ~v_100;
assign x_20882 = v_2520 | ~v_98;
assign x_20883 = v_2520 | ~v_97;
assign x_20884 = v_2519 | ~v_2423;
assign x_20885 = v_2519 | ~v_2424;
assign x_20886 = v_2519 | ~v_2425;
assign x_20887 = v_2519 | ~v_2426;
assign x_20888 = v_2519 | ~v_1681;
assign x_20889 = v_2519 | ~v_1682;
assign x_20890 = v_2519 | ~v_1683;
assign x_20891 = v_2519 | ~v_1684;
assign x_20892 = v_2519 | ~v_1601;
assign x_20893 = v_2519 | ~v_1602;
assign x_20894 = v_2519 | ~v_1603;
assign x_20895 = v_2519 | ~v_1604;
assign x_20896 = v_2519 | ~v_1605;
assign x_20897 = v_2519 | ~v_1606;
assign x_20898 = v_2519 | ~v_1032;
assign x_20899 = v_2519 | ~v_1033;
assign x_20900 = v_2519 | ~v_1034;
assign x_20901 = v_2519 | ~v_1035;
assign x_20902 = v_2519 | ~v_912;
assign x_20903 = v_2519 | ~v_913;
assign x_20904 = v_2519 | ~v_2475;
assign x_20905 = v_2519 | ~v_2476;
assign x_20906 = v_2519 | ~v_2477;
assign x_20907 = v_2519 | ~v_2478;
assign x_20908 = v_2519 | ~v_806;
assign x_20909 = v_2519 | ~v_2431;
assign x_20910 = v_2519 | ~v_2432;
assign x_20911 = v_2519 | ~v_2433;
assign x_20912 = v_2519 | ~v_2434;
assign x_20913 = v_2519 | ~v_2435;
assign x_20914 = v_2519 | ~v_2436;
assign x_20915 = v_2519 | ~v_807;
assign x_20916 = v_2519 | ~v_183;
assign x_20917 = v_2519 | ~v_166;
assign x_20918 = v_2519 | ~v_165;
assign x_20919 = v_2519 | ~v_146;
assign x_20920 = v_2519 | ~v_145;
assign x_20921 = v_2519 | ~v_143;
assign x_20922 = v_2519 | ~v_142;
assign x_20923 = v_2519 | ~v_61;
assign x_20924 = v_2519 | ~v_59;
assign x_20925 = v_2519 | ~v_58;
assign x_20926 = v_2519 | ~v_56;
assign x_20927 = v_2519 | ~v_55;
assign x_20928 = v_2518 | ~v_2408;
assign x_20929 = v_2518 | ~v_2409;
assign x_20930 = v_2518 | ~v_2410;
assign x_20931 = v_2518 | ~v_2411;
assign x_20932 = v_2518 | ~v_1672;
assign x_20933 = v_2518 | ~v_1673;
assign x_20934 = v_2518 | ~v_1674;
assign x_20935 = v_2518 | ~v_1675;
assign x_20936 = v_2518 | ~v_1576;
assign x_20937 = v_2518 | ~v_1577;
assign x_20938 = v_2518 | ~v_1578;
assign x_20939 = v_2518 | ~v_1579;
assign x_20940 = v_2518 | ~v_1580;
assign x_20941 = v_2518 | ~v_1581;
assign x_20942 = v_2518 | ~v_1027;
assign x_20943 = v_2518 | ~v_1028;
assign x_20944 = v_2518 | ~v_1029;
assign x_20945 = v_2518 | ~v_1030;
assign x_20946 = v_2518 | ~v_897;
assign x_20947 = v_2518 | ~v_898;
assign x_20948 = v_2518 | ~v_2470;
assign x_20949 = v_2518 | ~v_2471;
assign x_20950 = v_2518 | ~v_2472;
assign x_20951 = v_2518 | ~v_2473;
assign x_20952 = v_2518 | ~v_773;
assign x_20953 = v_2518 | ~v_774;
assign x_20954 = v_2518 | ~v_2416;
assign x_20955 = v_2518 | ~v_2417;
assign x_20956 = v_2518 | ~v_2418;
assign x_20957 = v_2518 | ~v_2419;
assign x_20958 = v_2518 | ~v_2420;
assign x_20959 = v_2518 | ~v_2421;
assign x_20960 = v_2518 | ~v_182;
assign x_20961 = v_2518 | ~v_162;
assign x_20962 = v_2518 | ~v_161;
assign x_20963 = v_2518 | ~v_138;
assign x_20964 = v_2518 | ~v_137;
assign x_20965 = v_2518 | ~v_135;
assign x_20966 = v_2518 | ~v_134;
assign x_20967 = v_2518 | ~v_18;
assign x_20968 = v_2518 | ~v_16;
assign x_20969 = v_2518 | ~v_15;
assign x_20970 = v_2518 | ~v_13;
assign x_20971 = v_2518 | ~v_12;
assign x_20972 = ~v_2516 | ~v_2511 | ~v_2506 | v_2517;
assign x_20973 = v_2516 | ~v_2438;
assign x_20974 = v_2516 | ~v_2439;
assign x_20975 = v_2516 | ~v_2440;
assign x_20976 = v_2516 | ~v_2441;
assign x_20977 = v_2516 | ~v_1662;
assign x_20978 = v_2516 | ~v_1663;
assign x_20979 = v_2516 | ~v_1664;
assign x_20980 = v_2516 | ~v_1665;
assign x_20981 = v_2516 | ~v_1626;
assign x_20982 = v_2516 | ~v_1746;
assign x_20983 = v_2516 | ~v_1747;
assign x_20984 = v_2516 | ~v_1629;
assign x_20985 = v_2516 | ~v_1748;
assign x_20986 = v_2516 | ~v_1749;
assign x_20987 = v_2516 | ~v_1193;
assign x_20988 = v_2516 | ~v_1241;
assign x_20989 = v_2516 | ~v_1194;
assign x_20990 = v_2516 | ~v_1242;
assign x_20991 = v_2516 | ~v_2464;
assign x_20992 = v_2516 | ~v_2465;
assign x_20993 = v_2516 | ~v_2466;
assign x_20994 = v_2516 | ~v_2467;
assign x_20995 = v_2516 | ~v_1023;
assign x_20996 = v_2516 | ~v_1024;
assign x_20997 = v_2516 | ~v_2446;
assign x_20998 = v_2516 | ~v_2512;
assign x_20999 = v_2516 | ~v_2513;
assign x_21000 = v_2516 | ~v_2449;
assign x_21001 = v_2516 | ~v_2514;
assign x_21002 = v_2516 | ~v_2515;
assign x_21003 = v_2516 | ~v_1243;
assign x_21004 = v_2516 | ~v_1244;
assign x_21005 = v_2516 | ~v_184;
assign x_21006 = v_2516 | ~v_171;
assign x_21007 = v_2516 | ~v_170;
assign x_21008 = v_2516 | ~v_169;
assign x_21009 = v_2516 | ~v_149;
assign x_21010 = v_2516 | ~v_148;
assign x_21011 = v_2516 | ~v_147;
assign x_21012 = v_2516 | ~v_103;
assign x_21013 = v_2516 | ~v_102;
assign x_21014 = v_2516 | ~v_101;
assign x_21015 = v_2516 | ~v_100;
assign x_21016 = v_2516 | ~v_99;
assign x_21017 = ~v_131 | ~v_139 | v_2515;
assign x_21018 = ~v_126 | ~v_140 | v_2514;
assign x_21019 = ~v_116 | v_139 | v_2513;
assign x_21020 = ~v_111 | v_140 | v_2512;
assign x_21021 = v_2511 | ~v_2423;
assign x_21022 = v_2511 | ~v_2424;
assign x_21023 = v_2511 | ~v_2425;
assign x_21024 = v_2511 | ~v_2426;
assign x_21025 = v_2511 | ~v_1653;
assign x_21026 = v_2511 | ~v_1654;
assign x_21027 = v_2511 | ~v_1655;
assign x_21028 = v_2511 | ~v_1656;
assign x_21029 = v_2511 | ~v_1601;
assign x_21030 = v_2511 | ~v_1737;
assign x_21031 = v_2511 | ~v_1738;
assign x_21032 = v_2511 | ~v_1604;
assign x_21033 = v_2511 | ~v_1739;
assign x_21034 = v_2511 | ~v_1740;
assign x_21035 = v_2511 | ~v_1178;
assign x_21036 = v_2511 | ~v_1236;
assign x_21037 = v_2511 | ~v_1179;
assign x_21038 = v_2511 | ~v_1237;
assign x_21039 = v_2511 | ~v_2459;
assign x_21040 = v_2511 | ~v_2460;
assign x_21041 = v_2511 | ~v_2461;
assign x_21042 = v_2511 | ~v_2462;
assign x_21043 = v_2511 | ~v_1008;
assign x_21044 = v_2511 | ~v_1009;
assign x_21045 = v_2511 | ~v_2431;
assign x_21046 = v_2511 | ~v_2507;
assign x_21047 = v_2511 | ~v_2508;
assign x_21048 = v_2511 | ~v_2434;
assign x_21049 = v_2511 | ~v_2509;
assign x_21050 = v_2511 | ~v_2510;
assign x_21051 = v_2511 | ~v_1238;
assign x_21052 = v_2511 | ~v_1239;
assign x_21053 = v_2511 | ~v_183;
assign x_21054 = v_2511 | ~v_167;
assign x_21055 = v_2511 | ~v_166;
assign x_21056 = v_2511 | ~v_165;
assign x_21057 = v_2511 | ~v_144;
assign x_21058 = v_2511 | ~v_143;
assign x_21059 = v_2511 | ~v_142;
assign x_21060 = v_2511 | ~v_61;
assign x_21061 = v_2511 | ~v_60;
assign x_21062 = v_2511 | ~v_59;
assign x_21063 = v_2511 | ~v_58;
assign x_21064 = v_2511 | ~v_57;
assign x_21065 = ~v_89 | ~v_139 | v_2510;
assign x_21066 = ~v_84 | ~v_140 | v_2509;
assign x_21067 = ~v_74 | v_139 | v_2508;
assign x_21068 = ~v_69 | v_140 | v_2507;
assign x_21069 = v_2506 | ~v_2408;
assign x_21070 = v_2506 | ~v_2409;
assign x_21071 = v_2506 | ~v_2410;
assign x_21072 = v_2506 | ~v_2411;
assign x_21073 = v_2506 | ~v_1644;
assign x_21074 = v_2506 | ~v_1645;
assign x_21075 = v_2506 | ~v_1646;
assign x_21076 = v_2506 | ~v_1647;
assign x_21077 = v_2506 | ~v_1576;
assign x_21078 = v_2506 | ~v_1728;
assign x_21079 = v_2506 | ~v_1729;
assign x_21080 = v_2506 | ~v_1579;
assign x_21081 = v_2506 | ~v_1730;
assign x_21082 = v_2506 | ~v_1731;
assign x_21083 = v_2506 | ~v_1163;
assign x_21084 = v_2506 | ~v_1231;
assign x_21085 = v_2506 | ~v_1164;
assign x_21086 = v_2506 | ~v_1232;
assign x_21087 = v_2506 | ~v_2454;
assign x_21088 = v_2506 | ~v_2455;
assign x_21089 = v_2506 | ~v_2456;
assign x_21090 = v_2506 | ~v_2457;
assign x_21091 = v_2506 | ~v_2416;
assign x_21092 = v_2506 | ~v_2502;
assign x_21093 = v_2506 | ~v_2503;
assign x_21094 = v_2506 | ~v_2419;
assign x_21095 = v_2506 | ~v_2504;
assign x_21096 = v_2506 | ~v_2505;
assign x_21097 = v_2506 | ~v_1233;
assign x_21098 = v_2506 | ~v_1234;
assign x_21099 = v_2506 | ~v_182;
assign x_21100 = v_2506 | ~v_163;
assign x_21101 = v_2506 | ~v_162;
assign x_21102 = v_2506 | ~v_161;
assign x_21103 = v_2506 | ~v_136;
assign x_21104 = v_2506 | ~v_135;
assign x_21105 = v_2506 | ~v_134;
assign x_21106 = v_2506 | ~v_993;
assign x_21107 = v_2506 | ~v_994;
assign x_21108 = v_2506 | ~v_18;
assign x_21109 = v_2506 | ~v_17;
assign x_21110 = v_2506 | ~v_16;
assign x_21111 = v_2506 | ~v_15;
assign x_21112 = v_2506 | ~v_14;
assign x_21113 = ~v_47 | ~v_139 | v_2505;
assign x_21114 = ~v_42 | ~v_140 | v_2504;
assign x_21115 = ~v_32 | v_139 | v_2503;
assign x_21116 = ~v_27 | v_140 | v_2502;
assign x_21117 = ~v_2500 | ~v_2495 | ~v_2490 | v_2501;
assign x_21118 = v_2500 | ~v_2438;
assign x_21119 = v_2500 | ~v_2439;
assign x_21120 = v_2500 | ~v_2440;
assign x_21121 = v_2500 | ~v_2441;
assign x_21122 = v_2500 | ~v_1662;
assign x_21123 = v_2500 | ~v_1663;
assign x_21124 = v_2500 | ~v_1664;
assign x_21125 = v_2500 | ~v_1665;
assign x_21126 = v_2500 | ~v_1718;
assign x_21127 = v_2500 | ~v_1719;
assign x_21128 = v_2500 | ~v_1720;
assign x_21129 = v_2500 | ~v_1721;
assign x_21130 = v_2500 | ~v_1626;
assign x_21131 = v_2500 | ~v_1629;
assign x_21132 = v_2500 | ~v_1191;
assign x_21133 = v_2500 | ~v_1192;
assign x_21134 = v_2500 | ~v_1193;
assign x_21135 = v_2500 | ~v_1194;
assign x_21136 = v_2500 | ~v_2464;
assign x_21137 = v_2500 | ~v_2465;
assign x_21138 = v_2500 | ~v_2466;
assign x_21139 = v_2500 | ~v_2467;
assign x_21140 = v_2500 | ~v_837;
assign x_21141 = v_2500 | ~v_838;
assign x_21142 = v_2500 | ~v_2496;
assign x_21143 = v_2500 | ~v_2497;
assign x_21144 = v_2500 | ~v_2498;
assign x_21145 = v_2500 | ~v_2499;
assign x_21146 = v_2500 | ~v_2446;
assign x_21147 = v_2500 | ~v_2449;
assign x_21148 = v_2500 | ~v_1195;
assign x_21149 = v_2500 | ~v_1196;
assign x_21150 = v_2500 | ~v_184;
assign x_21151 = v_2500 | ~v_171;
assign x_21152 = v_2500 | ~v_170;
assign x_21153 = v_2500 | ~v_169;
assign x_21154 = v_2500 | ~v_160;
assign x_21155 = v_2500 | ~v_151;
assign x_21156 = v_2500 | ~v_150;
assign x_21157 = v_2500 | ~v_149;
assign x_21158 = v_2500 | ~v_147;
assign x_21159 = v_2500 | ~v_103;
assign x_21160 = v_2500 | ~v_100;
assign x_21161 = v_2500 | ~v_96;
assign x_21162 = ~v_131 | ~v_176 | v_2499;
assign x_21163 = ~v_126 | ~v_175 | v_2498;
assign x_21164 = ~v_116 | v_176 | v_2497;
assign x_21165 = ~v_111 | v_175 | v_2496;
assign x_21166 = v_2495 | ~v_2423;
assign x_21167 = v_2495 | ~v_2424;
assign x_21168 = v_2495 | ~v_2425;
assign x_21169 = v_2495 | ~v_2426;
assign x_21170 = v_2495 | ~v_1653;
assign x_21171 = v_2495 | ~v_1654;
assign x_21172 = v_2495 | ~v_1655;
assign x_21173 = v_2495 | ~v_1656;
assign x_21174 = v_2495 | ~v_1709;
assign x_21175 = v_2495 | ~v_1710;
assign x_21176 = v_2495 | ~v_1711;
assign x_21177 = v_2495 | ~v_1712;
assign x_21178 = v_2495 | ~v_1601;
assign x_21179 = v_2495 | ~v_1604;
assign x_21180 = v_2495 | ~v_1176;
assign x_21181 = v_2495 | ~v_1177;
assign x_21182 = v_2495 | ~v_1178;
assign x_21183 = v_2495 | ~v_1179;
assign x_21184 = v_2495 | ~v_2459;
assign x_21185 = v_2495 | ~v_2460;
assign x_21186 = v_2495 | ~v_2461;
assign x_21187 = v_2495 | ~v_2462;
assign x_21188 = v_2495 | ~v_804;
assign x_21189 = v_2495 | ~v_805;
assign x_21190 = v_2495 | ~v_2491;
assign x_21191 = v_2495 | ~v_2492;
assign x_21192 = v_2495 | ~v_2493;
assign x_21193 = v_2495 | ~v_2494;
assign x_21194 = v_2495 | ~v_2431;
assign x_21195 = v_2495 | ~v_2434;
assign x_21196 = v_2495 | ~v_1180;
assign x_21197 = v_2495 | ~v_1181;
assign x_21198 = v_2495 | ~v_183;
assign x_21199 = v_2495 | ~v_167;
assign x_21200 = v_2495 | ~v_166;
assign x_21201 = v_2495 | ~v_165;
assign x_21202 = v_2495 | ~v_159;
assign x_21203 = v_2495 | ~v_146;
assign x_21204 = v_2495 | ~v_145;
assign x_21205 = v_2495 | ~v_144;
assign x_21206 = v_2495 | ~v_142;
assign x_21207 = v_2495 | ~v_61;
assign x_21208 = v_2495 | ~v_58;
assign x_21209 = v_2495 | ~v_54;
assign x_21210 = ~v_89 | ~v_176 | v_2494;
assign x_21211 = ~v_84 | ~v_175 | v_2493;
assign x_21212 = ~v_74 | v_176 | v_2492;
assign x_21213 = ~v_69 | v_175 | v_2491;
assign x_21214 = v_2490 | ~v_2408;
assign x_21215 = v_2490 | ~v_2409;
assign x_21216 = v_2490 | ~v_2410;
assign x_21217 = v_2490 | ~v_2411;
assign x_21218 = v_2490 | ~v_1644;
assign x_21219 = v_2490 | ~v_1645;
assign x_21220 = v_2490 | ~v_1646;
assign x_21221 = v_2490 | ~v_1647;
assign x_21222 = v_2490 | ~v_1700;
assign x_21223 = v_2490 | ~v_1701;
assign x_21224 = v_2490 | ~v_1702;
assign x_21225 = v_2490 | ~v_1703;
assign x_21226 = v_2490 | ~v_1576;
assign x_21227 = v_2490 | ~v_1579;
assign x_21228 = v_2490 | ~v_1161;
assign x_21229 = v_2490 | ~v_1162;
assign x_21230 = v_2490 | ~v_1163;
assign x_21231 = v_2490 | ~v_1164;
assign x_21232 = v_2490 | ~v_2454;
assign x_21233 = v_2490 | ~v_2455;
assign x_21234 = v_2490 | ~v_2456;
assign x_21235 = v_2490 | ~v_2457;
assign x_21236 = v_2490 | ~v_771;
assign x_21237 = v_2490 | ~v_772;
assign x_21238 = v_2490 | ~v_2486;
assign x_21239 = v_2490 | ~v_2487;
assign x_21240 = v_2490 | ~v_2488;
assign x_21241 = v_2490 | ~v_2489;
assign x_21242 = v_2490 | ~v_2416;
assign x_21243 = v_2490 | ~v_2419;
assign x_21244 = v_2490 | ~v_1165;
assign x_21245 = v_2490 | ~v_1166;
assign x_21246 = v_2490 | ~v_182;
assign x_21247 = v_2490 | ~v_163;
assign x_21248 = v_2490 | ~v_162;
assign x_21249 = v_2490 | ~v_161;
assign x_21250 = v_2490 | ~v_155;
assign x_21251 = v_2490 | ~v_138;
assign x_21252 = v_2490 | ~v_137;
assign x_21253 = v_2490 | ~v_136;
assign x_21254 = v_2490 | ~v_134;
assign x_21255 = v_2490 | ~v_18;
assign x_21256 = v_2490 | ~v_15;
assign x_21257 = v_2490 | ~v_11;
assign x_21258 = ~v_47 | ~v_176 | v_2489;
assign x_21259 = ~v_42 | ~v_175 | v_2488;
assign x_21260 = ~v_32 | v_176 | v_2487;
assign x_21261 = ~v_27 | v_175 | v_2486;
assign x_21262 = ~v_2484 | ~v_2479 | ~v_2474 | v_2485;
assign x_21263 = v_2484 | ~v_2438;
assign x_21264 = v_2484 | ~v_2439;
assign x_21265 = v_2484 | ~v_2440;
assign x_21266 = v_2484 | ~v_2441;
assign x_21267 = v_2484 | ~v_1662;
assign x_21268 = v_2484 | ~v_1663;
assign x_21269 = v_2484 | ~v_1664;
assign x_21270 = v_2484 | ~v_1665;
assign x_21271 = v_2484 | ~v_1690;
assign x_21272 = v_2484 | ~v_1691;
assign x_21273 = v_2484 | ~v_1692;
assign x_21274 = v_2484 | ~v_1693;
assign x_21275 = v_2484 | ~v_1626;
assign x_21276 = v_2484 | ~v_1629;
assign x_21277 = v_2484 | ~v_1209;
assign x_21278 = v_2484 | ~v_1210;
assign x_21279 = v_2484 | ~v_1193;
assign x_21280 = v_2484 | ~v_1194;
assign x_21281 = v_2484 | ~v_2464;
assign x_21282 = v_2484 | ~v_2465;
assign x_21283 = v_2484 | ~v_2466;
assign x_21284 = v_2484 | ~v_2467;
assign x_21285 = v_2484 | ~v_927;
assign x_21286 = v_2484 | ~v_928;
assign x_21287 = v_2484 | ~v_2480;
assign x_21288 = v_2484 | ~v_2481;
assign x_21289 = v_2484 | ~v_2482;
assign x_21290 = v_2484 | ~v_2483;
assign x_21291 = v_2484 | ~v_2446;
assign x_21292 = v_2484 | ~v_2449;
assign x_21293 = v_2484 | ~v_1211;
assign x_21294 = v_2484 | ~v_1212;
assign x_21295 = v_2484 | ~v_184;
assign x_21296 = v_2484 | ~v_172;
assign x_21297 = v_2484 | ~v_171;
assign x_21298 = v_2484 | ~v_170;
assign x_21299 = v_2484 | ~v_169;
assign x_21300 = v_2484 | ~v_150;
assign x_21301 = v_2484 | ~v_148;
assign x_21302 = v_2484 | ~v_147;
assign x_21303 = v_2484 | ~v_102;
assign x_21304 = v_2484 | ~v_101;
assign x_21305 = v_2484 | ~v_100;
assign x_21306 = v_2484 | ~v_97;
assign x_21307 = ~v_131 | ~v_141 | v_2483;
assign x_21308 = ~v_126 | ~v_141 | v_2482;
assign x_21309 = ~v_116 | v_141 | v_2481;
assign x_21310 = ~v_111 | v_141 | v_2480;
assign x_21311 = v_2479 | ~v_2423;
assign x_21312 = v_2479 | ~v_2424;
assign x_21313 = v_2479 | ~v_2425;
assign x_21314 = v_2479 | ~v_2426;
assign x_21315 = v_2479 | ~v_1653;
assign x_21316 = v_2479 | ~v_1654;
assign x_21317 = v_2479 | ~v_1655;
assign x_21318 = v_2479 | ~v_1656;
assign x_21319 = v_2479 | ~v_1681;
assign x_21320 = v_2479 | ~v_1682;
assign x_21321 = v_2479 | ~v_1683;
assign x_21322 = v_2479 | ~v_1684;
assign x_21323 = v_2479 | ~v_1601;
assign x_21324 = v_2479 | ~v_1604;
assign x_21325 = v_2479 | ~v_1204;
assign x_21326 = v_2479 | ~v_1205;
assign x_21327 = v_2479 | ~v_1178;
assign x_21328 = v_2479 | ~v_1179;
assign x_21329 = v_2479 | ~v_2459;
assign x_21330 = v_2479 | ~v_2460;
assign x_21331 = v_2479 | ~v_2461;
assign x_21332 = v_2479 | ~v_2462;
assign x_21333 = v_2479 | ~v_912;
assign x_21334 = v_2479 | ~v_913;
assign x_21335 = v_2479 | ~v_2475;
assign x_21336 = v_2479 | ~v_2476;
assign x_21337 = v_2479 | ~v_2477;
assign x_21338 = v_2479 | ~v_2478;
assign x_21339 = v_2479 | ~v_2431;
assign x_21340 = v_2479 | ~v_2434;
assign x_21341 = v_2479 | ~v_1206;
assign x_21342 = v_2479 | ~v_1207;
assign x_21343 = v_2479 | ~v_183;
assign x_21344 = v_2479 | ~v_168;
assign x_21345 = v_2479 | ~v_167;
assign x_21346 = v_2479 | ~v_166;
assign x_21347 = v_2479 | ~v_165;
assign x_21348 = v_2479 | ~v_145;
assign x_21349 = v_2479 | ~v_143;
assign x_21350 = v_2479 | ~v_142;
assign x_21351 = v_2479 | ~v_60;
assign x_21352 = v_2479 | ~v_59;
assign x_21353 = v_2479 | ~v_58;
assign x_21354 = v_2479 | ~v_55;
assign x_21355 = ~v_89 | ~v_141 | v_2478;
assign x_21356 = ~v_84 | ~v_141 | v_2477;
assign x_21357 = ~v_74 | v_141 | v_2476;
assign x_21358 = ~v_69 | v_141 | v_2475;
assign x_21359 = v_2474 | ~v_2408;
assign x_21360 = v_2474 | ~v_2409;
assign x_21361 = v_2474 | ~v_2410;
assign x_21362 = v_2474 | ~v_2411;
assign x_21363 = v_2474 | ~v_1644;
assign x_21364 = v_2474 | ~v_1645;
assign x_21365 = v_2474 | ~v_1646;
assign x_21366 = v_2474 | ~v_1647;
assign x_21367 = v_2474 | ~v_1672;
assign x_21368 = v_2474 | ~v_1673;
assign x_21369 = v_2474 | ~v_1674;
assign x_21370 = v_2474 | ~v_1675;
assign x_21371 = v_2474 | ~v_1576;
assign x_21372 = v_2474 | ~v_1579;
assign x_21373 = v_2474 | ~v_1199;
assign x_21374 = v_2474 | ~v_1200;
assign x_21375 = v_2474 | ~v_1163;
assign x_21376 = v_2474 | ~v_1164;
assign x_21377 = v_2474 | ~v_2454;
assign x_21378 = v_2474 | ~v_2455;
assign x_21379 = v_2474 | ~v_2456;
assign x_21380 = v_2474 | ~v_2457;
assign x_21381 = v_2474 | ~v_897;
assign x_21382 = v_2474 | ~v_898;
assign x_21383 = v_2474 | ~v_2470;
assign x_21384 = v_2474 | ~v_2471;
assign x_21385 = v_2474 | ~v_2472;
assign x_21386 = v_2474 | ~v_2473;
assign x_21387 = v_2474 | ~v_2416;
assign x_21388 = v_2474 | ~v_2419;
assign x_21389 = v_2474 | ~v_1201;
assign x_21390 = v_2474 | ~v_1202;
assign x_21391 = v_2474 | ~v_182;
assign x_21392 = v_2474 | ~v_164;
assign x_21393 = v_2474 | ~v_163;
assign x_21394 = v_2474 | ~v_162;
assign x_21395 = v_2474 | ~v_161;
assign x_21396 = v_2474 | ~v_137;
assign x_21397 = v_2474 | ~v_135;
assign x_21398 = v_2474 | ~v_134;
assign x_21399 = v_2474 | ~v_17;
assign x_21400 = v_2474 | ~v_16;
assign x_21401 = v_2474 | ~v_15;
assign x_21402 = v_2474 | ~v_12;
assign x_21403 = ~v_47 | ~v_141 | v_2473;
assign x_21404 = ~v_42 | ~v_141 | v_2472;
assign x_21405 = ~v_32 | v_141 | v_2471;
assign x_21406 = ~v_27 | v_141 | v_2470;
assign x_21407 = ~v_2468 | ~v_2463 | ~v_2458 | v_2469;
assign x_21408 = v_2468 | ~v_2438;
assign x_21409 = v_2468 | ~v_2439;
assign x_21410 = v_2468 | ~v_2440;
assign x_21411 = v_2468 | ~v_2441;
assign x_21412 = v_2468 | ~v_1662;
assign x_21413 = v_2468 | ~v_1663;
assign x_21414 = v_2468 | ~v_1664;
assign x_21415 = v_2468 | ~v_1665;
assign x_21416 = v_2468 | ~v_1622;
assign x_21417 = v_2468 | ~v_1623;
assign x_21418 = v_2468 | ~v_1624;
assign x_21419 = v_2468 | ~v_1625;
assign x_21420 = v_2468 | ~v_1626;
assign x_21421 = v_2468 | ~v_1629;
assign x_21422 = v_2468 | ~v_1225;
assign x_21423 = v_2468 | ~v_1226;
assign x_21424 = v_2468 | ~v_1227;
assign x_21425 = v_2468 | ~v_1228;
assign x_21426 = v_2468 | ~v_1193;
assign x_21427 = v_2468 | ~v_1194;
assign x_21428 = v_2468 | ~v_2464;
assign x_21429 = v_2468 | ~v_2465;
assign x_21430 = v_2468 | ~v_2466;
assign x_21431 = v_2468 | ~v_2467;
assign x_21432 = v_2468 | ~v_975;
assign x_21433 = v_2468 | ~v_976;
assign x_21434 = v_2468 | ~v_2442;
assign x_21435 = v_2468 | ~v_2443;
assign x_21436 = v_2468 | ~v_2444;
assign x_21437 = v_2468 | ~v_2445;
assign x_21438 = v_2468 | ~v_2446;
assign x_21439 = v_2468 | ~v_2449;
assign x_21440 = v_2468 | ~v_184;
assign x_21441 = v_2468 | ~v_171;
assign x_21442 = v_2468 | ~v_170;
assign x_21443 = v_2468 | ~v_169;
assign x_21444 = v_2468 | ~v_150;
assign x_21445 = v_2468 | ~v_149;
assign x_21446 = v_2468 | ~v_148;
assign x_21447 = v_2468 | ~v_103;
assign x_21448 = v_2468 | ~v_102;
assign x_21449 = v_2468 | ~v_101;
assign x_21450 = v_2468 | ~v_100;
assign x_21451 = v_2468 | ~v_95;
assign x_21452 = ~v_128 | ~v_174 | v_2467;
assign x_21453 = ~v_125 | ~v_173 | v_2466;
assign x_21454 = ~v_113 | v_174 | v_2465;
assign x_21455 = ~v_110 | v_173 | v_2464;
assign x_21456 = v_2463 | ~v_2423;
assign x_21457 = v_2463 | ~v_2424;
assign x_21458 = v_2463 | ~v_2425;
assign x_21459 = v_2463 | ~v_2426;
assign x_21460 = v_2463 | ~v_1653;
assign x_21461 = v_2463 | ~v_1654;
assign x_21462 = v_2463 | ~v_1655;
assign x_21463 = v_2463 | ~v_1656;
assign x_21464 = v_2463 | ~v_1597;
assign x_21465 = v_2463 | ~v_1598;
assign x_21466 = v_2463 | ~v_1599;
assign x_21467 = v_2463 | ~v_1600;
assign x_21468 = v_2463 | ~v_1601;
assign x_21469 = v_2463 | ~v_1604;
assign x_21470 = v_2463 | ~v_1220;
assign x_21471 = v_2463 | ~v_1221;
assign x_21472 = v_2463 | ~v_1222;
assign x_21473 = v_2463 | ~v_1223;
assign x_21474 = v_2463 | ~v_1178;
assign x_21475 = v_2463 | ~v_1179;
assign x_21476 = v_2463 | ~v_2459;
assign x_21477 = v_2463 | ~v_2460;
assign x_21478 = v_2463 | ~v_2461;
assign x_21479 = v_2463 | ~v_2462;
assign x_21480 = v_2463 | ~v_960;
assign x_21481 = v_2463 | ~v_961;
assign x_21482 = v_2463 | ~v_2427;
assign x_21483 = v_2463 | ~v_2428;
assign x_21484 = v_2463 | ~v_2429;
assign x_21485 = v_2463 | ~v_2430;
assign x_21486 = v_2463 | ~v_2431;
assign x_21487 = v_2463 | ~v_2434;
assign x_21488 = v_2463 | ~v_183;
assign x_21489 = v_2463 | ~v_167;
assign x_21490 = v_2463 | ~v_166;
assign x_21491 = v_2463 | ~v_165;
assign x_21492 = v_2463 | ~v_145;
assign x_21493 = v_2463 | ~v_144;
assign x_21494 = v_2463 | ~v_143;
assign x_21495 = v_2463 | ~v_61;
assign x_21496 = v_2463 | ~v_60;
assign x_21497 = v_2463 | ~v_59;
assign x_21498 = v_2463 | ~v_58;
assign x_21499 = v_2463 | ~v_53;
assign x_21500 = ~v_86 | ~v_174 | v_2462;
assign x_21501 = ~v_83 | ~v_173 | v_2461;
assign x_21502 = ~v_71 | v_174 | v_2460;
assign x_21503 = ~v_68 | v_173 | v_2459;
assign x_21504 = v_2458 | ~v_2408;
assign x_21505 = v_2458 | ~v_2409;
assign x_21506 = v_2458 | ~v_2410;
assign x_21507 = v_2458 | ~v_2411;
assign x_21508 = v_2458 | ~v_1644;
assign x_21509 = v_2458 | ~v_1645;
assign x_21510 = v_2458 | ~v_1646;
assign x_21511 = v_2458 | ~v_1647;
assign x_21512 = v_2458 | ~v_1572;
assign x_21513 = v_2458 | ~v_1573;
assign x_21514 = v_2458 | ~v_1574;
assign x_21515 = v_2458 | ~v_1575;
assign x_21516 = v_2458 | ~v_1576;
assign x_21517 = v_2458 | ~v_1579;
assign x_21518 = v_2458 | ~v_1215;
assign x_21519 = v_2458 | ~v_1216;
assign x_21520 = v_2458 | ~v_1217;
assign x_21521 = v_2458 | ~v_1218;
assign x_21522 = v_2458 | ~v_1163;
assign x_21523 = v_2458 | ~v_1164;
assign x_21524 = v_2458 | ~v_2454;
assign x_21525 = v_2458 | ~v_2455;
assign x_21526 = v_2458 | ~v_2456;
assign x_21527 = v_2458 | ~v_2457;
assign x_21528 = v_2458 | ~v_945;
assign x_21529 = v_2458 | ~v_946;
assign x_21530 = v_2458 | ~v_2412;
assign x_21531 = v_2458 | ~v_2413;
assign x_21532 = v_2458 | ~v_2414;
assign x_21533 = v_2458 | ~v_2415;
assign x_21534 = v_2458 | ~v_2416;
assign x_21535 = v_2458 | ~v_2419;
assign x_21536 = v_2458 | ~v_182;
assign x_21537 = v_2458 | ~v_163;
assign x_21538 = v_2458 | ~v_162;
assign x_21539 = v_2458 | ~v_161;
assign x_21540 = v_2458 | ~v_137;
assign x_21541 = v_2458 | ~v_136;
assign x_21542 = v_2458 | ~v_135;
assign x_21543 = v_2458 | ~v_18;
assign x_21544 = v_2458 | ~v_17;
assign x_21545 = v_2458 | ~v_16;
assign x_21546 = v_2458 | ~v_15;
assign x_21547 = v_2458 | ~v_10;
assign x_21548 = ~v_44 | ~v_174 | v_2457;
assign x_21549 = ~v_41 | ~v_173 | v_2456;
assign x_21550 = ~v_29 | v_174 | v_2455;
assign x_21551 = ~v_26 | v_173 | v_2454;
assign x_21552 = ~v_2452 | ~v_2437 | ~v_2422 | v_2453;
assign x_21553 = v_2452 | ~v_2438;
assign x_21554 = v_2452 | ~v_2439;
assign x_21555 = v_2452 | ~v_2440;
assign x_21556 = v_2452 | ~v_2441;
assign x_21557 = v_2452 | ~v_1622;
assign x_21558 = v_2452 | ~v_1623;
assign x_21559 = v_2452 | ~v_1624;
assign x_21560 = v_2452 | ~v_1625;
assign x_21561 = v_2452 | ~v_1626;
assign x_21562 = v_2452 | ~v_1627;
assign x_21563 = v_2452 | ~v_1628;
assign x_21564 = v_2452 | ~v_1629;
assign x_21565 = v_2452 | ~v_1630;
assign x_21566 = v_2452 | ~v_1631;
assign x_21567 = v_2452 | ~v_1147;
assign x_21568 = v_2452 | ~v_1148;
assign x_21569 = v_2452 | ~v_975;
assign x_21570 = v_2452 | ~v_976;
assign x_21571 = v_2452 | ~v_2442;
assign x_21572 = v_2452 | ~v_2443;
assign x_21573 = v_2452 | ~v_2444;
assign x_21574 = v_2452 | ~v_2445;
assign x_21575 = v_2452 | ~v_839;
assign x_21576 = v_2452 | ~v_840;
assign x_21577 = v_2452 | ~v_2446;
assign x_21578 = v_2452 | ~v_2447;
assign x_21579 = v_2452 | ~v_2448;
assign x_21580 = v_2452 | ~v_2449;
assign x_21581 = v_2452 | ~v_2450;
assign x_21582 = v_2452 | ~v_2451;
assign x_21583 = v_2452 | ~v_1149;
assign x_21584 = v_2452 | ~v_1150;
assign x_21585 = v_2452 | ~v_184;
assign x_21586 = v_2452 | ~v_170;
assign x_21587 = v_2452 | ~v_169;
assign x_21588 = v_2452 | ~v_150;
assign x_21589 = v_2452 | ~v_149;
assign x_21590 = v_2452 | ~v_148;
assign x_21591 = v_2452 | ~v_147;
assign x_21592 = v_2452 | ~v_103;
assign x_21593 = v_2452 | ~v_102;
assign x_21594 = v_2452 | ~v_101;
assign x_21595 = v_2452 | ~v_100;
assign x_21596 = v_2452 | ~v_98;
assign x_21597 = ~v_128 | ~v_139 | v_2451;
assign x_21598 = ~v_125 | ~v_140 | v_2450;
assign x_21599 = ~v_124 | ~v_141 | v_2449;
assign x_21600 = ~v_113 | v_139 | v_2448;
assign x_21601 = ~v_110 | v_140 | v_2447;
assign x_21602 = ~v_109 | v_141 | v_2446;
assign x_21603 = ~v_131 | ~v_174 | v_2445;
assign x_21604 = ~v_126 | ~v_173 | v_2444;
assign x_21605 = ~v_116 | v_174 | v_2443;
assign x_21606 = ~v_111 | v_173 | v_2442;
assign x_21607 = ~v_123 | ~v_175 | v_2441;
assign x_21608 = ~v_120 | ~v_176 | v_2440;
assign x_21609 = ~v_108 | v_175 | v_2439;
assign x_21610 = ~v_105 | v_176 | v_2438;
assign x_21611 = v_2437 | ~v_2423;
assign x_21612 = v_2437 | ~v_2424;
assign x_21613 = v_2437 | ~v_2425;
assign x_21614 = v_2437 | ~v_2426;
assign x_21615 = v_2437 | ~v_1597;
assign x_21616 = v_2437 | ~v_1598;
assign x_21617 = v_2437 | ~v_1599;
assign x_21618 = v_2437 | ~v_1600;
assign x_21619 = v_2437 | ~v_1601;
assign x_21620 = v_2437 | ~v_1602;
assign x_21621 = v_2437 | ~v_1603;
assign x_21622 = v_2437 | ~v_1604;
assign x_21623 = v_2437 | ~v_1605;
assign x_21624 = v_2437 | ~v_1606;
assign x_21625 = v_2437 | ~v_1142;
assign x_21626 = v_2437 | ~v_1143;
assign x_21627 = v_2437 | ~v_960;
assign x_21628 = v_2437 | ~v_961;
assign x_21629 = v_2437 | ~v_2427;
assign x_21630 = v_2437 | ~v_2428;
assign x_21631 = v_2437 | ~v_2429;
assign x_21632 = v_2437 | ~v_2430;
assign x_21633 = v_2437 | ~v_806;
assign x_21634 = v_2437 | ~v_2431;
assign x_21635 = v_2437 | ~v_2432;
assign x_21636 = v_2437 | ~v_2433;
assign x_21637 = v_2437 | ~v_2434;
assign x_21638 = v_2437 | ~v_2435;
assign x_21639 = v_2437 | ~v_2436;
assign x_21640 = v_2437 | ~v_807;
assign x_21641 = v_2437 | ~v_1144;
assign x_21642 = v_2437 | ~v_1145;
assign x_21643 = v_2437 | ~v_183;
assign x_21644 = v_2437 | ~v_166;
assign x_21645 = v_2437 | ~v_165;
assign x_21646 = v_2437 | ~v_145;
assign x_21647 = v_2437 | ~v_144;
assign x_21648 = v_2437 | ~v_143;
assign x_21649 = v_2437 | ~v_142;
assign x_21650 = v_2437 | ~v_61;
assign x_21651 = v_2437 | ~v_60;
assign x_21652 = v_2437 | ~v_59;
assign x_21653 = v_2437 | ~v_58;
assign x_21654 = v_2437 | ~v_56;
assign x_21655 = ~v_86 | ~v_139 | v_2436;
assign x_21656 = ~v_83 | ~v_140 | v_2435;
assign x_21657 = ~v_82 | ~v_141 | v_2434;
assign x_21658 = ~v_71 | v_139 | v_2433;
assign x_21659 = ~v_68 | v_140 | v_2432;
assign x_21660 = ~v_67 | v_141 | v_2431;
assign x_21661 = ~v_89 | ~v_174 | v_2430;
assign x_21662 = ~v_84 | ~v_173 | v_2429;
assign x_21663 = ~v_74 | v_174 | v_2428;
assign x_21664 = ~v_69 | v_173 | v_2427;
assign x_21665 = ~v_81 | ~v_175 | v_2426;
assign x_21666 = ~v_78 | ~v_176 | v_2425;
assign x_21667 = ~v_66 | v_175 | v_2424;
assign x_21668 = ~v_63 | v_176 | v_2423;
assign x_21669 = v_2422 | ~v_2408;
assign x_21670 = v_2422 | ~v_2409;
assign x_21671 = v_2422 | ~v_2410;
assign x_21672 = v_2422 | ~v_2411;
assign x_21673 = v_2422 | ~v_1572;
assign x_21674 = v_2422 | ~v_1573;
assign x_21675 = v_2422 | ~v_1574;
assign x_21676 = v_2422 | ~v_1575;
assign x_21677 = v_2422 | ~v_1576;
assign x_21678 = v_2422 | ~v_1577;
assign x_21679 = v_2422 | ~v_1578;
assign x_21680 = v_2422 | ~v_1579;
assign x_21681 = v_2422 | ~v_1580;
assign x_21682 = v_2422 | ~v_1581;
assign x_21683 = v_2422 | ~v_1137;
assign x_21684 = v_2422 | ~v_1138;
assign x_21685 = v_2422 | ~v_945;
assign x_21686 = v_2422 | ~v_946;
assign x_21687 = v_2422 | ~v_2412;
assign x_21688 = v_2422 | ~v_2413;
assign x_21689 = v_2422 | ~v_2414;
assign x_21690 = v_2422 | ~v_2415;
assign x_21691 = v_2422 | ~v_773;
assign x_21692 = v_2422 | ~v_774;
assign x_21693 = v_2422 | ~v_2416;
assign x_21694 = v_2422 | ~v_2417;
assign x_21695 = v_2422 | ~v_2418;
assign x_21696 = v_2422 | ~v_2419;
assign x_21697 = v_2422 | ~v_2420;
assign x_21698 = v_2422 | ~v_2421;
assign x_21699 = v_2422 | ~v_1139;
assign x_21700 = v_2422 | ~v_1140;
assign x_21701 = v_2422 | ~v_182;
assign x_21702 = v_2422 | ~v_162;
assign x_21703 = v_2422 | ~v_161;
assign x_21704 = v_2422 | ~v_137;
assign x_21705 = v_2422 | ~v_136;
assign x_21706 = v_2422 | ~v_135;
assign x_21707 = v_2422 | ~v_134;
assign x_21708 = v_2422 | ~v_18;
assign x_21709 = v_2422 | ~v_17;
assign x_21710 = v_2422 | ~v_16;
assign x_21711 = v_2422 | ~v_15;
assign x_21712 = v_2422 | ~v_13;
assign x_21713 = ~v_44 | ~v_139 | v_2421;
assign x_21714 = ~v_41 | ~v_140 | v_2420;
assign x_21715 = ~v_40 | ~v_141 | v_2419;
assign x_21716 = ~v_29 | v_139 | v_2418;
assign x_21717 = ~v_26 | v_140 | v_2417;
assign x_21718 = ~v_25 | v_141 | v_2416;
assign x_21719 = ~v_47 | ~v_174 | v_2415;
assign x_21720 = ~v_42 | ~v_173 | v_2414;
assign x_21721 = ~v_32 | v_174 | v_2413;
assign x_21722 = ~v_27 | v_173 | v_2412;
assign x_21723 = ~v_39 | ~v_175 | v_2411;
assign x_21724 = ~v_36 | ~v_176 | v_2410;
assign x_21725 = ~v_24 | v_175 | v_2409;
assign x_21726 = ~v_21 | v_176 | v_2408;
assign x_21727 = v_2407 | ~v_2406;
assign x_21728 = v_2407 | ~v_727;
assign x_21729 = v_140 | v_139 | ~v_2405 | ~v_2404 | v_2406;
assign x_21730 = v_2405 | ~v_737;
assign x_21731 = v_2405 | ~v_731;
assign x_21732 = v_2404 | ~v_735;
assign x_21733 = v_2404 | ~v_727;
assign x_21734 = v_2403 | ~v_1562;
assign x_21735 = v_2403 | ~v_730;
assign x_21736 = ~v_725 | ~v_724 | ~v_723 | ~v_722 | ~v_2401 | ~v_2397 | ~v_2393 | ~v_2389 | ~v_2385 | ~v_2369 | ~v_2365 | ~v_2361 | ~v_2357 | ~v_2353 | ~v_2337 | ~v_2333 | ~v_2317 | ~v_2301 | ~v_2285 | ~v_2269 | ~v_2223 | v_2402;
assign x_21737 = v_2401 | ~v_2398;
assign x_21738 = v_2401 | ~v_2399;
assign x_21739 = v_2401 | ~v_2400;
assign x_21740 = v_98 | v_103 | v_101 | v_100 | v_95 | v_99 | v_102 | ~v_719 | ~v_718 | v_170 | v_169 | v_149 | v_148 | v_184 | ~v_2331 | ~v_2267 | ~v_2330 | ~v_2266 | ~v_2265 | ~v_2329 | ~v_2264 | ~v_2328 | ~v_2263 | ~v_2262 | ~v_483 | ~v_717 | ~v_299 | ~v_482 | ~v_716 | ~v_298 | ~v_1460 | ~v_1342 | ~v_1459 | ~v_1341 | ~v_1340 | ~v_1458 | ~v_1339 | ~v_1457 | ~v_1338 | ~v_1337 | ~v_2257 | ~v_2256 | ~v_2255 | ~v_2254 | v_2400;
assign x_21741 = v_53 | v_56 | v_61 | v_60 | v_59 | v_58 | v_57 | ~v_714 | ~v_713 | v_144 | v_143 | v_166 | v_165 | v_183 | ~v_266 | ~v_2326 | ~v_2252 | ~v_2325 | ~v_2251 | ~v_2250 | ~v_2324 | ~v_2249 | ~v_2323 | ~v_2248 | ~v_2247 | ~v_468 | ~v_712 | ~v_467 | ~v_711 | ~v_265 | ~v_1451 | ~v_1317 | ~v_1450 | ~v_1316 | ~v_1315 | ~v_1449 | ~v_1314 | ~v_1448 | ~v_1313 | ~v_1312 | ~v_2242 | ~v_2241 | ~v_2240 | ~v_2239 | v_2399;
assign x_21742 = v_13 | v_18 | v_17 | v_16 | v_15 | v_14 | v_10 | ~v_453 | ~v_709 | ~v_452 | ~v_708 | v_136 | v_135 | ~v_707 | ~v_706 | v_162 | v_161 | v_182 | ~v_2321 | ~v_2237 | ~v_2320 | ~v_2236 | ~v_2235 | ~v_2319 | ~v_2234 | ~v_2318 | ~v_2233 | ~v_2232 | ~v_233 | ~v_232 | ~v_1442 | ~v_1292 | ~v_1441 | ~v_1291 | ~v_1290 | ~v_1440 | ~v_1289 | ~v_1439 | ~v_1288 | ~v_1287 | ~v_2227 | ~v_2226 | ~v_2225 | ~v_2224 | v_2398;
assign x_21743 = v_2397 | ~v_2394;
assign x_21744 = v_2397 | ~v_2395;
assign x_21745 = v_2397 | ~v_2396;
assign x_21746 = v_103 | v_101 | v_99 | v_93 | v_102 | v_171 | v_170 | v_149 | v_148 | v_147 | v_184 | v_181 | ~v_2331 | ~v_2330 | ~v_2265 | ~v_2329 | ~v_2328 | ~v_2262 | ~v_483 | ~v_482 | ~v_2383 | ~v_2382 | ~v_2381 | ~v_2380 | ~v_481 | ~v_480 | ~v_345 | ~v_479 | ~v_478 | ~v_344 | ~v_1460 | ~v_1459 | ~v_1340 | ~v_1458 | ~v_1457 | ~v_1337 | ~v_1536 | ~v_1535 | ~v_1534 | ~v_1533 | ~v_2257 | ~v_2256 | ~v_2255 | ~v_2254 | v_2396;
assign x_21747 = v_61 | v_51 | v_60 | v_59 | v_57 | v_144 | v_180 | v_143 | v_142 | v_167 | v_166 | v_183 | ~v_2326 | ~v_2325 | ~v_2250 | ~v_2324 | ~v_2323 | ~v_2247 | ~v_468 | ~v_467 | ~v_2378 | ~v_2377 | ~v_2376 | ~v_2375 | ~v_466 | ~v_465 | ~v_330 | ~v_464 | ~v_463 | ~v_329 | ~v_1451 | ~v_1450 | ~v_1315 | ~v_1449 | ~v_1448 | ~v_1312 | ~v_1527 | ~v_1526 | ~v_1525 | ~v_1524 | ~v_2242 | ~v_2241 | ~v_2240 | ~v_2239 | v_2395;
assign x_21748 = v_18 | v_17 | v_16 | v_8 | v_14 | ~v_453 | ~v_452 | v_136 | v_135 | v_134 | v_179 | v_163 | v_162 | v_182 | ~v_2321 | ~v_2320 | ~v_2235 | ~v_2319 | ~v_2318 | ~v_2232 | ~v_2373 | ~v_2372 | ~v_2371 | ~v_2370 | ~v_451 | ~v_450 | ~v_315 | ~v_449 | ~v_448 | ~v_314 | ~v_1442 | ~v_1441 | ~v_1290 | ~v_1440 | ~v_1439 | ~v_1287 | ~v_1518 | ~v_1517 | ~v_1516 | ~v_1515 | ~v_2227 | ~v_2226 | ~v_2225 | ~v_2224 | v_2394;
assign x_21749 = v_2393 | ~v_2390;
assign x_21750 = v_2393 | ~v_2391;
assign x_21751 = v_2393 | ~v_2392;
assign x_21752 = v_103 | v_96 | v_95 | v_93 | v_102 | v_171 | v_170 | v_160 | v_150 | v_149 | v_184 | v_181 | ~v_2265 | ~v_2262 | ~v_2315 | ~v_2314 | ~v_2313 | ~v_2312 | ~v_297 | ~v_296 | ~v_2383 | ~v_2382 | ~v_2381 | ~v_2380 | ~v_345 | ~v_344 | ~v_343 | ~v_342 | ~v_341 | ~v_340 | ~v_1340 | ~v_1337 | ~v_1536 | ~v_1535 | ~v_1534 | ~v_1533 | ~v_1432 | ~v_1431 | ~v_1430 | ~v_1429 | ~v_2257 | ~v_2256 | ~v_2255 | ~v_2254 | v_2392;
assign x_21753 = v_54 | v_53 | v_61 | v_51 | v_60 | v_144 | v_180 | v_159 | v_145 | v_167 | v_166 | v_183 | ~v_2250 | ~v_2247 | ~v_2310 | ~v_2309 | ~v_2308 | ~v_2307 | ~v_264 | ~v_263 | ~v_2378 | ~v_2377 | ~v_2376 | ~v_2375 | ~v_330 | ~v_329 | ~v_328 | ~v_327 | ~v_326 | ~v_325 | ~v_1315 | ~v_1312 | ~v_1527 | ~v_1526 | ~v_1525 | ~v_1524 | ~v_1423 | ~v_1422 | ~v_1421 | ~v_1420 | ~v_2242 | ~v_2241 | ~v_2240 | ~v_2239 | v_2391;
assign x_21754 = v_18 | v_17 | v_8 | v_11 | v_10 | v_136 | v_137 | v_179 | v_163 | v_162 | v_155 | v_182 | ~v_2235 | ~v_2232 | ~v_2305 | ~v_2304 | ~v_2303 | ~v_2302 | ~v_231 | ~v_230 | ~v_2373 | ~v_2372 | ~v_2371 | ~v_2370 | ~v_315 | ~v_314 | ~v_313 | ~v_312 | ~v_311 | ~v_310 | ~v_1290 | ~v_1287 | ~v_1518 | ~v_1517 | ~v_1516 | ~v_1515 | ~v_1414 | ~v_1413 | ~v_1412 | ~v_1411 | ~v_2227 | ~v_2226 | ~v_2225 | ~v_2224 | v_2390;
assign x_21755 = v_2389 | ~v_2386;
assign x_21756 = v_2389 | ~v_2387;
assign x_21757 = v_2389 | ~v_2388;
assign x_21758 = v_103 | v_101 | v_97 | v_93 | v_102 | v_171 | v_170 | v_150 | v_148 | v_147 | v_184 | v_181 | ~v_391 | ~v_390 | ~v_2265 | ~v_2262 | ~v_2299 | ~v_2298 | ~v_2297 | ~v_2296 | ~v_387 | ~v_386 | ~v_2383 | ~v_2382 | ~v_2381 | ~v_2380 | ~v_345 | ~v_344 | ~v_385 | ~v_384 | ~v_1340 | ~v_1337 | ~v_1536 | ~v_1535 | ~v_1534 | ~v_1533 | ~v_1404 | ~v_1403 | ~v_1402 | ~v_1401 | ~v_2257 | ~v_2256 | ~v_2255 | ~v_2254 | v_2388;
assign x_21759 = v_55 | v_61 | v_51 | v_60 | v_59 | v_180 | v_145 | v_143 | v_142 | v_167 | v_166 | v_183 | ~v_376 | ~v_375 | ~v_2250 | ~v_2247 | ~v_2294 | ~v_2293 | ~v_2292 | ~v_2291 | ~v_372 | ~v_371 | ~v_2378 | ~v_2377 | ~v_2376 | ~v_2375 | ~v_330 | ~v_329 | ~v_370 | ~v_369 | ~v_1315 | ~v_1312 | ~v_1527 | ~v_1526 | ~v_1525 | ~v_1524 | ~v_1395 | ~v_1394 | ~v_1393 | ~v_1392 | ~v_2242 | ~v_2241 | ~v_2240 | ~v_2239 | v_2387;
assign x_21760 = v_18 | v_17 | v_16 | v_8 | v_12 | v_135 | v_134 | v_137 | v_179 | v_163 | v_162 | v_182 | ~v_361 | ~v_360 | ~v_2235 | ~v_2232 | ~v_2289 | ~v_2288 | ~v_2287 | ~v_2286 | ~v_357 | ~v_356 | ~v_2373 | ~v_2372 | ~v_2371 | ~v_2370 | ~v_315 | ~v_314 | ~v_355 | ~v_354 | ~v_1290 | ~v_1287 | ~v_1518 | ~v_1517 | ~v_1516 | ~v_1515 | ~v_1386 | ~v_1385 | ~v_1384 | ~v_1383 | ~v_2227 | ~v_2226 | ~v_2225 | ~v_2224 | v_2386;
assign x_21761 = v_2385 | ~v_2374;
assign x_21762 = v_2385 | ~v_2379;
assign x_21763 = v_2385 | ~v_2384;
assign x_21764 = v_101 | v_93 | v_102 | v_172 | v_171 | v_170 | v_150 | v_149 | v_148 | v_147 | v_184 | v_181 | ~v_437 | ~v_436 | ~v_2265 | ~v_2262 | ~v_2261 | ~v_2260 | ~v_2259 | ~v_2258 | ~v_435 | ~v_434 | ~v_2383 | ~v_2382 | ~v_2381 | ~v_2380 | ~v_345 | ~v_344 | ~v_433 | ~v_432 | ~v_1340 | ~v_1337 | ~v_1536 | ~v_1535 | ~v_1534 | ~v_1533 | ~v_1336 | ~v_1335 | ~v_1334 | ~v_1333 | ~v_2257 | ~v_2256 | ~v_2255 | ~v_2254 | v_2384;
assign x_21765 = v_2383 | v_176;
assign x_21766 = v_2383 | v_128;
assign x_21767 = v_2382 | v_175;
assign x_21768 = v_2382 | v_125;
assign x_21769 = v_2381 | ~v_176;
assign x_21770 = v_2381 | v_113;
assign x_21771 = v_2380 | ~v_175;
assign x_21772 = v_2380 | v_110;
assign x_21773 = v_51 | v_60 | v_59 | v_144 | v_180 | v_145 | v_143 | v_142 | v_168 | v_167 | v_166 | v_183 | ~v_422 | ~v_421 | ~v_2250 | ~v_2247 | ~v_2246 | ~v_2245 | ~v_2244 | ~v_2243 | ~v_420 | ~v_419 | ~v_2378 | ~v_2377 | ~v_2376 | ~v_2375 | ~v_330 | ~v_329 | ~v_418 | ~v_417 | ~v_1315 | ~v_1312 | ~v_1527 | ~v_1526 | ~v_1525 | ~v_1524 | ~v_1311 | ~v_1310 | ~v_1309 | ~v_1308 | ~v_2242 | ~v_2241 | ~v_2240 | ~v_2239 | v_2379;
assign x_21774 = v_2378 | v_176;
assign x_21775 = v_2378 | v_86;
assign x_21776 = v_2377 | v_175;
assign x_21777 = v_2377 | v_83;
assign x_21778 = v_2376 | ~v_176;
assign x_21779 = v_2376 | v_71;
assign x_21780 = v_2375 | ~v_175;
assign x_21781 = v_2375 | v_68;
assign x_21782 = v_17 | v_16 | v_8 | v_136 | v_135 | v_134 | v_137 | v_179 | v_164 | v_163 | v_162 | v_182 | ~v_407 | ~v_406 | ~v_2235 | ~v_2232 | ~v_2231 | ~v_2230 | ~v_2229 | ~v_2228 | ~v_405 | ~v_404 | ~v_2373 | ~v_2372 | ~v_2371 | ~v_2370 | ~v_315 | ~v_314 | ~v_403 | ~v_402 | ~v_1290 | ~v_1287 | ~v_1518 | ~v_1517 | ~v_1516 | ~v_1515 | ~v_1286 | ~v_1285 | ~v_1284 | ~v_1283 | ~v_2227 | ~v_2226 | ~v_2225 | ~v_2224 | v_2374;
assign x_21783 = v_2373 | v_176;
assign x_21784 = v_2373 | v_44;
assign x_21785 = v_2372 | v_175;
assign x_21786 = v_2372 | v_41;
assign x_21787 = v_2371 | ~v_176;
assign x_21788 = v_2371 | v_29;
assign x_21789 = v_2370 | ~v_175;
assign x_21790 = v_2370 | v_26;
assign x_21791 = v_2369 | ~v_2366;
assign x_21792 = v_2369 | ~v_2367;
assign x_21793 = v_2369 | ~v_2368;
assign x_21794 = v_98 | v_103 | v_96 | v_100 | v_102 | v_170 | v_169 | v_160 | v_150 | v_149 | v_147 | v_184 | ~v_2267 | ~v_2266 | ~v_2265 | ~v_2264 | ~v_2263 | ~v_2262 | ~v_299 | ~v_298 | ~v_2315 | ~v_2314 | ~v_2313 | ~v_2312 | ~v_297 | ~v_296 | ~v_295 | ~v_294 | ~v_293 | ~v_292 | ~v_1342 | ~v_1341 | ~v_1340 | ~v_1339 | ~v_1338 | ~v_1337 | ~v_1432 | ~v_1431 | ~v_1430 | ~v_1429 | ~v_2257 | ~v_2256 | ~v_2255 | ~v_2254 | v_2368;
assign x_21795 = v_54 | v_56 | v_61 | v_60 | v_58 | v_144 | v_159 | v_145 | v_142 | v_166 | v_165 | v_183 | ~v_266 | ~v_2252 | ~v_2251 | ~v_2250 | ~v_2249 | ~v_2248 | ~v_2247 | ~v_265 | ~v_2310 | ~v_2309 | ~v_2308 | ~v_2307 | ~v_264 | ~v_263 | ~v_262 | ~v_261 | ~v_260 | ~v_259 | ~v_1317 | ~v_1316 | ~v_1315 | ~v_1314 | ~v_1313 | ~v_1312 | ~v_1423 | ~v_1422 | ~v_1421 | ~v_1420 | ~v_2242 | ~v_2241 | ~v_2240 | ~v_2239 | v_2367;
assign x_21796 = v_13 | v_18 | v_17 | v_15 | v_11 | v_136 | v_134 | v_137 | v_162 | v_161 | v_155 | v_182 | ~v_2237 | ~v_2236 | ~v_2235 | ~v_2234 | ~v_2233 | ~v_2232 | ~v_233 | ~v_232 | ~v_2305 | ~v_2304 | ~v_2303 | ~v_2302 | ~v_231 | ~v_230 | ~v_229 | ~v_228 | ~v_227 | ~v_226 | ~v_1292 | ~v_1291 | ~v_1290 | ~v_1289 | ~v_1288 | ~v_1287 | ~v_1414 | ~v_1413 | ~v_1412 | ~v_1411 | ~v_2227 | ~v_2226 | ~v_2225 | ~v_2224 | v_2366;
assign x_21797 = v_2365 | ~v_2362;
assign x_21798 = v_2365 | ~v_2363;
assign x_21799 = v_2365 | ~v_2364;
assign x_21800 = v_101 | v_100 | v_94 | v_99 | v_102 | v_172 | v_171 | v_169 | v_149 | v_148 | v_147 | v_184 | ~v_2331 | ~v_2330 | ~v_2265 | ~v_2329 | ~v_2328 | ~v_2262 | ~v_483 | ~v_482 | ~v_2351 | ~v_2350 | ~v_2349 | ~v_2348 | ~v_593 | ~v_592 | ~v_545 | ~v_591 | ~v_590 | ~v_544 | ~v_1460 | ~v_1459 | ~v_1340 | ~v_1458 | ~v_1457 | ~v_1337 | ~v_1492 | ~v_1491 | ~v_1490 | ~v_1489 | ~v_2257 | ~v_2256 | ~v_2255 | ~v_2254 | v_2364;
assign x_21801 = v_52 | v_60 | v_59 | v_58 | v_57 | v_144 | v_143 | v_142 | v_168 | v_167 | v_165 | v_183 | ~v_2326 | ~v_2325 | ~v_2250 | ~v_2324 | ~v_2323 | ~v_2247 | ~v_468 | ~v_467 | ~v_2346 | ~v_2345 | ~v_2344 | ~v_2343 | ~v_588 | ~v_587 | ~v_530 | ~v_586 | ~v_585 | ~v_529 | ~v_1451 | ~v_1450 | ~v_1315 | ~v_1449 | ~v_1448 | ~v_1312 | ~v_1483 | ~v_1482 | ~v_1481 | ~v_1480 | ~v_2242 | ~v_2241 | ~v_2240 | ~v_2239 | v_2363;
assign x_21802 = v_9 | v_17 | v_16 | v_15 | v_14 | ~v_453 | ~v_452 | v_136 | v_135 | v_134 | v_164 | v_163 | v_161 | v_182 | ~v_2321 | ~v_2320 | ~v_2235 | ~v_2319 | ~v_2318 | ~v_2232 | ~v_2341 | ~v_2340 | ~v_2339 | ~v_2338 | ~v_583 | ~v_582 | ~v_515 | ~v_581 | ~v_580 | ~v_514 | ~v_1442 | ~v_1441 | ~v_1290 | ~v_1440 | ~v_1439 | ~v_1287 | ~v_1474 | ~v_1473 | ~v_1472 | ~v_1471 | ~v_2227 | ~v_2226 | ~v_2225 | ~v_2224 | v_2362;
assign x_21803 = v_2361 | ~v_2358;
assign x_21804 = v_2361 | ~v_2359;
assign x_21805 = v_2361 | ~v_2360;
assign x_21806 = v_103 | v_96 | v_100 | v_94 | v_102 | v_171 | v_169 | v_160 | v_150 | v_149 | v_147 | v_184 | ~v_2265 | ~v_2262 | ~v_2351 | ~v_2350 | ~v_2349 | ~v_2348 | ~v_545 | ~v_544 | ~v_2315 | ~v_2314 | ~v_2313 | ~v_2312 | ~v_543 | ~v_542 | ~v_541 | ~v_540 | ~v_297 | ~v_296 | ~v_1340 | ~v_1337 | ~v_1432 | ~v_1431 | ~v_1430 | ~v_1429 | ~v_1492 | ~v_1491 | ~v_1490 | ~v_1489 | ~v_2257 | ~v_2256 | ~v_2255 | ~v_2254 | v_2360;
assign x_21807 = v_54 | v_61 | v_52 | v_60 | v_58 | v_144 | v_159 | v_145 | v_142 | v_167 | v_165 | v_183 | ~v_2250 | ~v_2247 | ~v_2346 | ~v_2345 | ~v_2344 | ~v_2343 | ~v_530 | ~v_529 | ~v_2310 | ~v_2309 | ~v_2308 | ~v_2307 | ~v_528 | ~v_527 | ~v_526 | ~v_525 | ~v_264 | ~v_263 | ~v_1315 | ~v_1312 | ~v_1423 | ~v_1422 | ~v_1421 | ~v_1420 | ~v_1483 | ~v_1482 | ~v_1481 | ~v_1480 | ~v_2242 | ~v_2241 | ~v_2240 | ~v_2239 | v_2359;
assign x_21808 = v_9 | v_18 | v_17 | v_15 | v_11 | v_136 | v_134 | v_137 | v_163 | v_161 | v_155 | v_182 | ~v_2235 | ~v_2232 | ~v_2341 | ~v_2340 | ~v_2339 | ~v_2338 | ~v_515 | ~v_514 | ~v_2305 | ~v_2304 | ~v_2303 | ~v_2302 | ~v_513 | ~v_512 | ~v_511 | ~v_510 | ~v_231 | ~v_230 | ~v_1290 | ~v_1287 | ~v_1414 | ~v_1413 | ~v_1412 | ~v_1411 | ~v_1474 | ~v_1473 | ~v_1472 | ~v_1471 | ~v_2227 | ~v_2226 | ~v_2225 | ~v_2224 | v_2358;
assign x_21809 = v_2357 | ~v_2354;
assign x_21810 = v_2357 | ~v_2355;
assign x_21811 = v_2357 | ~v_2356;
assign x_21812 = v_103 | v_101 | v_97 | v_100 | v_95 | v_94 | v_102 | v_171 | v_169 | v_150 | v_148 | v_184 | ~v_2265 | ~v_2262 | ~v_2351 | ~v_2350 | ~v_2349 | ~v_2348 | ~v_545 | ~v_544 | ~v_2299 | ~v_2298 | ~v_2297 | ~v_2296 | ~v_561 | ~v_560 | ~v_559 | ~v_558 | ~v_387 | ~v_386 | ~v_1340 | ~v_1337 | ~v_1404 | ~v_1403 | ~v_1402 | ~v_1401 | ~v_1492 | ~v_1491 | ~v_1490 | ~v_1489 | ~v_2257 | ~v_2256 | ~v_2255 | ~v_2254 | v_2356;
assign x_21813 = v_53 | v_55 | v_61 | v_52 | v_60 | v_59 | v_58 | v_145 | v_143 | v_167 | v_165 | v_183 | ~v_2250 | ~v_2247 | ~v_2346 | ~v_2345 | ~v_2344 | ~v_2343 | ~v_530 | ~v_529 | ~v_2294 | ~v_2293 | ~v_2292 | ~v_2291 | ~v_556 | ~v_555 | ~v_554 | ~v_553 | ~v_372 | ~v_371 | ~v_1315 | ~v_1312 | ~v_1395 | ~v_1394 | ~v_1393 | ~v_1392 | ~v_1483 | ~v_1482 | ~v_1481 | ~v_1480 | ~v_2242 | ~v_2241 | ~v_2240 | ~v_2239 | v_2355;
assign x_21814 = v_9 | v_18 | v_17 | v_16 | v_15 | v_12 | v_10 | v_135 | v_137 | v_163 | v_161 | v_182 | ~v_2235 | ~v_2232 | ~v_2341 | ~v_2340 | ~v_2339 | ~v_2338 | ~v_515 | ~v_514 | ~v_2289 | ~v_2288 | ~v_2287 | ~v_2286 | ~v_551 | ~v_550 | ~v_549 | ~v_548 | ~v_357 | ~v_356 | ~v_1290 | ~v_1287 | ~v_1386 | ~v_1385 | ~v_1384 | ~v_1383 | ~v_1474 | ~v_1473 | ~v_1472 | ~v_1471 | ~v_2227 | ~v_2226 | ~v_2225 | ~v_2224 | v_2354;
assign x_21815 = v_2353 | ~v_2342;
assign x_21816 = v_2353 | ~v_2347;
assign x_21817 = v_2353 | ~v_2352;
assign x_21818 = v_103 | v_101 | v_100 | v_94 | v_151 | v_171 | v_169 | v_150 | v_149 | v_148 | v_147 | v_184 | ~v_577 | ~v_576 | ~v_2265 | ~v_2262 | ~v_2351 | ~v_2350 | ~v_2349 | ~v_2348 | ~v_545 | ~v_544 | ~v_2261 | ~v_2260 | ~v_2259 | ~v_2258 | ~v_575 | ~v_574 | ~v_435 | ~v_434 | ~v_1340 | ~v_1337 | ~v_1336 | ~v_1335 | ~v_1334 | ~v_1333 | ~v_1492 | ~v_1491 | ~v_1490 | ~v_1489 | ~v_2257 | ~v_2256 | ~v_2255 | ~v_2254 | v_2352;
assign x_21819 = v_2351 | v_141;
assign x_21820 = v_2351 | v_128;
assign x_21821 = v_2350 | v_141;
assign x_21822 = v_2350 | v_125;
assign x_21823 = v_2349 | ~v_141;
assign x_21824 = v_2349 | v_113;
assign x_21825 = v_2348 | ~v_141;
assign x_21826 = v_2348 | v_110;
assign x_21827 = v_61 | v_52 | v_59 | v_58 | v_144 | v_145 | v_143 | v_142 | v_167 | v_165 | v_146 | v_183 | ~v_572 | ~v_571 | ~v_2250 | ~v_2247 | ~v_2346 | ~v_2345 | ~v_2344 | ~v_2343 | ~v_530 | ~v_529 | ~v_2246 | ~v_2245 | ~v_2244 | ~v_2243 | ~v_570 | ~v_569 | ~v_420 | ~v_419 | ~v_1315 | ~v_1312 | ~v_1311 | ~v_1310 | ~v_1309 | ~v_1308 | ~v_1483 | ~v_1482 | ~v_1481 | ~v_1480 | ~v_2242 | ~v_2241 | ~v_2240 | ~v_2239 | v_2347;
assign x_21828 = v_2346 | v_141;
assign x_21829 = v_2346 | v_86;
assign x_21830 = v_2345 | v_141;
assign x_21831 = v_2345 | v_83;
assign x_21832 = v_2344 | ~v_141;
assign x_21833 = v_2344 | v_71;
assign x_21834 = v_2343 | ~v_141;
assign x_21835 = v_2343 | v_68;
assign x_21836 = v_9 | v_18 | v_16 | v_15 | v_136 | v_135 | v_134 | v_137 | v_138 | v_163 | v_161 | v_182 | ~v_567 | ~v_566 | ~v_2235 | ~v_2232 | ~v_2341 | ~v_2340 | ~v_2339 | ~v_2338 | ~v_515 | ~v_514 | ~v_2231 | ~v_2230 | ~v_2229 | ~v_2228 | ~v_565 | ~v_564 | ~v_405 | ~v_404 | ~v_1290 | ~v_1287 | ~v_1286 | ~v_1285 | ~v_1284 | ~v_1283 | ~v_1474 | ~v_1473 | ~v_1472 | ~v_1471 | ~v_2227 | ~v_2226 | ~v_2225 | ~v_2224 | v_2342;
assign x_21837 = v_2341 | v_141;
assign x_21838 = v_2341 | v_44;
assign x_21839 = v_2340 | v_141;
assign x_21840 = v_2340 | v_41;
assign x_21841 = v_2339 | ~v_141;
assign x_21842 = v_2339 | v_29;
assign x_21843 = v_2338 | ~v_141;
assign x_21844 = v_2338 | v_26;
assign x_21845 = v_2337 | ~v_2334;
assign x_21846 = v_2337 | ~v_2335;
assign x_21847 = v_2337 | ~v_2336;
assign x_21848 = v_98 | v_103 | v_101 | v_97 | v_100 | v_151 | v_170 | v_169 | v_150 | v_148 | v_147 | v_184 | ~v_2267 | ~v_2266 | ~v_2265 | ~v_2264 | ~v_2263 | ~v_2262 | ~v_299 | ~v_298 | ~v_2299 | ~v_2298 | ~v_2297 | ~v_2296 | ~v_387 | ~v_386 | ~v_499 | ~v_498 | ~v_497 | ~v_496 | ~v_1342 | ~v_1341 | ~v_1340 | ~v_1339 | ~v_1338 | ~v_1337 | ~v_1404 | ~v_1403 | ~v_1402 | ~v_1401 | ~v_2257 | ~v_2256 | ~v_2255 | ~v_2254 | v_2336;
assign x_21849 = v_56 | v_55 | v_61 | v_59 | v_58 | v_145 | v_143 | v_142 | v_166 | v_165 | v_146 | v_183 | ~v_266 | ~v_2252 | ~v_2251 | ~v_2250 | ~v_2249 | ~v_2248 | ~v_2247 | ~v_265 | ~v_2294 | ~v_2293 | ~v_2292 | ~v_2291 | ~v_372 | ~v_371 | ~v_494 | ~v_493 | ~v_492 | ~v_491 | ~v_1317 | ~v_1316 | ~v_1315 | ~v_1314 | ~v_1313 | ~v_1312 | ~v_1395 | ~v_1394 | ~v_1393 | ~v_1392 | ~v_2242 | ~v_2241 | ~v_2240 | ~v_2239 | v_2335;
assign x_21850 = v_13 | v_18 | v_16 | v_15 | v_12 | v_135 | v_134 | v_137 | v_138 | v_162 | v_161 | v_182 | ~v_2237 | ~v_2236 | ~v_2235 | ~v_2234 | ~v_2233 | ~v_2232 | ~v_233 | ~v_232 | ~v_2289 | ~v_2288 | ~v_2287 | ~v_2286 | ~v_357 | ~v_356 | ~v_489 | ~v_488 | ~v_487 | ~v_486 | ~v_1292 | ~v_1291 | ~v_1290 | ~v_1289 | ~v_1288 | ~v_1287 | ~v_1386 | ~v_1385 | ~v_1384 | ~v_1383 | ~v_2227 | ~v_2226 | ~v_2225 | ~v_2224 | v_2334;
assign x_21851 = v_2333 | ~v_2322;
assign x_21852 = v_2333 | ~v_2327;
assign x_21853 = v_2333 | ~v_2332;
assign x_21854 = v_103 | v_101 | v_100 | v_99 | v_102 | v_171 | v_170 | v_169 | v_149 | v_148 | v_147 | v_184 | ~v_703 | ~v_702 | ~v_2331 | ~v_2330 | ~v_2265 | ~v_2329 | ~v_2328 | ~v_2262 | ~v_483 | ~v_482 | ~v_2283 | ~v_2282 | ~v_2281 | ~v_2280 | ~v_701 | ~v_653 | ~v_700 | ~v_652 | ~v_1460 | ~v_1459 | ~v_1340 | ~v_1458 | ~v_1457 | ~v_1337 | ~v_1376 | ~v_1375 | ~v_1374 | ~v_1373 | ~v_2257 | ~v_2256 | ~v_2255 | ~v_2254 | v_2332;
assign x_21855 = v_2331 | v_139;
assign x_21856 = v_2331 | v_131;
assign x_21857 = v_2330 | v_140;
assign x_21858 = v_2330 | v_126;
assign x_21859 = v_2329 | ~v_139;
assign x_21860 = v_2329 | v_116;
assign x_21861 = v_2328 | ~v_140;
assign x_21862 = v_2328 | v_111;
assign x_21863 = v_61 | v_60 | v_59 | v_58 | v_57 | v_144 | v_143 | v_142 | v_167 | v_166 | v_165 | v_183 | ~v_698 | ~v_697 | ~v_2326 | ~v_2325 | ~v_2250 | ~v_2324 | ~v_2323 | ~v_2247 | ~v_468 | ~v_467 | ~v_2278 | ~v_2277 | ~v_2276 | ~v_2275 | ~v_696 | ~v_638 | ~v_695 | ~v_637 | ~v_1451 | ~v_1450 | ~v_1315 | ~v_1449 | ~v_1448 | ~v_1312 | ~v_1367 | ~v_1366 | ~v_1365 | ~v_1364 | ~v_2242 | ~v_2241 | ~v_2240 | ~v_2239 | v_2327;
assign x_21864 = v_2326 | v_139;
assign x_21865 = v_2326 | v_89;
assign x_21866 = v_2325 | v_140;
assign x_21867 = v_2325 | v_84;
assign x_21868 = v_2324 | ~v_139;
assign x_21869 = v_2324 | v_74;
assign x_21870 = v_2323 | ~v_140;
assign x_21871 = v_2323 | v_69;
assign x_21872 = v_18 | v_17 | v_16 | v_15 | v_14 | ~v_453 | ~v_452 | v_136 | v_135 | v_134 | v_163 | v_162 | v_161 | v_182 | ~v_693 | ~v_692 | ~v_2321 | ~v_2320 | ~v_2235 | ~v_2319 | ~v_2318 | ~v_2232 | ~v_2273 | ~v_2272 | ~v_2271 | ~v_2270 | ~v_691 | ~v_623 | ~v_690 | ~v_622 | ~v_1442 | ~v_1441 | ~v_1290 | ~v_1440 | ~v_1439 | ~v_1287 | ~v_1358 | ~v_1357 | ~v_1356 | ~v_1355 | ~v_2227 | ~v_2226 | ~v_2225 | ~v_2224 | v_2322;
assign x_21873 = v_2321 | v_139;
assign x_21874 = v_2321 | v_47;
assign x_21875 = v_2320 | v_140;
assign x_21876 = v_2320 | v_42;
assign x_21877 = v_2319 | ~v_139;
assign x_21878 = v_2319 | v_32;
assign x_21879 = v_2318 | ~v_140;
assign x_21880 = v_2318 | v_27;
assign x_21881 = v_2317 | ~v_2306;
assign x_21882 = v_2317 | ~v_2311;
assign x_21883 = v_2317 | ~v_2316;
assign x_21884 = v_103 | v_96 | v_100 | v_151 | v_171 | v_170 | v_169 | v_160 | v_150 | v_149 | v_147 | v_184 | ~v_655 | ~v_654 | ~v_2265 | ~v_2262 | ~v_2315 | ~v_2314 | ~v_2313 | ~v_2312 | ~v_297 | ~v_296 | ~v_2283 | ~v_2282 | ~v_2281 | ~v_2280 | ~v_653 | ~v_652 | ~v_651 | ~v_650 | ~v_1340 | ~v_1337 | ~v_1432 | ~v_1431 | ~v_1430 | ~v_1429 | ~v_1376 | ~v_1375 | ~v_1374 | ~v_1373 | ~v_2257 | ~v_2256 | ~v_2255 | ~v_2254 | v_2316;
assign x_21885 = v_2315 | v_176;
assign x_21886 = v_2315 | v_131;
assign x_21887 = v_2314 | v_175;
assign x_21888 = v_2314 | v_126;
assign x_21889 = v_2313 | ~v_176;
assign x_21890 = v_2313 | v_116;
assign x_21891 = v_2312 | ~v_175;
assign x_21892 = v_2312 | v_111;
assign x_21893 = v_54 | v_61 | v_58 | v_144 | v_159 | v_145 | v_142 | v_167 | v_166 | v_165 | v_146 | v_183 | ~v_640 | ~v_639 | ~v_2250 | ~v_2247 | ~v_2310 | ~v_2309 | ~v_2308 | ~v_2307 | ~v_264 | ~v_263 | ~v_2278 | ~v_2277 | ~v_2276 | ~v_2275 | ~v_638 | ~v_637 | ~v_636 | ~v_635 | ~v_1315 | ~v_1312 | ~v_1423 | ~v_1422 | ~v_1421 | ~v_1420 | ~v_1367 | ~v_1366 | ~v_1365 | ~v_1364 | ~v_2242 | ~v_2241 | ~v_2240 | ~v_2239 | v_2311;
assign x_21894 = v_2310 | v_176;
assign x_21895 = v_2310 | v_89;
assign x_21896 = v_2309 | v_175;
assign x_21897 = v_2309 | v_84;
assign x_21898 = v_2308 | ~v_176;
assign x_21899 = v_2308 | v_74;
assign x_21900 = v_2307 | ~v_175;
assign x_21901 = v_2307 | v_69;
assign x_21902 = v_18 | v_15 | v_11 | v_136 | v_134 | v_137 | v_138 | v_163 | v_162 | v_161 | v_155 | v_182 | ~v_625 | ~v_624 | ~v_2235 | ~v_2232 | ~v_2305 | ~v_2304 | ~v_2303 | ~v_2302 | ~v_231 | ~v_230 | ~v_2273 | ~v_2272 | ~v_2271 | ~v_2270 | ~v_623 | ~v_622 | ~v_621 | ~v_620 | ~v_1290 | ~v_1287 | ~v_1414 | ~v_1413 | ~v_1412 | ~v_1411 | ~v_1358 | ~v_1357 | ~v_1356 | ~v_1355 | ~v_2227 | ~v_2226 | ~v_2225 | ~v_2224 | v_2306;
assign x_21903 = v_2305 | v_176;
assign x_21904 = v_2305 | v_47;
assign x_21905 = v_2304 | v_175;
assign x_21906 = v_2304 | v_42;
assign x_21907 = v_2303 | ~v_176;
assign x_21908 = v_2303 | v_32;
assign x_21909 = v_2302 | ~v_175;
assign x_21910 = v_2302 | v_27;
assign x_21911 = v_2301 | ~v_2290;
assign x_21912 = v_2301 | ~v_2295;
assign x_21913 = v_2301 | ~v_2300;
assign x_21914 = v_101 | v_97 | v_100 | v_102 | v_172 | v_171 | v_170 | v_169 | v_150 | v_148 | v_147 | v_184 | ~v_671 | ~v_670 | ~v_2265 | ~v_2262 | ~v_2299 | ~v_2298 | ~v_2297 | ~v_2296 | ~v_387 | ~v_386 | ~v_2283 | ~v_2282 | ~v_2281 | ~v_2280 | ~v_653 | ~v_652 | ~v_669 | ~v_668 | ~v_1340 | ~v_1337 | ~v_1404 | ~v_1403 | ~v_1402 | ~v_1401 | ~v_1376 | ~v_1375 | ~v_1374 | ~v_1373 | ~v_2257 | ~v_2256 | ~v_2255 | ~v_2254 | v_2300;
assign x_21915 = v_2299 | v_141;
assign x_21916 = v_2299 | v_131;
assign x_21917 = v_2298 | v_141;
assign x_21918 = v_2298 | v_126;
assign x_21919 = v_2297 | ~v_141;
assign x_21920 = v_2297 | v_116;
assign x_21921 = v_2296 | ~v_141;
assign x_21922 = v_2296 | v_111;
assign x_21923 = v_55 | v_60 | v_59 | v_58 | v_145 | v_143 | v_142 | v_168 | v_167 | v_166 | v_165 | v_183 | ~v_666 | ~v_665 | ~v_2250 | ~v_2247 | ~v_2294 | ~v_2293 | ~v_2292 | ~v_2291 | ~v_372 | ~v_371 | ~v_2278 | ~v_2277 | ~v_2276 | ~v_2275 | ~v_638 | ~v_637 | ~v_664 | ~v_663 | ~v_1315 | ~v_1312 | ~v_1395 | ~v_1394 | ~v_1393 | ~v_1392 | ~v_1367 | ~v_1366 | ~v_1365 | ~v_1364 | ~v_2242 | ~v_2241 | ~v_2240 | ~v_2239 | v_2295;
assign x_21924 = v_2294 | v_141;
assign x_21925 = v_2294 | v_89;
assign x_21926 = v_2293 | v_141;
assign x_21927 = v_2293 | v_84;
assign x_21928 = v_2292 | ~v_141;
assign x_21929 = v_2292 | v_74;
assign x_21930 = v_2291 | ~v_141;
assign x_21931 = v_2291 | v_69;
assign x_21932 = v_17 | v_16 | v_15 | v_12 | v_135 | v_134 | v_137 | v_164 | v_163 | v_162 | v_161 | v_182 | ~v_661 | ~v_660 | ~v_2235 | ~v_2232 | ~v_2289 | ~v_2288 | ~v_2287 | ~v_2286 | ~v_357 | ~v_356 | ~v_2273 | ~v_2272 | ~v_2271 | ~v_2270 | ~v_623 | ~v_622 | ~v_659 | ~v_658 | ~v_1290 | ~v_1287 | ~v_1386 | ~v_1385 | ~v_1384 | ~v_1383 | ~v_1358 | ~v_1357 | ~v_1356 | ~v_1355 | ~v_2227 | ~v_2226 | ~v_2225 | ~v_2224 | v_2290;
assign x_21933 = v_2289 | v_141;
assign x_21934 = v_2289 | v_47;
assign x_21935 = v_2288 | v_141;
assign x_21936 = v_2288 | v_42;
assign x_21937 = v_2287 | ~v_141;
assign x_21938 = v_2287 | v_32;
assign x_21939 = v_2286 | ~v_141;
assign x_21940 = v_2286 | v_27;
assign x_21941 = v_2285 | ~v_2274;
assign x_21942 = v_2285 | ~v_2279;
assign x_21943 = v_2285 | ~v_2284;
assign x_21944 = v_103 | v_101 | v_100 | v_95 | v_102 | v_171 | v_170 | v_169 | v_150 | v_149 | v_148 | v_184 | ~v_2265 | ~v_2262 | ~v_2261 | ~v_2260 | ~v_2259 | ~v_2258 | ~v_435 | ~v_434 | ~v_2283 | ~v_2282 | ~v_2281 | ~v_2280 | ~v_653 | ~v_652 | ~v_687 | ~v_686 | ~v_685 | ~v_684 | ~v_1340 | ~v_1337 | ~v_1336 | ~v_1335 | ~v_1334 | ~v_1333 | ~v_1376 | ~v_1375 | ~v_1374 | ~v_1373 | ~v_2257 | ~v_2256 | ~v_2255 | ~v_2254 | v_2284;
assign x_21945 = v_2283 | v_174;
assign x_21946 = v_2283 | v_128;
assign x_21947 = v_2282 | v_173;
assign x_21948 = v_2282 | v_125;
assign x_21949 = v_2281 | ~v_174;
assign x_21950 = v_2281 | v_113;
assign x_21951 = v_2280 | ~v_173;
assign x_21952 = v_2280 | v_110;
assign x_21953 = v_53 | v_61 | v_60 | v_59 | v_58 | v_144 | v_145 | v_143 | v_167 | v_166 | v_165 | v_183 | ~v_2250 | ~v_2247 | ~v_2246 | ~v_2245 | ~v_2244 | ~v_2243 | ~v_420 | ~v_419 | ~v_2278 | ~v_2277 | ~v_2276 | ~v_2275 | ~v_638 | ~v_637 | ~v_682 | ~v_681 | ~v_680 | ~v_679 | ~v_1315 | ~v_1312 | ~v_1311 | ~v_1310 | ~v_1309 | ~v_1308 | ~v_1367 | ~v_1366 | ~v_1365 | ~v_1364 | ~v_2242 | ~v_2241 | ~v_2240 | ~v_2239 | v_2279;
assign x_21954 = v_2278 | v_174;
assign x_21955 = v_2278 | v_86;
assign x_21956 = v_2277 | v_173;
assign x_21957 = v_2277 | v_83;
assign x_21958 = v_2276 | ~v_174;
assign x_21959 = v_2276 | v_71;
assign x_21960 = v_2275 | ~v_173;
assign x_21961 = v_2275 | v_68;
assign x_21962 = v_18 | v_17 | v_16 | v_15 | v_10 | v_136 | v_135 | v_137 | v_163 | v_162 | v_161 | v_182 | ~v_2235 | ~v_2232 | ~v_2231 | ~v_2230 | ~v_2229 | ~v_2228 | ~v_405 | ~v_404 | ~v_2273 | ~v_2272 | ~v_2271 | ~v_2270 | ~v_623 | ~v_622 | ~v_677 | ~v_676 | ~v_675 | ~v_674 | ~v_1290 | ~v_1287 | ~v_1286 | ~v_1285 | ~v_1284 | ~v_1283 | ~v_1358 | ~v_1357 | ~v_1356 | ~v_1355 | ~v_2227 | ~v_2226 | ~v_2225 | ~v_2224 | v_2274;
assign x_21963 = v_2273 | v_174;
assign x_21964 = v_2273 | v_44;
assign x_21965 = v_2272 | v_173;
assign x_21966 = v_2272 | v_41;
assign x_21967 = v_2271 | ~v_174;
assign x_21968 = v_2271 | v_29;
assign x_21969 = v_2270 | ~v_173;
assign x_21970 = v_2270 | v_26;
assign x_21971 = v_2269 | ~v_2238;
assign x_21972 = v_2269 | ~v_2253;
assign x_21973 = v_2269 | ~v_2268;
assign x_21974 = v_98 | v_103 | v_101 | v_100 | v_102 | v_170 | v_169 | v_150 | v_149 | v_148 | v_147 | v_184 | ~v_609 | ~v_608 | ~v_2267 | ~v_2266 | ~v_2265 | ~v_2264 | ~v_2263 | ~v_2262 | ~v_299 | ~v_298 | ~v_2261 | ~v_2260 | ~v_2259 | ~v_2258 | ~v_435 | ~v_434 | ~v_607 | ~v_606 | ~v_1342 | ~v_1341 | ~v_1340 | ~v_1339 | ~v_1338 | ~v_1337 | ~v_1336 | ~v_1335 | ~v_1334 | ~v_1333 | ~v_2257 | ~v_2256 | ~v_2255 | ~v_2254 | v_2268;
assign x_21975 = v_2267 | v_139;
assign x_21976 = v_2267 | v_128;
assign x_21977 = v_2266 | v_140;
assign x_21978 = v_2266 | v_125;
assign x_21979 = v_2265 | v_141;
assign x_21980 = v_2265 | v_124;
assign x_21981 = v_2264 | ~v_139;
assign x_21982 = v_2264 | v_113;
assign x_21983 = v_2263 | ~v_140;
assign x_21984 = v_2263 | v_110;
assign x_21985 = v_2262 | ~v_141;
assign x_21986 = v_2262 | v_109;
assign x_21987 = v_2261 | v_174;
assign x_21988 = v_2261 | v_131;
assign x_21989 = v_2260 | v_173;
assign x_21990 = v_2260 | v_126;
assign x_21991 = v_2259 | ~v_174;
assign x_21992 = v_2259 | v_116;
assign x_21993 = v_2258 | ~v_173;
assign x_21994 = v_2258 | v_111;
assign x_21995 = v_2257 | v_175;
assign x_21996 = v_2257 | v_123;
assign x_21997 = v_2256 | v_176;
assign x_21998 = v_2256 | v_120;
assign x_21999 = v_2255 | ~v_175;
assign x_22000 = v_2255 | v_108;
assign x_22001 = v_2254 | ~v_176;
assign x_22002 = v_2254 | v_105;
assign x_22003 = v_56 | v_61 | v_60 | v_59 | v_58 | v_144 | v_145 | v_143 | v_142 | v_166 | v_165 | v_183 | ~v_604 | ~v_603 | ~v_266 | ~v_2252 | ~v_2251 | ~v_2250 | ~v_2249 | ~v_2248 | ~v_2247 | ~v_265 | ~v_2246 | ~v_2245 | ~v_2244 | ~v_2243 | ~v_420 | ~v_419 | ~v_602 | ~v_601 | ~v_1317 | ~v_1316 | ~v_1315 | ~v_1314 | ~v_1313 | ~v_1312 | ~v_1311 | ~v_1310 | ~v_1309 | ~v_1308 | ~v_2242 | ~v_2241 | ~v_2240 | ~v_2239 | v_2253;
assign x_22004 = v_2252 | v_139;
assign x_22005 = v_2252 | v_86;
assign x_22006 = v_2251 | v_140;
assign x_22007 = v_2251 | v_83;
assign x_22008 = v_2250 | v_141;
assign x_22009 = v_2250 | v_82;
assign x_22010 = v_2249 | ~v_139;
assign x_22011 = v_2249 | v_71;
assign x_22012 = v_2248 | ~v_140;
assign x_22013 = v_2248 | v_68;
assign x_22014 = v_2247 | ~v_141;
assign x_22015 = v_2247 | v_67;
assign x_22016 = v_2246 | v_174;
assign x_22017 = v_2246 | v_89;
assign x_22018 = v_2245 | v_173;
assign x_22019 = v_2245 | v_84;
assign x_22020 = v_2244 | ~v_174;
assign x_22021 = v_2244 | v_74;
assign x_22022 = v_2243 | ~v_173;
assign x_22023 = v_2243 | v_69;
assign x_22024 = v_2242 | v_175;
assign x_22025 = v_2242 | v_81;
assign x_22026 = v_2241 | v_176;
assign x_22027 = v_2241 | v_78;
assign x_22028 = v_2240 | ~v_175;
assign x_22029 = v_2240 | v_66;
assign x_22030 = v_2239 | ~v_176;
assign x_22031 = v_2239 | v_63;
assign x_22032 = v_13 | v_18 | v_17 | v_16 | v_15 | v_136 | v_135 | v_134 | v_137 | v_162 | v_161 | v_182 | ~v_599 | ~v_598 | ~v_2237 | ~v_2236 | ~v_2235 | ~v_2234 | ~v_2233 | ~v_2232 | ~v_233 | ~v_232 | ~v_2231 | ~v_2230 | ~v_2229 | ~v_2228 | ~v_405 | ~v_404 | ~v_597 | ~v_596 | ~v_1292 | ~v_1291 | ~v_1290 | ~v_1289 | ~v_1288 | ~v_1287 | ~v_1286 | ~v_1285 | ~v_1284 | ~v_1283 | ~v_2227 | ~v_2226 | ~v_2225 | ~v_2224 | v_2238;
assign x_22033 = v_2237 | v_139;
assign x_22034 = v_2237 | v_44;
assign x_22035 = v_2236 | v_140;
assign x_22036 = v_2236 | v_41;
assign x_22037 = v_2235 | v_141;
assign x_22038 = v_2235 | v_40;
assign x_22039 = v_2234 | ~v_139;
assign x_22040 = v_2234 | v_29;
assign x_22041 = v_2233 | ~v_140;
assign x_22042 = v_2233 | v_26;
assign x_22043 = v_2232 | ~v_141;
assign x_22044 = v_2232 | v_25;
assign x_22045 = v_2231 | v_174;
assign x_22046 = v_2231 | v_47;
assign x_22047 = v_2230 | v_173;
assign x_22048 = v_2230 | v_42;
assign x_22049 = v_2229 | ~v_174;
assign x_22050 = v_2229 | v_32;
assign x_22051 = v_2228 | ~v_173;
assign x_22052 = v_2228 | v_27;
assign x_22053 = v_2227 | v_175;
assign x_22054 = v_2227 | v_39;
assign x_22055 = v_2226 | v_176;
assign x_22056 = v_2226 | v_36;
assign x_22057 = v_2225 | ~v_175;
assign x_22058 = v_2225 | v_24;
assign x_22059 = v_2224 | ~v_176;
assign x_22060 = v_2224 | v_21;
assign x_22061 = v_2223 | ~v_2218;
assign x_22062 = v_2223 | ~v_2222;
assign x_22063 = v_2223 | ~v_187;
assign x_22064 = v_2223 | ~v_190;
assign x_22065 = v_2223 | ~v_176;
assign x_22066 = v_2223 | ~v_175;
assign x_22067 = ~v_185 | ~v_2221 | v_2222;
assign x_22068 = v_2221 | ~v_2219;
assign x_22069 = v_2221 | ~v_2220;
assign x_22070 = v_2221 | ~v_140;
assign x_22071 = v_2221 | ~v_139;
assign x_22072 = ~v_189 | ~v_193 | v_2220;
assign x_22073 = ~v_185 | ~v_195 | v_2219;
assign x_22074 = ~v_188 | ~v_1272 | v_2218;
assign x_22075 = v_2217 | ~v_2033;
assign x_22076 = v_2217 | ~v_2216;
assign x_22077 = v_176 | v_175 | ~v_2215 | ~v_732 | ~v_729 | ~v_2036 | ~v_2035 | v_2216;
assign x_22078 = v_2215 | ~v_2082;
assign x_22079 = v_2215 | ~v_2098;
assign x_22080 = v_2215 | ~v_2114;
assign x_22081 = v_2215 | ~v_2130;
assign x_22082 = v_2215 | ~v_2146;
assign x_22083 = v_2215 | ~v_2150;
assign x_22084 = v_2215 | ~v_2166;
assign x_22085 = v_2215 | ~v_2170;
assign x_22086 = v_2215 | ~v_2174;
assign x_22087 = v_2215 | ~v_2178;
assign x_22088 = v_2215 | ~v_2182;
assign x_22089 = v_2215 | ~v_2198;
assign x_22090 = v_2215 | ~v_2202;
assign x_22091 = v_2215 | ~v_2206;
assign x_22092 = v_2215 | ~v_2210;
assign x_22093 = v_2215 | ~v_2214;
assign x_22094 = v_2215 | ~v_1263;
assign x_22095 = v_2215 | ~v_1264;
assign x_22096 = v_2215 | ~v_1265;
assign x_22097 = v_2215 | ~v_1266;
assign x_22098 = ~v_2213 | ~v_2212 | ~v_2211 | v_2214;
assign x_22099 = v_2213 | ~v_2067;
assign x_22100 = v_2213 | ~v_2068;
assign x_22101 = v_2213 | ~v_2069;
assign x_22102 = v_2213 | ~v_2070;
assign x_22103 = v_2213 | ~v_817;
assign x_22104 = v_2213 | ~v_818;
assign x_22105 = v_2213 | ~v_1011;
assign x_22106 = v_2213 | ~v_819;
assign x_22107 = v_2213 | ~v_1012;
assign x_22108 = v_2213 | ~v_820;
assign x_22109 = v_2213 | ~v_821;
assign x_22110 = v_2213 | ~v_1013;
assign x_22111 = v_2213 | ~v_822;
assign x_22112 = v_2213 | ~v_1014;
assign x_22113 = v_2213 | ~v_2075;
assign x_22114 = v_2213 | ~v_2076;
assign x_22115 = v_2213 | ~v_2141;
assign x_22116 = v_2213 | ~v_2077;
assign x_22117 = v_2213 | ~v_2142;
assign x_22118 = v_2213 | ~v_2078;
assign x_22119 = v_2213 | ~v_2079;
assign x_22120 = v_2213 | ~v_2143;
assign x_22121 = v_2213 | ~v_2080;
assign x_22122 = v_2213 | ~v_2144;
assign x_22123 = v_2213 | ~v_839;
assign x_22124 = v_2213 | ~v_1257;
assign x_22125 = v_2213 | ~v_1023;
assign x_22126 = v_2213 | ~v_840;
assign x_22127 = v_2213 | ~v_1258;
assign x_22128 = v_2213 | ~v_1024;
assign x_22129 = v_2213 | ~v_184;
assign x_22130 = v_2213 | ~v_170;
assign x_22131 = v_2213 | ~v_169;
assign x_22132 = v_2213 | ~v_149;
assign x_22133 = v_2213 | ~v_148;
assign x_22134 = v_2213 | ~v_1259;
assign x_22135 = v_2213 | ~v_1260;
assign x_22136 = v_2213 | ~v_103;
assign x_22137 = v_2213 | ~v_102;
assign x_22138 = v_2213 | ~v_101;
assign x_22139 = v_2213 | ~v_100;
assign x_22140 = v_2213 | ~v_99;
assign x_22141 = v_2213 | ~v_98;
assign x_22142 = v_2213 | ~v_95;
assign x_22143 = v_2212 | ~v_2052;
assign x_22144 = v_2212 | ~v_2053;
assign x_22145 = v_2212 | ~v_2054;
assign x_22146 = v_2212 | ~v_2055;
assign x_22147 = v_2212 | ~v_784;
assign x_22148 = v_2212 | ~v_785;
assign x_22149 = v_2212 | ~v_996;
assign x_22150 = v_2212 | ~v_786;
assign x_22151 = v_2212 | ~v_997;
assign x_22152 = v_2212 | ~v_787;
assign x_22153 = v_2212 | ~v_788;
assign x_22154 = v_2212 | ~v_998;
assign x_22155 = v_2212 | ~v_789;
assign x_22156 = v_2212 | ~v_999;
assign x_22157 = v_2212 | ~v_2060;
assign x_22158 = v_2212 | ~v_2061;
assign x_22159 = v_2212 | ~v_2136;
assign x_22160 = v_2212 | ~v_2062;
assign x_22161 = v_2212 | ~v_2137;
assign x_22162 = v_2212 | ~v_2063;
assign x_22163 = v_2212 | ~v_2064;
assign x_22164 = v_2212 | ~v_2138;
assign x_22165 = v_2212 | ~v_2065;
assign x_22166 = v_2212 | ~v_2139;
assign x_22167 = v_2212 | ~v_806;
assign x_22168 = v_2212 | ~v_1252;
assign x_22169 = v_2212 | ~v_1008;
assign x_22170 = v_2212 | ~v_1253;
assign x_22171 = v_2212 | ~v_1009;
assign x_22172 = v_2212 | ~v_807;
assign x_22173 = v_2212 | ~v_183;
assign x_22174 = v_2212 | ~v_166;
assign x_22175 = v_2212 | ~v_165;
assign x_22176 = v_2212 | ~v_144;
assign x_22177 = v_2212 | ~v_143;
assign x_22178 = v_2212 | ~v_1254;
assign x_22179 = v_2212 | ~v_1255;
assign x_22180 = v_2212 | ~v_61;
assign x_22181 = v_2212 | ~v_60;
assign x_22182 = v_2212 | ~v_59;
assign x_22183 = v_2212 | ~v_58;
assign x_22184 = v_2212 | ~v_57;
assign x_22185 = v_2212 | ~v_56;
assign x_22186 = v_2212 | ~v_53;
assign x_22187 = v_2211 | ~v_2037;
assign x_22188 = v_2211 | ~v_2038;
assign x_22189 = v_2211 | ~v_2039;
assign x_22190 = v_2211 | ~v_2040;
assign x_22191 = v_2211 | ~v_751;
assign x_22192 = v_2211 | ~v_752;
assign x_22193 = v_2211 | ~v_981;
assign x_22194 = v_2211 | ~v_753;
assign x_22195 = v_2211 | ~v_982;
assign x_22196 = v_2211 | ~v_754;
assign x_22197 = v_2211 | ~v_755;
assign x_22198 = v_2211 | ~v_983;
assign x_22199 = v_2211 | ~v_756;
assign x_22200 = v_2211 | ~v_984;
assign x_22201 = v_2211 | ~v_2045;
assign x_22202 = v_2211 | ~v_2046;
assign x_22203 = v_2211 | ~v_2131;
assign x_22204 = v_2211 | ~v_2047;
assign x_22205 = v_2211 | ~v_2132;
assign x_22206 = v_2211 | ~v_2048;
assign x_22207 = v_2211 | ~v_2049;
assign x_22208 = v_2211 | ~v_2133;
assign x_22209 = v_2211 | ~v_2050;
assign x_22210 = v_2211 | ~v_2134;
assign x_22211 = v_2211 | ~v_773;
assign x_22212 = v_2211 | ~v_774;
assign x_22213 = v_2211 | ~v_182;
assign x_22214 = v_2211 | ~v_162;
assign x_22215 = v_2211 | ~v_161;
assign x_22216 = v_2211 | ~v_1247;
assign x_22217 = v_2211 | ~v_1248;
assign x_22218 = v_2211 | ~v_136;
assign x_22219 = v_2211 | ~v_135;
assign x_22220 = v_2211 | ~v_1249;
assign x_22221 = v_2211 | ~v_993;
assign x_22222 = v_2211 | ~v_1250;
assign x_22223 = v_2211 | ~v_994;
assign x_22224 = v_2211 | ~v_18;
assign x_22225 = v_2211 | ~v_17;
assign x_22226 = v_2211 | ~v_16;
assign x_22227 = v_2211 | ~v_15;
assign x_22228 = v_2211 | ~v_14;
assign x_22229 = v_2211 | ~v_13;
assign x_22230 = v_2211 | ~v_10;
assign x_22231 = ~v_2209 | ~v_2208 | ~v_2207 | v_2210;
assign x_22232 = v_2209 | ~v_2067;
assign x_22233 = v_2209 | ~v_2068;
assign x_22234 = v_2209 | ~v_2069;
assign x_22235 = v_2209 | ~v_2070;
assign x_22236 = v_2209 | ~v_1073;
assign x_22237 = v_2209 | ~v_1074;
assign x_22238 = v_2209 | ~v_1075;
assign x_22239 = v_2209 | ~v_1076;
assign x_22240 = v_2209 | ~v_817;
assign x_22241 = v_2209 | ~v_1011;
assign x_22242 = v_2209 | ~v_1012;
assign x_22243 = v_2209 | ~v_820;
assign x_22244 = v_2209 | ~v_1013;
assign x_22245 = v_2209 | ~v_1014;
assign x_22246 = v_2209 | ~v_2193;
assign x_22247 = v_2209 | ~v_2194;
assign x_22248 = v_2209 | ~v_2195;
assign x_22249 = v_2209 | ~v_2196;
assign x_22250 = v_2209 | ~v_2075;
assign x_22251 = v_2209 | ~v_2141;
assign x_22252 = v_2209 | ~v_2142;
assign x_22253 = v_2209 | ~v_2078;
assign x_22254 = v_2209 | ~v_2143;
assign x_22255 = v_2209 | ~v_2144;
assign x_22256 = v_2209 | ~v_1085;
assign x_22257 = v_2209 | ~v_1131;
assign x_22258 = v_2209 | ~v_1132;
assign x_22259 = v_2209 | ~v_1086;
assign x_22260 = v_2209 | ~v_1133;
assign x_22261 = v_2209 | ~v_1134;
assign x_22262 = v_2209 | ~v_1023;
assign x_22263 = v_2209 | ~v_1024;
assign x_22264 = v_2209 | ~v_184;
assign x_22265 = v_2209 | ~v_172;
assign x_22266 = v_2209 | ~v_171;
assign x_22267 = v_2209 | ~v_170;
assign x_22268 = v_2209 | ~v_149;
assign x_22269 = v_2209 | ~v_148;
assign x_22270 = v_2209 | ~v_147;
assign x_22271 = v_2209 | ~v_102;
assign x_22272 = v_2209 | ~v_101;
assign x_22273 = v_2209 | ~v_100;
assign x_22274 = v_2209 | ~v_99;
assign x_22275 = v_2209 | ~v_93;
assign x_22276 = v_2208 | ~v_2052;
assign x_22277 = v_2208 | ~v_2053;
assign x_22278 = v_2208 | ~v_2054;
assign x_22279 = v_2208 | ~v_2055;
assign x_22280 = v_2208 | ~v_1058;
assign x_22281 = v_2208 | ~v_1059;
assign x_22282 = v_2208 | ~v_1060;
assign x_22283 = v_2208 | ~v_1061;
assign x_22284 = v_2208 | ~v_784;
assign x_22285 = v_2208 | ~v_996;
assign x_22286 = v_2208 | ~v_997;
assign x_22287 = v_2208 | ~v_787;
assign x_22288 = v_2208 | ~v_998;
assign x_22289 = v_2208 | ~v_999;
assign x_22290 = v_2208 | ~v_2188;
assign x_22291 = v_2208 | ~v_2189;
assign x_22292 = v_2208 | ~v_2190;
assign x_22293 = v_2208 | ~v_2191;
assign x_22294 = v_2208 | ~v_2060;
assign x_22295 = v_2208 | ~v_2136;
assign x_22296 = v_2208 | ~v_2137;
assign x_22297 = v_2208 | ~v_2063;
assign x_22298 = v_2208 | ~v_2138;
assign x_22299 = v_2208 | ~v_2139;
assign x_22300 = v_2208 | ~v_1070;
assign x_22301 = v_2208 | ~v_1126;
assign x_22302 = v_2208 | ~v_1127;
assign x_22303 = v_2208 | ~v_1071;
assign x_22304 = v_2208 | ~v_1128;
assign x_22305 = v_2208 | ~v_1129;
assign x_22306 = v_2208 | ~v_1008;
assign x_22307 = v_2208 | ~v_1009;
assign x_22308 = v_2208 | ~v_183;
assign x_22309 = v_2208 | ~v_168;
assign x_22310 = v_2208 | ~v_167;
assign x_22311 = v_2208 | ~v_166;
assign x_22312 = v_2208 | ~v_144;
assign x_22313 = v_2208 | ~v_143;
assign x_22314 = v_2208 | ~v_142;
assign x_22315 = v_2208 | ~v_60;
assign x_22316 = v_2208 | ~v_59;
assign x_22317 = v_2208 | ~v_58;
assign x_22318 = v_2208 | ~v_57;
assign x_22319 = v_2208 | ~v_51;
assign x_22320 = v_2207 | ~v_2037;
assign x_22321 = v_2207 | ~v_2038;
assign x_22322 = v_2207 | ~v_2039;
assign x_22323 = v_2207 | ~v_2040;
assign x_22324 = v_2207 | ~v_1043;
assign x_22325 = v_2207 | ~v_1044;
assign x_22326 = v_2207 | ~v_1045;
assign x_22327 = v_2207 | ~v_1046;
assign x_22328 = v_2207 | ~v_751;
assign x_22329 = v_2207 | ~v_981;
assign x_22330 = v_2207 | ~v_982;
assign x_22331 = v_2207 | ~v_754;
assign x_22332 = v_2207 | ~v_983;
assign x_22333 = v_2207 | ~v_984;
assign x_22334 = v_2207 | ~v_2183;
assign x_22335 = v_2207 | ~v_2184;
assign x_22336 = v_2207 | ~v_2185;
assign x_22337 = v_2207 | ~v_2186;
assign x_22338 = v_2207 | ~v_2045;
assign x_22339 = v_2207 | ~v_2131;
assign x_22340 = v_2207 | ~v_2132;
assign x_22341 = v_2207 | ~v_2048;
assign x_22342 = v_2207 | ~v_2133;
assign x_22343 = v_2207 | ~v_2134;
assign x_22344 = v_2207 | ~v_1055;
assign x_22345 = v_2207 | ~v_1121;
assign x_22346 = v_2207 | ~v_1122;
assign x_22347 = v_2207 | ~v_1056;
assign x_22348 = v_2207 | ~v_1123;
assign x_22349 = v_2207 | ~v_1124;
assign x_22350 = v_2207 | ~v_182;
assign x_22351 = v_2207 | ~v_164;
assign x_22352 = v_2207 | ~v_163;
assign x_22353 = v_2207 | ~v_162;
assign x_22354 = v_2207 | ~v_136;
assign x_22355 = v_2207 | ~v_135;
assign x_22356 = v_2207 | ~v_134;
assign x_22357 = v_2207 | ~v_993;
assign x_22358 = v_2207 | ~v_994;
assign x_22359 = v_2207 | ~v_17;
assign x_22360 = v_2207 | ~v_16;
assign x_22361 = v_2207 | ~v_15;
assign x_22362 = v_2207 | ~v_14;
assign x_22363 = v_2207 | ~v_8;
assign x_22364 = ~v_2205 | ~v_2204 | ~v_2203 | v_2206;
assign x_22365 = v_2205 | ~v_2067;
assign x_22366 = v_2205 | ~v_2068;
assign x_22367 = v_2205 | ~v_2069;
assign x_22368 = v_2205 | ~v_2070;
assign x_22369 = v_2205 | ~v_1073;
assign x_22370 = v_2205 | ~v_1074;
assign x_22371 = v_2205 | ~v_1075;
assign x_22372 = v_2205 | ~v_1076;
assign x_22373 = v_2205 | ~v_919;
assign x_22374 = v_2205 | ~v_920;
assign x_22375 = v_2205 | ~v_817;
assign x_22376 = v_2205 | ~v_820;
assign x_22377 = v_2205 | ~v_2125;
assign x_22378 = v_2205 | ~v_2126;
assign x_22379 = v_2205 | ~v_2127;
assign x_22380 = v_2205 | ~v_2128;
assign x_22381 = v_2205 | ~v_2193;
assign x_22382 = v_2205 | ~v_2194;
assign x_22383 = v_2205 | ~v_2195;
assign x_22384 = v_2205 | ~v_2196;
assign x_22385 = v_2205 | ~v_2075;
assign x_22386 = v_2205 | ~v_2078;
assign x_22387 = v_2205 | ~v_927;
assign x_22388 = v_2205 | ~v_928;
assign x_22389 = v_2205 | ~v_1099;
assign x_22390 = v_2205 | ~v_1100;
assign x_22391 = v_2205 | ~v_1101;
assign x_22392 = v_2205 | ~v_1102;
assign x_22393 = v_2205 | ~v_1085;
assign x_22394 = v_2205 | ~v_1086;
assign x_22395 = v_2205 | ~v_931;
assign x_22396 = v_2205 | ~v_932;
assign x_22397 = v_2205 | ~v_184;
assign x_22398 = v_2205 | ~v_171;
assign x_22399 = v_2205 | ~v_170;
assign x_22400 = v_2205 | ~v_150;
assign x_22401 = v_2205 | ~v_149;
assign x_22402 = v_2205 | ~v_103;
assign x_22403 = v_2205 | ~v_102;
assign x_22404 = v_2205 | ~v_101;
assign x_22405 = v_2205 | ~v_100;
assign x_22406 = v_2205 | ~v_96;
assign x_22407 = v_2205 | ~v_95;
assign x_22408 = v_2205 | ~v_93;
assign x_22409 = v_2204 | ~v_2052;
assign x_22410 = v_2204 | ~v_2053;
assign x_22411 = v_2204 | ~v_2054;
assign x_22412 = v_2204 | ~v_2055;
assign x_22413 = v_2204 | ~v_1058;
assign x_22414 = v_2204 | ~v_1059;
assign x_22415 = v_2204 | ~v_1060;
assign x_22416 = v_2204 | ~v_1061;
assign x_22417 = v_2204 | ~v_904;
assign x_22418 = v_2204 | ~v_905;
assign x_22419 = v_2204 | ~v_784;
assign x_22420 = v_2204 | ~v_787;
assign x_22421 = v_2204 | ~v_2120;
assign x_22422 = v_2204 | ~v_2121;
assign x_22423 = v_2204 | ~v_2122;
assign x_22424 = v_2204 | ~v_2123;
assign x_22425 = v_2204 | ~v_2188;
assign x_22426 = v_2204 | ~v_2189;
assign x_22427 = v_2204 | ~v_2190;
assign x_22428 = v_2204 | ~v_2191;
assign x_22429 = v_2204 | ~v_2060;
assign x_22430 = v_2204 | ~v_2063;
assign x_22431 = v_2204 | ~v_912;
assign x_22432 = v_2204 | ~v_913;
assign x_22433 = v_2204 | ~v_1094;
assign x_22434 = v_2204 | ~v_1095;
assign x_22435 = v_2204 | ~v_1096;
assign x_22436 = v_2204 | ~v_1097;
assign x_22437 = v_2204 | ~v_1070;
assign x_22438 = v_2204 | ~v_1071;
assign x_22439 = v_2204 | ~v_916;
assign x_22440 = v_2204 | ~v_917;
assign x_22441 = v_2204 | ~v_183;
assign x_22442 = v_2204 | ~v_167;
assign x_22443 = v_2204 | ~v_166;
assign x_22444 = v_2204 | ~v_145;
assign x_22445 = v_2204 | ~v_144;
assign x_22446 = v_2204 | ~v_61;
assign x_22447 = v_2204 | ~v_60;
assign x_22448 = v_2204 | ~v_59;
assign x_22449 = v_2204 | ~v_58;
assign x_22450 = v_2204 | ~v_54;
assign x_22451 = v_2204 | ~v_53;
assign x_22452 = v_2204 | ~v_51;
assign x_22453 = v_2203 | ~v_2037;
assign x_22454 = v_2203 | ~v_2038;
assign x_22455 = v_2203 | ~v_2039;
assign x_22456 = v_2203 | ~v_2040;
assign x_22457 = v_2203 | ~v_1043;
assign x_22458 = v_2203 | ~v_1044;
assign x_22459 = v_2203 | ~v_1045;
assign x_22460 = v_2203 | ~v_1046;
assign x_22461 = v_2203 | ~v_889;
assign x_22462 = v_2203 | ~v_890;
assign x_22463 = v_2203 | ~v_751;
assign x_22464 = v_2203 | ~v_754;
assign x_22465 = v_2203 | ~v_2115;
assign x_22466 = v_2203 | ~v_2116;
assign x_22467 = v_2203 | ~v_2117;
assign x_22468 = v_2203 | ~v_2118;
assign x_22469 = v_2203 | ~v_2183;
assign x_22470 = v_2203 | ~v_2184;
assign x_22471 = v_2203 | ~v_2185;
assign x_22472 = v_2203 | ~v_2186;
assign x_22473 = v_2203 | ~v_2045;
assign x_22474 = v_2203 | ~v_2048;
assign x_22475 = v_2203 | ~v_897;
assign x_22476 = v_2203 | ~v_898;
assign x_22477 = v_2203 | ~v_1089;
assign x_22478 = v_2203 | ~v_1090;
assign x_22479 = v_2203 | ~v_1091;
assign x_22480 = v_2203 | ~v_1092;
assign x_22481 = v_2203 | ~v_1055;
assign x_22482 = v_2203 | ~v_1056;
assign x_22483 = v_2203 | ~v_901;
assign x_22484 = v_2203 | ~v_902;
assign x_22485 = v_2203 | ~v_182;
assign x_22486 = v_2203 | ~v_163;
assign x_22487 = v_2203 | ~v_162;
assign x_22488 = v_2203 | ~v_137;
assign x_22489 = v_2203 | ~v_136;
assign x_22490 = v_2203 | ~v_18;
assign x_22491 = v_2203 | ~v_17;
assign x_22492 = v_2203 | ~v_16;
assign x_22493 = v_2203 | ~v_15;
assign x_22494 = v_2203 | ~v_11;
assign x_22495 = v_2203 | ~v_10;
assign x_22496 = v_2203 | ~v_8;
assign x_22497 = ~v_2201 | ~v_2200 | ~v_2199 | v_2202;
assign x_22498 = v_2201 | ~v_2067;
assign x_22499 = v_2201 | ~v_2068;
assign x_22500 = v_2201 | ~v_2069;
assign x_22501 = v_2201 | ~v_2070;
assign x_22502 = v_2201 | ~v_1073;
assign x_22503 = v_2201 | ~v_1074;
assign x_22504 = v_2201 | ~v_1075;
assign x_22505 = v_2201 | ~v_1076;
assign x_22506 = v_2201 | ~v_965;
assign x_22507 = v_2201 | ~v_966;
assign x_22508 = v_2201 | ~v_967;
assign x_22509 = v_2201 | ~v_968;
assign x_22510 = v_2201 | ~v_817;
assign x_22511 = v_2201 | ~v_820;
assign x_22512 = v_2201 | ~v_2109;
assign x_22513 = v_2201 | ~v_2110;
assign x_22514 = v_2201 | ~v_2111;
assign x_22515 = v_2201 | ~v_2112;
assign x_22516 = v_2201 | ~v_2193;
assign x_22517 = v_2201 | ~v_2194;
assign x_22518 = v_2201 | ~v_2195;
assign x_22519 = v_2201 | ~v_2196;
assign x_22520 = v_2201 | ~v_2075;
assign x_22521 = v_2201 | ~v_2078;
assign x_22522 = v_2201 | ~v_975;
assign x_22523 = v_2201 | ~v_976;
assign x_22524 = v_2201 | ~v_1115;
assign x_22525 = v_2201 | ~v_1116;
assign x_22526 = v_2201 | ~v_1085;
assign x_22527 = v_2201 | ~v_1086;
assign x_22528 = v_2201 | ~v_1117;
assign x_22529 = v_2201 | ~v_1118;
assign x_22530 = v_2201 | ~v_184;
assign x_22531 = v_2201 | ~v_171;
assign x_22532 = v_2201 | ~v_170;
assign x_22533 = v_2201 | ~v_151;
assign x_22534 = v_2201 | ~v_150;
assign x_22535 = v_2201 | ~v_149;
assign x_22536 = v_2201 | ~v_148;
assign x_22537 = v_2201 | ~v_147;
assign x_22538 = v_2201 | ~v_103;
assign x_22539 = v_2201 | ~v_101;
assign x_22540 = v_2201 | ~v_100;
assign x_22541 = v_2201 | ~v_93;
assign x_22542 = v_2200 | ~v_2052;
assign x_22543 = v_2200 | ~v_2053;
assign x_22544 = v_2200 | ~v_2054;
assign x_22545 = v_2200 | ~v_2055;
assign x_22546 = v_2200 | ~v_1058;
assign x_22547 = v_2200 | ~v_1059;
assign x_22548 = v_2200 | ~v_1060;
assign x_22549 = v_2200 | ~v_1061;
assign x_22550 = v_2200 | ~v_950;
assign x_22551 = v_2200 | ~v_951;
assign x_22552 = v_2200 | ~v_952;
assign x_22553 = v_2200 | ~v_953;
assign x_22554 = v_2200 | ~v_784;
assign x_22555 = v_2200 | ~v_787;
assign x_22556 = v_2200 | ~v_2104;
assign x_22557 = v_2200 | ~v_2105;
assign x_22558 = v_2200 | ~v_2106;
assign x_22559 = v_2200 | ~v_2107;
assign x_22560 = v_2200 | ~v_2188;
assign x_22561 = v_2200 | ~v_2189;
assign x_22562 = v_2200 | ~v_2190;
assign x_22563 = v_2200 | ~v_2191;
assign x_22564 = v_2200 | ~v_2060;
assign x_22565 = v_2200 | ~v_2063;
assign x_22566 = v_2200 | ~v_960;
assign x_22567 = v_2200 | ~v_961;
assign x_22568 = v_2200 | ~v_1110;
assign x_22569 = v_2200 | ~v_1111;
assign x_22570 = v_2200 | ~v_1070;
assign x_22571 = v_2200 | ~v_1071;
assign x_22572 = v_2200 | ~v_1112;
assign x_22573 = v_2200 | ~v_1113;
assign x_22574 = v_2200 | ~v_183;
assign x_22575 = v_2200 | ~v_167;
assign x_22576 = v_2200 | ~v_166;
assign x_22577 = v_2200 | ~v_146;
assign x_22578 = v_2200 | ~v_145;
assign x_22579 = v_2200 | ~v_144;
assign x_22580 = v_2200 | ~v_143;
assign x_22581 = v_2200 | ~v_142;
assign x_22582 = v_2200 | ~v_61;
assign x_22583 = v_2200 | ~v_59;
assign x_22584 = v_2200 | ~v_58;
assign x_22585 = v_2200 | ~v_51;
assign x_22586 = v_2199 | ~v_2037;
assign x_22587 = v_2199 | ~v_2038;
assign x_22588 = v_2199 | ~v_2039;
assign x_22589 = v_2199 | ~v_2040;
assign x_22590 = v_2199 | ~v_1043;
assign x_22591 = v_2199 | ~v_1044;
assign x_22592 = v_2199 | ~v_1045;
assign x_22593 = v_2199 | ~v_1046;
assign x_22594 = v_2199 | ~v_935;
assign x_22595 = v_2199 | ~v_936;
assign x_22596 = v_2199 | ~v_937;
assign x_22597 = v_2199 | ~v_938;
assign x_22598 = v_2199 | ~v_751;
assign x_22599 = v_2199 | ~v_754;
assign x_22600 = v_2199 | ~v_2099;
assign x_22601 = v_2199 | ~v_2100;
assign x_22602 = v_2199 | ~v_2101;
assign x_22603 = v_2199 | ~v_2102;
assign x_22604 = v_2199 | ~v_2183;
assign x_22605 = v_2199 | ~v_2184;
assign x_22606 = v_2199 | ~v_2185;
assign x_22607 = v_2199 | ~v_2186;
assign x_22608 = v_2199 | ~v_2045;
assign x_22609 = v_2199 | ~v_2048;
assign x_22610 = v_2199 | ~v_945;
assign x_22611 = v_2199 | ~v_946;
assign x_22612 = v_2199 | ~v_1105;
assign x_22613 = v_2199 | ~v_1106;
assign x_22614 = v_2199 | ~v_1055;
assign x_22615 = v_2199 | ~v_1056;
assign x_22616 = v_2199 | ~v_1107;
assign x_22617 = v_2199 | ~v_1108;
assign x_22618 = v_2199 | ~v_182;
assign x_22619 = v_2199 | ~v_163;
assign x_22620 = v_2199 | ~v_162;
assign x_22621 = v_2199 | ~v_138;
assign x_22622 = v_2199 | ~v_137;
assign x_22623 = v_2199 | ~v_136;
assign x_22624 = v_2199 | ~v_135;
assign x_22625 = v_2199 | ~v_134;
assign x_22626 = v_2199 | ~v_18;
assign x_22627 = v_2199 | ~v_16;
assign x_22628 = v_2199 | ~v_15;
assign x_22629 = v_2199 | ~v_8;
assign x_22630 = ~v_2197 | ~v_2192 | ~v_2187 | v_2198;
assign x_22631 = v_2197 | ~v_2067;
assign x_22632 = v_2197 | ~v_2068;
assign x_22633 = v_2197 | ~v_2069;
assign x_22634 = v_2197 | ~v_2070;
assign x_22635 = v_2197 | ~v_1073;
assign x_22636 = v_2197 | ~v_1074;
assign x_22637 = v_2197 | ~v_1075;
assign x_22638 = v_2197 | ~v_1076;
assign x_22639 = v_2197 | ~v_813;
assign x_22640 = v_2197 | ~v_814;
assign x_22641 = v_2197 | ~v_815;
assign x_22642 = v_2197 | ~v_816;
assign x_22643 = v_2197 | ~v_817;
assign x_22644 = v_2197 | ~v_820;
assign x_22645 = v_2197 | ~v_2071;
assign x_22646 = v_2197 | ~v_2072;
assign x_22647 = v_2197 | ~v_2073;
assign x_22648 = v_2197 | ~v_2074;
assign x_22649 = v_2197 | ~v_2193;
assign x_22650 = v_2197 | ~v_2194;
assign x_22651 = v_2197 | ~v_2195;
assign x_22652 = v_2197 | ~v_2196;
assign x_22653 = v_2197 | ~v_2075;
assign x_22654 = v_2197 | ~v_2078;
assign x_22655 = v_2197 | ~v_837;
assign x_22656 = v_2197 | ~v_838;
assign x_22657 = v_2197 | ~v_1081;
assign x_22658 = v_2197 | ~v_1082;
assign x_22659 = v_2197 | ~v_1083;
assign x_22660 = v_2197 | ~v_1084;
assign x_22661 = v_2197 | ~v_1085;
assign x_22662 = v_2197 | ~v_1086;
assign x_22663 = v_2197 | ~v_184;
assign x_22664 = v_2197 | ~v_171;
assign x_22665 = v_2197 | ~v_170;
assign x_22666 = v_2197 | ~v_160;
assign x_22667 = v_2197 | ~v_150;
assign x_22668 = v_2197 | ~v_148;
assign x_22669 = v_2197 | ~v_147;
assign x_22670 = v_2197 | ~v_103;
assign x_22671 = v_2197 | ~v_102;
assign x_22672 = v_2197 | ~v_100;
assign x_22673 = v_2197 | ~v_97;
assign x_22674 = v_2197 | ~v_93;
assign x_22675 = ~v_127 | ~v_141 | v_2196;
assign x_22676 = ~v_121 | ~v_141 | v_2195;
assign x_22677 = ~v_112 | v_141 | v_2194;
assign x_22678 = ~v_106 | v_141 | v_2193;
assign x_22679 = v_2192 | ~v_2052;
assign x_22680 = v_2192 | ~v_2053;
assign x_22681 = v_2192 | ~v_2054;
assign x_22682 = v_2192 | ~v_2055;
assign x_22683 = v_2192 | ~v_1058;
assign x_22684 = v_2192 | ~v_1059;
assign x_22685 = v_2192 | ~v_1060;
assign x_22686 = v_2192 | ~v_1061;
assign x_22687 = v_2192 | ~v_780;
assign x_22688 = v_2192 | ~v_781;
assign x_22689 = v_2192 | ~v_782;
assign x_22690 = v_2192 | ~v_783;
assign x_22691 = v_2192 | ~v_784;
assign x_22692 = v_2192 | ~v_787;
assign x_22693 = v_2192 | ~v_2056;
assign x_22694 = v_2192 | ~v_2057;
assign x_22695 = v_2192 | ~v_2058;
assign x_22696 = v_2192 | ~v_2059;
assign x_22697 = v_2192 | ~v_2188;
assign x_22698 = v_2192 | ~v_2189;
assign x_22699 = v_2192 | ~v_2190;
assign x_22700 = v_2192 | ~v_2191;
assign x_22701 = v_2192 | ~v_2060;
assign x_22702 = v_2192 | ~v_2063;
assign x_22703 = v_2192 | ~v_804;
assign x_22704 = v_2192 | ~v_805;
assign x_22705 = v_2192 | ~v_1066;
assign x_22706 = v_2192 | ~v_1067;
assign x_22707 = v_2192 | ~v_1068;
assign x_22708 = v_2192 | ~v_1069;
assign x_22709 = v_2192 | ~v_1070;
assign x_22710 = v_2192 | ~v_1071;
assign x_22711 = v_2192 | ~v_183;
assign x_22712 = v_2192 | ~v_167;
assign x_22713 = v_2192 | ~v_166;
assign x_22714 = v_2192 | ~v_159;
assign x_22715 = v_2192 | ~v_145;
assign x_22716 = v_2192 | ~v_143;
assign x_22717 = v_2192 | ~v_142;
assign x_22718 = v_2192 | ~v_61;
assign x_22719 = v_2192 | ~v_60;
assign x_22720 = v_2192 | ~v_58;
assign x_22721 = v_2192 | ~v_55;
assign x_22722 = v_2192 | ~v_51;
assign x_22723 = ~v_85 | ~v_141 | v_2191;
assign x_22724 = ~v_79 | ~v_141 | v_2190;
assign x_22725 = ~v_70 | v_141 | v_2189;
assign x_22726 = ~v_64 | v_141 | v_2188;
assign x_22727 = v_2187 | ~v_2037;
assign x_22728 = v_2187 | ~v_2038;
assign x_22729 = v_2187 | ~v_2039;
assign x_22730 = v_2187 | ~v_2040;
assign x_22731 = v_2187 | ~v_1043;
assign x_22732 = v_2187 | ~v_1044;
assign x_22733 = v_2187 | ~v_1045;
assign x_22734 = v_2187 | ~v_1046;
assign x_22735 = v_2187 | ~v_747;
assign x_22736 = v_2187 | ~v_748;
assign x_22737 = v_2187 | ~v_749;
assign x_22738 = v_2187 | ~v_750;
assign x_22739 = v_2187 | ~v_751;
assign x_22740 = v_2187 | ~v_754;
assign x_22741 = v_2187 | ~v_2041;
assign x_22742 = v_2187 | ~v_2042;
assign x_22743 = v_2187 | ~v_2043;
assign x_22744 = v_2187 | ~v_2044;
assign x_22745 = v_2187 | ~v_2183;
assign x_22746 = v_2187 | ~v_2184;
assign x_22747 = v_2187 | ~v_2185;
assign x_22748 = v_2187 | ~v_2186;
assign x_22749 = v_2187 | ~v_2045;
assign x_22750 = v_2187 | ~v_2048;
assign x_22751 = v_2187 | ~v_771;
assign x_22752 = v_2187 | ~v_772;
assign x_22753 = v_2187 | ~v_1051;
assign x_22754 = v_2187 | ~v_1052;
assign x_22755 = v_2187 | ~v_1053;
assign x_22756 = v_2187 | ~v_1054;
assign x_22757 = v_2187 | ~v_1055;
assign x_22758 = v_2187 | ~v_1056;
assign x_22759 = v_2187 | ~v_182;
assign x_22760 = v_2187 | ~v_163;
assign x_22761 = v_2187 | ~v_162;
assign x_22762 = v_2187 | ~v_155;
assign x_22763 = v_2187 | ~v_137;
assign x_22764 = v_2187 | ~v_135;
assign x_22765 = v_2187 | ~v_134;
assign x_22766 = v_2187 | ~v_18;
assign x_22767 = v_2187 | ~v_17;
assign x_22768 = v_2187 | ~v_15;
assign x_22769 = v_2187 | ~v_12;
assign x_22770 = v_2187 | ~v_8;
assign x_22771 = ~v_43 | ~v_141 | v_2186;
assign x_22772 = ~v_37 | ~v_141 | v_2185;
assign x_22773 = ~v_28 | v_141 | v_2184;
assign x_22774 = ~v_22 | v_141 | v_2183;
assign x_22775 = ~v_2181 | ~v_2180 | ~v_2179 | v_2182;
assign x_22776 = v_2181 | ~v_2067;
assign x_22777 = v_2181 | ~v_2068;
assign x_22778 = v_2181 | ~v_2069;
assign x_22779 = v_2181 | ~v_2070;
assign x_22780 = v_2181 | ~v_919;
assign x_22781 = v_2181 | ~v_920;
assign x_22782 = v_2181 | ~v_817;
assign x_22783 = v_2181 | ~v_818;
assign x_22784 = v_2181 | ~v_819;
assign x_22785 = v_2181 | ~v_820;
assign x_22786 = v_2181 | ~v_821;
assign x_22787 = v_2181 | ~v_822;
assign x_22788 = v_2181 | ~v_2125;
assign x_22789 = v_2181 | ~v_2126;
assign x_22790 = v_2181 | ~v_2127;
assign x_22791 = v_2181 | ~v_2128;
assign x_22792 = v_2181 | ~v_2075;
assign x_22793 = v_2181 | ~v_2076;
assign x_22794 = v_2181 | ~v_2077;
assign x_22795 = v_2181 | ~v_2078;
assign x_22796 = v_2181 | ~v_2079;
assign x_22797 = v_2181 | ~v_2080;
assign x_22798 = v_2181 | ~v_1037;
assign x_22799 = v_2181 | ~v_1038;
assign x_22800 = v_2181 | ~v_1039;
assign x_22801 = v_2181 | ~v_1040;
assign x_22802 = v_2181 | ~v_927;
assign x_22803 = v_2181 | ~v_928;
assign x_22804 = v_2181 | ~v_839;
assign x_22805 = v_2181 | ~v_840;
assign x_22806 = v_2181 | ~v_931;
assign x_22807 = v_2181 | ~v_932;
assign x_22808 = v_2181 | ~v_184;
assign x_22809 = v_2181 | ~v_170;
assign x_22810 = v_2181 | ~v_169;
assign x_22811 = v_2181 | ~v_151;
assign x_22812 = v_2181 | ~v_150;
assign x_22813 = v_2181 | ~v_149;
assign x_22814 = v_2181 | ~v_147;
assign x_22815 = v_2181 | ~v_103;
assign x_22816 = v_2181 | ~v_101;
assign x_22817 = v_2181 | ~v_100;
assign x_22818 = v_2181 | ~v_98;
assign x_22819 = v_2181 | ~v_96;
assign x_22820 = v_2180 | ~v_2052;
assign x_22821 = v_2180 | ~v_2053;
assign x_22822 = v_2180 | ~v_2054;
assign x_22823 = v_2180 | ~v_2055;
assign x_22824 = v_2180 | ~v_904;
assign x_22825 = v_2180 | ~v_905;
assign x_22826 = v_2180 | ~v_784;
assign x_22827 = v_2180 | ~v_785;
assign x_22828 = v_2180 | ~v_786;
assign x_22829 = v_2180 | ~v_787;
assign x_22830 = v_2180 | ~v_788;
assign x_22831 = v_2180 | ~v_789;
assign x_22832 = v_2180 | ~v_2120;
assign x_22833 = v_2180 | ~v_2121;
assign x_22834 = v_2180 | ~v_2122;
assign x_22835 = v_2180 | ~v_2123;
assign x_22836 = v_2180 | ~v_2060;
assign x_22837 = v_2180 | ~v_2061;
assign x_22838 = v_2180 | ~v_2062;
assign x_22839 = v_2180 | ~v_2063;
assign x_22840 = v_2180 | ~v_2064;
assign x_22841 = v_2180 | ~v_2065;
assign x_22842 = v_2180 | ~v_1032;
assign x_22843 = v_2180 | ~v_1033;
assign x_22844 = v_2180 | ~v_1034;
assign x_22845 = v_2180 | ~v_1035;
assign x_22846 = v_2180 | ~v_912;
assign x_22847 = v_2180 | ~v_913;
assign x_22848 = v_2180 | ~v_806;
assign x_22849 = v_2180 | ~v_807;
assign x_22850 = v_2180 | ~v_916;
assign x_22851 = v_2180 | ~v_917;
assign x_22852 = v_2180 | ~v_183;
assign x_22853 = v_2180 | ~v_166;
assign x_22854 = v_2180 | ~v_165;
assign x_22855 = v_2180 | ~v_146;
assign x_22856 = v_2180 | ~v_145;
assign x_22857 = v_2180 | ~v_144;
assign x_22858 = v_2180 | ~v_142;
assign x_22859 = v_2180 | ~v_61;
assign x_22860 = v_2180 | ~v_59;
assign x_22861 = v_2180 | ~v_58;
assign x_22862 = v_2180 | ~v_56;
assign x_22863 = v_2180 | ~v_54;
assign x_22864 = v_2179 | ~v_2037;
assign x_22865 = v_2179 | ~v_2038;
assign x_22866 = v_2179 | ~v_2039;
assign x_22867 = v_2179 | ~v_2040;
assign x_22868 = v_2179 | ~v_889;
assign x_22869 = v_2179 | ~v_890;
assign x_22870 = v_2179 | ~v_751;
assign x_22871 = v_2179 | ~v_752;
assign x_22872 = v_2179 | ~v_753;
assign x_22873 = v_2179 | ~v_754;
assign x_22874 = v_2179 | ~v_755;
assign x_22875 = v_2179 | ~v_756;
assign x_22876 = v_2179 | ~v_2115;
assign x_22877 = v_2179 | ~v_2116;
assign x_22878 = v_2179 | ~v_2117;
assign x_22879 = v_2179 | ~v_2118;
assign x_22880 = v_2179 | ~v_2045;
assign x_22881 = v_2179 | ~v_2046;
assign x_22882 = v_2179 | ~v_2047;
assign x_22883 = v_2179 | ~v_2048;
assign x_22884 = v_2179 | ~v_2049;
assign x_22885 = v_2179 | ~v_2050;
assign x_22886 = v_2179 | ~v_1027;
assign x_22887 = v_2179 | ~v_1028;
assign x_22888 = v_2179 | ~v_1029;
assign x_22889 = v_2179 | ~v_1030;
assign x_22890 = v_2179 | ~v_897;
assign x_22891 = v_2179 | ~v_898;
assign x_22892 = v_2179 | ~v_773;
assign x_22893 = v_2179 | ~v_774;
assign x_22894 = v_2179 | ~v_901;
assign x_22895 = v_2179 | ~v_902;
assign x_22896 = v_2179 | ~v_182;
assign x_22897 = v_2179 | ~v_162;
assign x_22898 = v_2179 | ~v_161;
assign x_22899 = v_2179 | ~v_138;
assign x_22900 = v_2179 | ~v_137;
assign x_22901 = v_2179 | ~v_136;
assign x_22902 = v_2179 | ~v_134;
assign x_22903 = v_2179 | ~v_18;
assign x_22904 = v_2179 | ~v_16;
assign x_22905 = v_2179 | ~v_15;
assign x_22906 = v_2179 | ~v_13;
assign x_22907 = v_2179 | ~v_11;
assign x_22908 = ~v_2177 | ~v_2176 | ~v_2175 | v_2178;
assign x_22909 = v_2177 | ~v_2067;
assign x_22910 = v_2177 | ~v_2068;
assign x_22911 = v_2177 | ~v_2069;
assign x_22912 = v_2177 | ~v_2070;
assign x_22913 = v_2177 | ~v_1183;
assign x_22914 = v_2177 | ~v_1184;
assign x_22915 = v_2177 | ~v_1185;
assign x_22916 = v_2177 | ~v_1186;
assign x_22917 = v_2177 | ~v_817;
assign x_22918 = v_2177 | ~v_1011;
assign x_22919 = v_2177 | ~v_1012;
assign x_22920 = v_2177 | ~v_820;
assign x_22921 = v_2177 | ~v_1013;
assign x_22922 = v_2177 | ~v_1014;
assign x_22923 = v_2177 | ~v_2161;
assign x_22924 = v_2177 | ~v_2162;
assign x_22925 = v_2177 | ~v_2163;
assign x_22926 = v_2177 | ~v_2164;
assign x_22927 = v_2177 | ~v_2075;
assign x_22928 = v_2177 | ~v_2141;
assign x_22929 = v_2177 | ~v_2142;
assign x_22930 = v_2177 | ~v_2078;
assign x_22931 = v_2177 | ~v_2143;
assign x_22932 = v_2177 | ~v_2144;
assign x_22933 = v_2177 | ~v_1193;
assign x_22934 = v_2177 | ~v_1241;
assign x_22935 = v_2177 | ~v_1194;
assign x_22936 = v_2177 | ~v_1242;
assign x_22937 = v_2177 | ~v_1023;
assign x_22938 = v_2177 | ~v_1024;
assign x_22939 = v_2177 | ~v_1243;
assign x_22940 = v_2177 | ~v_1244;
assign x_22941 = v_2177 | ~v_184;
assign x_22942 = v_2177 | ~v_171;
assign x_22943 = v_2177 | ~v_170;
assign x_22944 = v_2177 | ~v_169;
assign x_22945 = v_2177 | ~v_149;
assign x_22946 = v_2177 | ~v_148;
assign x_22947 = v_2177 | ~v_147;
assign x_22948 = v_2177 | ~v_103;
assign x_22949 = v_2177 | ~v_102;
assign x_22950 = v_2177 | ~v_101;
assign x_22951 = v_2177 | ~v_100;
assign x_22952 = v_2177 | ~v_99;
assign x_22953 = v_2176 | ~v_2052;
assign x_22954 = v_2176 | ~v_2053;
assign x_22955 = v_2176 | ~v_2054;
assign x_22956 = v_2176 | ~v_2055;
assign x_22957 = v_2176 | ~v_1168;
assign x_22958 = v_2176 | ~v_1169;
assign x_22959 = v_2176 | ~v_1170;
assign x_22960 = v_2176 | ~v_1171;
assign x_22961 = v_2176 | ~v_784;
assign x_22962 = v_2176 | ~v_996;
assign x_22963 = v_2176 | ~v_997;
assign x_22964 = v_2176 | ~v_787;
assign x_22965 = v_2176 | ~v_998;
assign x_22966 = v_2176 | ~v_999;
assign x_22967 = v_2176 | ~v_2156;
assign x_22968 = v_2176 | ~v_2157;
assign x_22969 = v_2176 | ~v_2158;
assign x_22970 = v_2176 | ~v_2159;
assign x_22971 = v_2176 | ~v_2060;
assign x_22972 = v_2176 | ~v_2136;
assign x_22973 = v_2176 | ~v_2137;
assign x_22974 = v_2176 | ~v_2063;
assign x_22975 = v_2176 | ~v_2138;
assign x_22976 = v_2176 | ~v_2139;
assign x_22977 = v_2176 | ~v_1178;
assign x_22978 = v_2176 | ~v_1236;
assign x_22979 = v_2176 | ~v_1179;
assign x_22980 = v_2176 | ~v_1237;
assign x_22981 = v_2176 | ~v_1008;
assign x_22982 = v_2176 | ~v_1009;
assign x_22983 = v_2176 | ~v_1238;
assign x_22984 = v_2176 | ~v_1239;
assign x_22985 = v_2176 | ~v_183;
assign x_22986 = v_2176 | ~v_167;
assign x_22987 = v_2176 | ~v_166;
assign x_22988 = v_2176 | ~v_165;
assign x_22989 = v_2176 | ~v_144;
assign x_22990 = v_2176 | ~v_143;
assign x_22991 = v_2176 | ~v_142;
assign x_22992 = v_2176 | ~v_61;
assign x_22993 = v_2176 | ~v_60;
assign x_22994 = v_2176 | ~v_59;
assign x_22995 = v_2176 | ~v_58;
assign x_22996 = v_2176 | ~v_57;
assign x_22997 = v_2175 | ~v_2037;
assign x_22998 = v_2175 | ~v_2038;
assign x_22999 = v_2175 | ~v_2039;
assign x_23000 = v_2175 | ~v_2040;
assign x_23001 = v_2175 | ~v_1153;
assign x_23002 = v_2175 | ~v_1154;
assign x_23003 = v_2175 | ~v_1155;
assign x_23004 = v_2175 | ~v_1156;
assign x_23005 = v_2175 | ~v_751;
assign x_23006 = v_2175 | ~v_981;
assign x_23007 = v_2175 | ~v_982;
assign x_23008 = v_2175 | ~v_754;
assign x_23009 = v_2175 | ~v_983;
assign x_23010 = v_2175 | ~v_984;
assign x_23011 = v_2175 | ~v_2151;
assign x_23012 = v_2175 | ~v_2152;
assign x_23013 = v_2175 | ~v_2153;
assign x_23014 = v_2175 | ~v_2154;
assign x_23015 = v_2175 | ~v_2045;
assign x_23016 = v_2175 | ~v_2131;
assign x_23017 = v_2175 | ~v_2132;
assign x_23018 = v_2175 | ~v_2048;
assign x_23019 = v_2175 | ~v_2133;
assign x_23020 = v_2175 | ~v_2134;
assign x_23021 = v_2175 | ~v_1163;
assign x_23022 = v_2175 | ~v_1231;
assign x_23023 = v_2175 | ~v_1164;
assign x_23024 = v_2175 | ~v_1232;
assign x_23025 = v_2175 | ~v_1233;
assign x_23026 = v_2175 | ~v_1234;
assign x_23027 = v_2175 | ~v_182;
assign x_23028 = v_2175 | ~v_163;
assign x_23029 = v_2175 | ~v_162;
assign x_23030 = v_2175 | ~v_161;
assign x_23031 = v_2175 | ~v_136;
assign x_23032 = v_2175 | ~v_135;
assign x_23033 = v_2175 | ~v_134;
assign x_23034 = v_2175 | ~v_993;
assign x_23035 = v_2175 | ~v_994;
assign x_23036 = v_2175 | ~v_18;
assign x_23037 = v_2175 | ~v_17;
assign x_23038 = v_2175 | ~v_16;
assign x_23039 = v_2175 | ~v_15;
assign x_23040 = v_2175 | ~v_14;
assign x_23041 = ~v_2173 | ~v_2172 | ~v_2171 | v_2174;
assign x_23042 = v_2173 | ~v_2067;
assign x_23043 = v_2173 | ~v_2068;
assign x_23044 = v_2173 | ~v_2069;
assign x_23045 = v_2173 | ~v_2070;
assign x_23046 = v_2173 | ~v_1183;
assign x_23047 = v_2173 | ~v_1184;
assign x_23048 = v_2173 | ~v_1185;
assign x_23049 = v_2173 | ~v_1186;
assign x_23050 = v_2173 | ~v_919;
assign x_23051 = v_2173 | ~v_920;
assign x_23052 = v_2173 | ~v_817;
assign x_23053 = v_2173 | ~v_820;
assign x_23054 = v_2173 | ~v_2161;
assign x_23055 = v_2173 | ~v_2162;
assign x_23056 = v_2173 | ~v_2163;
assign x_23057 = v_2173 | ~v_2164;
assign x_23058 = v_2173 | ~v_2125;
assign x_23059 = v_2173 | ~v_2126;
assign x_23060 = v_2173 | ~v_2127;
assign x_23061 = v_2173 | ~v_2128;
assign x_23062 = v_2173 | ~v_2075;
assign x_23063 = v_2173 | ~v_2078;
assign x_23064 = v_2173 | ~v_1209;
assign x_23065 = v_2173 | ~v_1210;
assign x_23066 = v_2173 | ~v_1193;
assign x_23067 = v_2173 | ~v_1194;
assign x_23068 = v_2173 | ~v_927;
assign x_23069 = v_2173 | ~v_928;
assign x_23070 = v_2173 | ~v_931;
assign x_23071 = v_2173 | ~v_932;
assign x_23072 = v_2173 | ~v_1211;
assign x_23073 = v_2173 | ~v_1212;
assign x_23074 = v_2173 | ~v_184;
assign x_23075 = v_2173 | ~v_172;
assign x_23076 = v_2173 | ~v_171;
assign x_23077 = v_2173 | ~v_170;
assign x_23078 = v_2173 | ~v_169;
assign x_23079 = v_2173 | ~v_150;
assign x_23080 = v_2173 | ~v_149;
assign x_23081 = v_2173 | ~v_147;
assign x_23082 = v_2173 | ~v_102;
assign x_23083 = v_2173 | ~v_101;
assign x_23084 = v_2173 | ~v_100;
assign x_23085 = v_2173 | ~v_96;
assign x_23086 = v_2172 | ~v_2052;
assign x_23087 = v_2172 | ~v_2053;
assign x_23088 = v_2172 | ~v_2054;
assign x_23089 = v_2172 | ~v_2055;
assign x_23090 = v_2172 | ~v_1168;
assign x_23091 = v_2172 | ~v_1169;
assign x_23092 = v_2172 | ~v_1170;
assign x_23093 = v_2172 | ~v_1171;
assign x_23094 = v_2172 | ~v_904;
assign x_23095 = v_2172 | ~v_905;
assign x_23096 = v_2172 | ~v_784;
assign x_23097 = v_2172 | ~v_787;
assign x_23098 = v_2172 | ~v_2156;
assign x_23099 = v_2172 | ~v_2157;
assign x_23100 = v_2172 | ~v_2158;
assign x_23101 = v_2172 | ~v_2159;
assign x_23102 = v_2172 | ~v_2120;
assign x_23103 = v_2172 | ~v_2121;
assign x_23104 = v_2172 | ~v_2122;
assign x_23105 = v_2172 | ~v_2123;
assign x_23106 = v_2172 | ~v_2060;
assign x_23107 = v_2172 | ~v_2063;
assign x_23108 = v_2172 | ~v_1204;
assign x_23109 = v_2172 | ~v_1205;
assign x_23110 = v_2172 | ~v_1178;
assign x_23111 = v_2172 | ~v_1179;
assign x_23112 = v_2172 | ~v_912;
assign x_23113 = v_2172 | ~v_913;
assign x_23114 = v_2172 | ~v_916;
assign x_23115 = v_2172 | ~v_917;
assign x_23116 = v_2172 | ~v_1206;
assign x_23117 = v_2172 | ~v_1207;
assign x_23118 = v_2172 | ~v_183;
assign x_23119 = v_2172 | ~v_168;
assign x_23120 = v_2172 | ~v_167;
assign x_23121 = v_2172 | ~v_166;
assign x_23122 = v_2172 | ~v_165;
assign x_23123 = v_2172 | ~v_145;
assign x_23124 = v_2172 | ~v_144;
assign x_23125 = v_2172 | ~v_142;
assign x_23126 = v_2172 | ~v_60;
assign x_23127 = v_2172 | ~v_59;
assign x_23128 = v_2172 | ~v_58;
assign x_23129 = v_2172 | ~v_54;
assign x_23130 = v_2171 | ~v_2037;
assign x_23131 = v_2171 | ~v_2038;
assign x_23132 = v_2171 | ~v_2039;
assign x_23133 = v_2171 | ~v_2040;
assign x_23134 = v_2171 | ~v_1153;
assign x_23135 = v_2171 | ~v_1154;
assign x_23136 = v_2171 | ~v_1155;
assign x_23137 = v_2171 | ~v_1156;
assign x_23138 = v_2171 | ~v_889;
assign x_23139 = v_2171 | ~v_890;
assign x_23140 = v_2171 | ~v_751;
assign x_23141 = v_2171 | ~v_754;
assign x_23142 = v_2171 | ~v_2151;
assign x_23143 = v_2171 | ~v_2152;
assign x_23144 = v_2171 | ~v_2153;
assign x_23145 = v_2171 | ~v_2154;
assign x_23146 = v_2171 | ~v_2115;
assign x_23147 = v_2171 | ~v_2116;
assign x_23148 = v_2171 | ~v_2117;
assign x_23149 = v_2171 | ~v_2118;
assign x_23150 = v_2171 | ~v_2045;
assign x_23151 = v_2171 | ~v_2048;
assign x_23152 = v_2171 | ~v_1199;
assign x_23153 = v_2171 | ~v_1200;
assign x_23154 = v_2171 | ~v_1163;
assign x_23155 = v_2171 | ~v_1164;
assign x_23156 = v_2171 | ~v_897;
assign x_23157 = v_2171 | ~v_898;
assign x_23158 = v_2171 | ~v_901;
assign x_23159 = v_2171 | ~v_902;
assign x_23160 = v_2171 | ~v_1201;
assign x_23161 = v_2171 | ~v_1202;
assign x_23162 = v_2171 | ~v_182;
assign x_23163 = v_2171 | ~v_164;
assign x_23164 = v_2171 | ~v_163;
assign x_23165 = v_2171 | ~v_162;
assign x_23166 = v_2171 | ~v_161;
assign x_23167 = v_2171 | ~v_137;
assign x_23168 = v_2171 | ~v_136;
assign x_23169 = v_2171 | ~v_134;
assign x_23170 = v_2171 | ~v_17;
assign x_23171 = v_2171 | ~v_16;
assign x_23172 = v_2171 | ~v_15;
assign x_23173 = v_2171 | ~v_11;
assign x_23174 = ~v_2169 | ~v_2168 | ~v_2167 | v_2170;
assign x_23175 = v_2169 | ~v_2067;
assign x_23176 = v_2169 | ~v_2068;
assign x_23177 = v_2169 | ~v_2069;
assign x_23178 = v_2169 | ~v_2070;
assign x_23179 = v_2169 | ~v_1183;
assign x_23180 = v_2169 | ~v_1184;
assign x_23181 = v_2169 | ~v_1185;
assign x_23182 = v_2169 | ~v_1186;
assign x_23183 = v_2169 | ~v_965;
assign x_23184 = v_2169 | ~v_966;
assign x_23185 = v_2169 | ~v_967;
assign x_23186 = v_2169 | ~v_968;
assign x_23187 = v_2169 | ~v_817;
assign x_23188 = v_2169 | ~v_820;
assign x_23189 = v_2169 | ~v_2161;
assign x_23190 = v_2169 | ~v_2162;
assign x_23191 = v_2169 | ~v_2163;
assign x_23192 = v_2169 | ~v_2164;
assign x_23193 = v_2169 | ~v_2109;
assign x_23194 = v_2169 | ~v_2110;
assign x_23195 = v_2169 | ~v_2111;
assign x_23196 = v_2169 | ~v_2112;
assign x_23197 = v_2169 | ~v_2075;
assign x_23198 = v_2169 | ~v_2078;
assign x_23199 = v_2169 | ~v_1225;
assign x_23200 = v_2169 | ~v_1226;
assign x_23201 = v_2169 | ~v_1227;
assign x_23202 = v_2169 | ~v_1228;
assign x_23203 = v_2169 | ~v_1193;
assign x_23204 = v_2169 | ~v_1194;
assign x_23205 = v_2169 | ~v_975;
assign x_23206 = v_2169 | ~v_976;
assign x_23207 = v_2169 | ~v_184;
assign x_23208 = v_2169 | ~v_171;
assign x_23209 = v_2169 | ~v_170;
assign x_23210 = v_2169 | ~v_169;
assign x_23211 = v_2169 | ~v_150;
assign x_23212 = v_2169 | ~v_149;
assign x_23213 = v_2169 | ~v_148;
assign x_23214 = v_2169 | ~v_103;
assign x_23215 = v_2169 | ~v_102;
assign x_23216 = v_2169 | ~v_101;
assign x_23217 = v_2169 | ~v_100;
assign x_23218 = v_2169 | ~v_95;
assign x_23219 = v_2168 | ~v_2052;
assign x_23220 = v_2168 | ~v_2053;
assign x_23221 = v_2168 | ~v_2054;
assign x_23222 = v_2168 | ~v_2055;
assign x_23223 = v_2168 | ~v_1168;
assign x_23224 = v_2168 | ~v_1169;
assign x_23225 = v_2168 | ~v_1170;
assign x_23226 = v_2168 | ~v_1171;
assign x_23227 = v_2168 | ~v_950;
assign x_23228 = v_2168 | ~v_951;
assign x_23229 = v_2168 | ~v_952;
assign x_23230 = v_2168 | ~v_953;
assign x_23231 = v_2168 | ~v_784;
assign x_23232 = v_2168 | ~v_787;
assign x_23233 = v_2168 | ~v_2156;
assign x_23234 = v_2168 | ~v_2157;
assign x_23235 = v_2168 | ~v_2158;
assign x_23236 = v_2168 | ~v_2159;
assign x_23237 = v_2168 | ~v_2104;
assign x_23238 = v_2168 | ~v_2105;
assign x_23239 = v_2168 | ~v_2106;
assign x_23240 = v_2168 | ~v_2107;
assign x_23241 = v_2168 | ~v_2060;
assign x_23242 = v_2168 | ~v_2063;
assign x_23243 = v_2168 | ~v_1220;
assign x_23244 = v_2168 | ~v_1221;
assign x_23245 = v_2168 | ~v_1222;
assign x_23246 = v_2168 | ~v_1223;
assign x_23247 = v_2168 | ~v_1178;
assign x_23248 = v_2168 | ~v_1179;
assign x_23249 = v_2168 | ~v_960;
assign x_23250 = v_2168 | ~v_961;
assign x_23251 = v_2168 | ~v_183;
assign x_23252 = v_2168 | ~v_167;
assign x_23253 = v_2168 | ~v_166;
assign x_23254 = v_2168 | ~v_165;
assign x_23255 = v_2168 | ~v_145;
assign x_23256 = v_2168 | ~v_144;
assign x_23257 = v_2168 | ~v_143;
assign x_23258 = v_2168 | ~v_61;
assign x_23259 = v_2168 | ~v_60;
assign x_23260 = v_2168 | ~v_59;
assign x_23261 = v_2168 | ~v_58;
assign x_23262 = v_2168 | ~v_53;
assign x_23263 = v_2167 | ~v_2037;
assign x_23264 = v_2167 | ~v_2038;
assign x_23265 = v_2167 | ~v_2039;
assign x_23266 = v_2167 | ~v_2040;
assign x_23267 = v_2167 | ~v_1153;
assign x_23268 = v_2167 | ~v_1154;
assign x_23269 = v_2167 | ~v_1155;
assign x_23270 = v_2167 | ~v_1156;
assign x_23271 = v_2167 | ~v_935;
assign x_23272 = v_2167 | ~v_936;
assign x_23273 = v_2167 | ~v_937;
assign x_23274 = v_2167 | ~v_938;
assign x_23275 = v_2167 | ~v_751;
assign x_23276 = v_2167 | ~v_754;
assign x_23277 = v_2167 | ~v_2151;
assign x_23278 = v_2167 | ~v_2152;
assign x_23279 = v_2167 | ~v_2153;
assign x_23280 = v_2167 | ~v_2154;
assign x_23281 = v_2167 | ~v_2099;
assign x_23282 = v_2167 | ~v_2100;
assign x_23283 = v_2167 | ~v_2101;
assign x_23284 = v_2167 | ~v_2102;
assign x_23285 = v_2167 | ~v_2045;
assign x_23286 = v_2167 | ~v_2048;
assign x_23287 = v_2167 | ~v_1215;
assign x_23288 = v_2167 | ~v_1216;
assign x_23289 = v_2167 | ~v_1217;
assign x_23290 = v_2167 | ~v_1218;
assign x_23291 = v_2167 | ~v_1163;
assign x_23292 = v_2167 | ~v_1164;
assign x_23293 = v_2167 | ~v_945;
assign x_23294 = v_2167 | ~v_946;
assign x_23295 = v_2167 | ~v_182;
assign x_23296 = v_2167 | ~v_163;
assign x_23297 = v_2167 | ~v_162;
assign x_23298 = v_2167 | ~v_161;
assign x_23299 = v_2167 | ~v_137;
assign x_23300 = v_2167 | ~v_136;
assign x_23301 = v_2167 | ~v_135;
assign x_23302 = v_2167 | ~v_18;
assign x_23303 = v_2167 | ~v_17;
assign x_23304 = v_2167 | ~v_16;
assign x_23305 = v_2167 | ~v_15;
assign x_23306 = v_2167 | ~v_10;
assign x_23307 = ~v_2165 | ~v_2160 | ~v_2155 | v_2166;
assign x_23308 = v_2165 | ~v_2067;
assign x_23309 = v_2165 | ~v_2068;
assign x_23310 = v_2165 | ~v_2069;
assign x_23311 = v_2165 | ~v_2070;
assign x_23312 = v_2165 | ~v_1183;
assign x_23313 = v_2165 | ~v_1184;
assign x_23314 = v_2165 | ~v_1185;
assign x_23315 = v_2165 | ~v_1186;
assign x_23316 = v_2165 | ~v_813;
assign x_23317 = v_2165 | ~v_814;
assign x_23318 = v_2165 | ~v_815;
assign x_23319 = v_2165 | ~v_816;
assign x_23320 = v_2165 | ~v_817;
assign x_23321 = v_2165 | ~v_820;
assign x_23322 = v_2165 | ~v_2161;
assign x_23323 = v_2165 | ~v_2162;
assign x_23324 = v_2165 | ~v_2163;
assign x_23325 = v_2165 | ~v_2164;
assign x_23326 = v_2165 | ~v_2071;
assign x_23327 = v_2165 | ~v_2072;
assign x_23328 = v_2165 | ~v_2073;
assign x_23329 = v_2165 | ~v_2074;
assign x_23330 = v_2165 | ~v_2075;
assign x_23331 = v_2165 | ~v_2078;
assign x_23332 = v_2165 | ~v_1191;
assign x_23333 = v_2165 | ~v_1192;
assign x_23334 = v_2165 | ~v_1193;
assign x_23335 = v_2165 | ~v_1194;
assign x_23336 = v_2165 | ~v_837;
assign x_23337 = v_2165 | ~v_838;
assign x_23338 = v_2165 | ~v_1195;
assign x_23339 = v_2165 | ~v_1196;
assign x_23340 = v_2165 | ~v_184;
assign x_23341 = v_2165 | ~v_171;
assign x_23342 = v_2165 | ~v_170;
assign x_23343 = v_2165 | ~v_169;
assign x_23344 = v_2165 | ~v_160;
assign x_23345 = v_2165 | ~v_151;
assign x_23346 = v_2165 | ~v_150;
assign x_23347 = v_2165 | ~v_148;
assign x_23348 = v_2165 | ~v_147;
assign x_23349 = v_2165 | ~v_103;
assign x_23350 = v_2165 | ~v_100;
assign x_23351 = v_2165 | ~v_97;
assign x_23352 = ~v_127 | ~v_174 | v_2164;
assign x_23353 = ~v_121 | ~v_173 | v_2163;
assign x_23354 = ~v_112 | v_174 | v_2162;
assign x_23355 = ~v_106 | v_173 | v_2161;
assign x_23356 = v_2160 | ~v_2052;
assign x_23357 = v_2160 | ~v_2053;
assign x_23358 = v_2160 | ~v_2054;
assign x_23359 = v_2160 | ~v_2055;
assign x_23360 = v_2160 | ~v_1168;
assign x_23361 = v_2160 | ~v_1169;
assign x_23362 = v_2160 | ~v_1170;
assign x_23363 = v_2160 | ~v_1171;
assign x_23364 = v_2160 | ~v_780;
assign x_23365 = v_2160 | ~v_781;
assign x_23366 = v_2160 | ~v_782;
assign x_23367 = v_2160 | ~v_783;
assign x_23368 = v_2160 | ~v_784;
assign x_23369 = v_2160 | ~v_787;
assign x_23370 = v_2160 | ~v_2156;
assign x_23371 = v_2160 | ~v_2157;
assign x_23372 = v_2160 | ~v_2158;
assign x_23373 = v_2160 | ~v_2159;
assign x_23374 = v_2160 | ~v_2056;
assign x_23375 = v_2160 | ~v_2057;
assign x_23376 = v_2160 | ~v_2058;
assign x_23377 = v_2160 | ~v_2059;
assign x_23378 = v_2160 | ~v_2060;
assign x_23379 = v_2160 | ~v_2063;
assign x_23380 = v_2160 | ~v_1176;
assign x_23381 = v_2160 | ~v_1177;
assign x_23382 = v_2160 | ~v_1178;
assign x_23383 = v_2160 | ~v_1179;
assign x_23384 = v_2160 | ~v_804;
assign x_23385 = v_2160 | ~v_805;
assign x_23386 = v_2160 | ~v_1180;
assign x_23387 = v_2160 | ~v_1181;
assign x_23388 = v_2160 | ~v_183;
assign x_23389 = v_2160 | ~v_167;
assign x_23390 = v_2160 | ~v_166;
assign x_23391 = v_2160 | ~v_165;
assign x_23392 = v_2160 | ~v_159;
assign x_23393 = v_2160 | ~v_146;
assign x_23394 = v_2160 | ~v_145;
assign x_23395 = v_2160 | ~v_143;
assign x_23396 = v_2160 | ~v_142;
assign x_23397 = v_2160 | ~v_61;
assign x_23398 = v_2160 | ~v_58;
assign x_23399 = v_2160 | ~v_55;
assign x_23400 = ~v_85 | ~v_174 | v_2159;
assign x_23401 = ~v_79 | ~v_173 | v_2158;
assign x_23402 = ~v_70 | v_174 | v_2157;
assign x_23403 = ~v_64 | v_173 | v_2156;
assign x_23404 = v_2155 | ~v_2037;
assign x_23405 = v_2155 | ~v_2038;
assign x_23406 = v_2155 | ~v_2039;
assign x_23407 = v_2155 | ~v_2040;
assign x_23408 = v_2155 | ~v_1153;
assign x_23409 = v_2155 | ~v_1154;
assign x_23410 = v_2155 | ~v_1155;
assign x_23411 = v_2155 | ~v_1156;
assign x_23412 = v_2155 | ~v_747;
assign x_23413 = v_2155 | ~v_748;
assign x_23414 = v_2155 | ~v_749;
assign x_23415 = v_2155 | ~v_750;
assign x_23416 = v_2155 | ~v_751;
assign x_23417 = v_2155 | ~v_754;
assign x_23418 = v_2155 | ~v_2151;
assign x_23419 = v_2155 | ~v_2152;
assign x_23420 = v_2155 | ~v_2153;
assign x_23421 = v_2155 | ~v_2154;
assign x_23422 = v_2155 | ~v_2041;
assign x_23423 = v_2155 | ~v_2042;
assign x_23424 = v_2155 | ~v_2043;
assign x_23425 = v_2155 | ~v_2044;
assign x_23426 = v_2155 | ~v_2045;
assign x_23427 = v_2155 | ~v_2048;
assign x_23428 = v_2155 | ~v_1161;
assign x_23429 = v_2155 | ~v_1162;
assign x_23430 = v_2155 | ~v_1163;
assign x_23431 = v_2155 | ~v_1164;
assign x_23432 = v_2155 | ~v_771;
assign x_23433 = v_2155 | ~v_772;
assign x_23434 = v_2155 | ~v_1165;
assign x_23435 = v_2155 | ~v_1166;
assign x_23436 = v_2155 | ~v_182;
assign x_23437 = v_2155 | ~v_163;
assign x_23438 = v_2155 | ~v_162;
assign x_23439 = v_2155 | ~v_161;
assign x_23440 = v_2155 | ~v_155;
assign x_23441 = v_2155 | ~v_138;
assign x_23442 = v_2155 | ~v_137;
assign x_23443 = v_2155 | ~v_135;
assign x_23444 = v_2155 | ~v_134;
assign x_23445 = v_2155 | ~v_18;
assign x_23446 = v_2155 | ~v_15;
assign x_23447 = v_2155 | ~v_12;
assign x_23448 = ~v_43 | ~v_174 | v_2154;
assign x_23449 = ~v_37 | ~v_173 | v_2153;
assign x_23450 = ~v_28 | v_174 | v_2152;
assign x_23451 = ~v_22 | v_173 | v_2151;
assign x_23452 = ~v_2149 | ~v_2148 | ~v_2147 | v_2150;
assign x_23453 = v_2149 | ~v_2067;
assign x_23454 = v_2149 | ~v_2068;
assign x_23455 = v_2149 | ~v_2069;
assign x_23456 = v_2149 | ~v_2070;
assign x_23457 = v_2149 | ~v_965;
assign x_23458 = v_2149 | ~v_966;
assign x_23459 = v_2149 | ~v_967;
assign x_23460 = v_2149 | ~v_968;
assign x_23461 = v_2149 | ~v_817;
assign x_23462 = v_2149 | ~v_818;
assign x_23463 = v_2149 | ~v_819;
assign x_23464 = v_2149 | ~v_820;
assign x_23465 = v_2149 | ~v_821;
assign x_23466 = v_2149 | ~v_822;
assign x_23467 = v_2149 | ~v_2109;
assign x_23468 = v_2149 | ~v_2110;
assign x_23469 = v_2149 | ~v_2111;
assign x_23470 = v_2149 | ~v_2112;
assign x_23471 = v_2149 | ~v_2075;
assign x_23472 = v_2149 | ~v_2076;
assign x_23473 = v_2149 | ~v_2077;
assign x_23474 = v_2149 | ~v_2078;
assign x_23475 = v_2149 | ~v_2079;
assign x_23476 = v_2149 | ~v_2080;
assign x_23477 = v_2149 | ~v_1147;
assign x_23478 = v_2149 | ~v_1148;
assign x_23479 = v_2149 | ~v_975;
assign x_23480 = v_2149 | ~v_976;
assign x_23481 = v_2149 | ~v_839;
assign x_23482 = v_2149 | ~v_840;
assign x_23483 = v_2149 | ~v_1149;
assign x_23484 = v_2149 | ~v_1150;
assign x_23485 = v_2149 | ~v_184;
assign x_23486 = v_2149 | ~v_170;
assign x_23487 = v_2149 | ~v_169;
assign x_23488 = v_2149 | ~v_150;
assign x_23489 = v_2149 | ~v_149;
assign x_23490 = v_2149 | ~v_148;
assign x_23491 = v_2149 | ~v_147;
assign x_23492 = v_2149 | ~v_103;
assign x_23493 = v_2149 | ~v_102;
assign x_23494 = v_2149 | ~v_101;
assign x_23495 = v_2149 | ~v_100;
assign x_23496 = v_2149 | ~v_98;
assign x_23497 = v_2148 | ~v_2052;
assign x_23498 = v_2148 | ~v_2053;
assign x_23499 = v_2148 | ~v_2054;
assign x_23500 = v_2148 | ~v_2055;
assign x_23501 = v_2148 | ~v_950;
assign x_23502 = v_2148 | ~v_951;
assign x_23503 = v_2148 | ~v_952;
assign x_23504 = v_2148 | ~v_953;
assign x_23505 = v_2148 | ~v_784;
assign x_23506 = v_2148 | ~v_785;
assign x_23507 = v_2148 | ~v_786;
assign x_23508 = v_2148 | ~v_787;
assign x_23509 = v_2148 | ~v_788;
assign x_23510 = v_2148 | ~v_789;
assign x_23511 = v_2148 | ~v_2104;
assign x_23512 = v_2148 | ~v_2105;
assign x_23513 = v_2148 | ~v_2106;
assign x_23514 = v_2148 | ~v_2107;
assign x_23515 = v_2148 | ~v_2060;
assign x_23516 = v_2148 | ~v_2061;
assign x_23517 = v_2148 | ~v_2062;
assign x_23518 = v_2148 | ~v_2063;
assign x_23519 = v_2148 | ~v_2064;
assign x_23520 = v_2148 | ~v_2065;
assign x_23521 = v_2148 | ~v_1142;
assign x_23522 = v_2148 | ~v_1143;
assign x_23523 = v_2148 | ~v_960;
assign x_23524 = v_2148 | ~v_961;
assign x_23525 = v_2148 | ~v_806;
assign x_23526 = v_2148 | ~v_807;
assign x_23527 = v_2148 | ~v_1144;
assign x_23528 = v_2148 | ~v_1145;
assign x_23529 = v_2148 | ~v_183;
assign x_23530 = v_2148 | ~v_166;
assign x_23531 = v_2148 | ~v_165;
assign x_23532 = v_2148 | ~v_145;
assign x_23533 = v_2148 | ~v_144;
assign x_23534 = v_2148 | ~v_143;
assign x_23535 = v_2148 | ~v_142;
assign x_23536 = v_2148 | ~v_61;
assign x_23537 = v_2148 | ~v_60;
assign x_23538 = v_2148 | ~v_59;
assign x_23539 = v_2148 | ~v_58;
assign x_23540 = v_2148 | ~v_56;
assign x_23541 = v_2147 | ~v_2037;
assign x_23542 = v_2147 | ~v_2038;
assign x_23543 = v_2147 | ~v_2039;
assign x_23544 = v_2147 | ~v_2040;
assign x_23545 = v_2147 | ~v_935;
assign x_23546 = v_2147 | ~v_936;
assign x_23547 = v_2147 | ~v_937;
assign x_23548 = v_2147 | ~v_938;
assign x_23549 = v_2147 | ~v_751;
assign x_23550 = v_2147 | ~v_752;
assign x_23551 = v_2147 | ~v_753;
assign x_23552 = v_2147 | ~v_754;
assign x_23553 = v_2147 | ~v_755;
assign x_23554 = v_2147 | ~v_756;
assign x_23555 = v_2147 | ~v_2099;
assign x_23556 = v_2147 | ~v_2100;
assign x_23557 = v_2147 | ~v_2101;
assign x_23558 = v_2147 | ~v_2102;
assign x_23559 = v_2147 | ~v_2045;
assign x_23560 = v_2147 | ~v_2046;
assign x_23561 = v_2147 | ~v_2047;
assign x_23562 = v_2147 | ~v_2048;
assign x_23563 = v_2147 | ~v_2049;
assign x_23564 = v_2147 | ~v_2050;
assign x_23565 = v_2147 | ~v_1137;
assign x_23566 = v_2147 | ~v_1138;
assign x_23567 = v_2147 | ~v_945;
assign x_23568 = v_2147 | ~v_946;
assign x_23569 = v_2147 | ~v_773;
assign x_23570 = v_2147 | ~v_774;
assign x_23571 = v_2147 | ~v_1139;
assign x_23572 = v_2147 | ~v_1140;
assign x_23573 = v_2147 | ~v_182;
assign x_23574 = v_2147 | ~v_162;
assign x_23575 = v_2147 | ~v_161;
assign x_23576 = v_2147 | ~v_137;
assign x_23577 = v_2147 | ~v_136;
assign x_23578 = v_2147 | ~v_135;
assign x_23579 = v_2147 | ~v_134;
assign x_23580 = v_2147 | ~v_18;
assign x_23581 = v_2147 | ~v_17;
assign x_23582 = v_2147 | ~v_16;
assign x_23583 = v_2147 | ~v_15;
assign x_23584 = v_2147 | ~v_13;
assign x_23585 = ~v_2145 | ~v_2140 | ~v_2135 | v_2146;
assign x_23586 = v_2145 | ~v_2067;
assign x_23587 = v_2145 | ~v_2068;
assign x_23588 = v_2145 | ~v_2069;
assign x_23589 = v_2145 | ~v_2070;
assign x_23590 = v_2145 | ~v_873;
assign x_23591 = v_2145 | ~v_874;
assign x_23592 = v_2145 | ~v_875;
assign x_23593 = v_2145 | ~v_876;
assign x_23594 = v_2145 | ~v_817;
assign x_23595 = v_2145 | ~v_1011;
assign x_23596 = v_2145 | ~v_1012;
assign x_23597 = v_2145 | ~v_820;
assign x_23598 = v_2145 | ~v_1013;
assign x_23599 = v_2145 | ~v_1014;
assign x_23600 = v_2145 | ~v_2093;
assign x_23601 = v_2145 | ~v_2094;
assign x_23602 = v_2145 | ~v_2095;
assign x_23603 = v_2145 | ~v_2096;
assign x_23604 = v_2145 | ~v_2075;
assign x_23605 = v_2145 | ~v_2141;
assign x_23606 = v_2145 | ~v_2142;
assign x_23607 = v_2145 | ~v_2078;
assign x_23608 = v_2145 | ~v_2143;
assign x_23609 = v_2145 | ~v_2144;
assign x_23610 = v_2145 | ~v_885;
assign x_23611 = v_2145 | ~v_1019;
assign x_23612 = v_2145 | ~v_1020;
assign x_23613 = v_2145 | ~v_886;
assign x_23614 = v_2145 | ~v_1021;
assign x_23615 = v_2145 | ~v_1022;
assign x_23616 = v_2145 | ~v_1023;
assign x_23617 = v_2145 | ~v_1024;
assign x_23618 = v_2145 | ~v_184;
assign x_23619 = v_2145 | ~v_181;
assign x_23620 = v_2145 | ~v_171;
assign x_23621 = v_2145 | ~v_169;
assign x_23622 = v_2145 | ~v_149;
assign x_23623 = v_2145 | ~v_148;
assign x_23624 = v_2145 | ~v_147;
assign x_23625 = v_2145 | ~v_103;
assign x_23626 = v_2145 | ~v_102;
assign x_23627 = v_2145 | ~v_101;
assign x_23628 = v_2145 | ~v_99;
assign x_23629 = v_2145 | ~v_94;
assign x_23630 = ~v_130 | ~v_139 | v_2144;
assign x_23631 = ~v_122 | ~v_140 | v_2143;
assign x_23632 = ~v_115 | v_139 | v_2142;
assign x_23633 = ~v_107 | v_140 | v_2141;
assign x_23634 = v_2140 | ~v_2052;
assign x_23635 = v_2140 | ~v_2053;
assign x_23636 = v_2140 | ~v_2054;
assign x_23637 = v_2140 | ~v_2055;
assign x_23638 = v_2140 | ~v_858;
assign x_23639 = v_2140 | ~v_859;
assign x_23640 = v_2140 | ~v_860;
assign x_23641 = v_2140 | ~v_861;
assign x_23642 = v_2140 | ~v_784;
assign x_23643 = v_2140 | ~v_996;
assign x_23644 = v_2140 | ~v_997;
assign x_23645 = v_2140 | ~v_787;
assign x_23646 = v_2140 | ~v_998;
assign x_23647 = v_2140 | ~v_999;
assign x_23648 = v_2140 | ~v_2088;
assign x_23649 = v_2140 | ~v_2089;
assign x_23650 = v_2140 | ~v_2090;
assign x_23651 = v_2140 | ~v_2091;
assign x_23652 = v_2140 | ~v_2060;
assign x_23653 = v_2140 | ~v_2136;
assign x_23654 = v_2140 | ~v_2137;
assign x_23655 = v_2140 | ~v_2063;
assign x_23656 = v_2140 | ~v_2138;
assign x_23657 = v_2140 | ~v_2139;
assign x_23658 = v_2140 | ~v_870;
assign x_23659 = v_2140 | ~v_1004;
assign x_23660 = v_2140 | ~v_1005;
assign x_23661 = v_2140 | ~v_871;
assign x_23662 = v_2140 | ~v_1006;
assign x_23663 = v_2140 | ~v_1007;
assign x_23664 = v_2140 | ~v_1008;
assign x_23665 = v_2140 | ~v_1009;
assign x_23666 = v_2140 | ~v_183;
assign x_23667 = v_2140 | ~v_180;
assign x_23668 = v_2140 | ~v_167;
assign x_23669 = v_2140 | ~v_165;
assign x_23670 = v_2140 | ~v_144;
assign x_23671 = v_2140 | ~v_143;
assign x_23672 = v_2140 | ~v_142;
assign x_23673 = v_2140 | ~v_61;
assign x_23674 = v_2140 | ~v_60;
assign x_23675 = v_2140 | ~v_59;
assign x_23676 = v_2140 | ~v_57;
assign x_23677 = v_2140 | ~v_52;
assign x_23678 = ~v_88 | ~v_139 | v_2139;
assign x_23679 = ~v_80 | ~v_140 | v_2138;
assign x_23680 = ~v_73 | v_139 | v_2137;
assign x_23681 = ~v_65 | v_140 | v_2136;
assign x_23682 = v_2135 | ~v_2037;
assign x_23683 = v_2135 | ~v_2038;
assign x_23684 = v_2135 | ~v_2039;
assign x_23685 = v_2135 | ~v_2040;
assign x_23686 = v_2135 | ~v_843;
assign x_23687 = v_2135 | ~v_844;
assign x_23688 = v_2135 | ~v_845;
assign x_23689 = v_2135 | ~v_846;
assign x_23690 = v_2135 | ~v_751;
assign x_23691 = v_2135 | ~v_981;
assign x_23692 = v_2135 | ~v_982;
assign x_23693 = v_2135 | ~v_754;
assign x_23694 = v_2135 | ~v_983;
assign x_23695 = v_2135 | ~v_984;
assign x_23696 = v_2135 | ~v_2083;
assign x_23697 = v_2135 | ~v_2084;
assign x_23698 = v_2135 | ~v_2085;
assign x_23699 = v_2135 | ~v_2086;
assign x_23700 = v_2135 | ~v_2045;
assign x_23701 = v_2135 | ~v_2131;
assign x_23702 = v_2135 | ~v_2132;
assign x_23703 = v_2135 | ~v_2048;
assign x_23704 = v_2135 | ~v_2133;
assign x_23705 = v_2135 | ~v_2134;
assign x_23706 = v_2135 | ~v_855;
assign x_23707 = v_2135 | ~v_989;
assign x_23708 = v_2135 | ~v_990;
assign x_23709 = v_2135 | ~v_856;
assign x_23710 = v_2135 | ~v_991;
assign x_23711 = v_2135 | ~v_992;
assign x_23712 = v_2135 | ~v_182;
assign x_23713 = v_2135 | ~v_179;
assign x_23714 = v_2135 | ~v_163;
assign x_23715 = v_2135 | ~v_161;
assign x_23716 = v_2135 | ~v_136;
assign x_23717 = v_2135 | ~v_135;
assign x_23718 = v_2135 | ~v_134;
assign x_23719 = v_2135 | ~v_993;
assign x_23720 = v_2135 | ~v_994;
assign x_23721 = v_2135 | ~v_18;
assign x_23722 = v_2135 | ~v_17;
assign x_23723 = v_2135 | ~v_16;
assign x_23724 = v_2135 | ~v_14;
assign x_23725 = v_2135 | ~v_9;
assign x_23726 = ~v_46 | ~v_139 | v_2134;
assign x_23727 = ~v_38 | ~v_140 | v_2133;
assign x_23728 = ~v_31 | v_139 | v_2132;
assign x_23729 = ~v_23 | v_140 | v_2131;
assign x_23730 = ~v_2129 | ~v_2124 | ~v_2119 | v_2130;
assign x_23731 = v_2129 | ~v_2067;
assign x_23732 = v_2129 | ~v_2068;
assign x_23733 = v_2129 | ~v_2069;
assign x_23734 = v_2129 | ~v_2070;
assign x_23735 = v_2129 | ~v_919;
assign x_23736 = v_2129 | ~v_920;
assign x_23737 = v_2129 | ~v_873;
assign x_23738 = v_2129 | ~v_874;
assign x_23739 = v_2129 | ~v_875;
assign x_23740 = v_2129 | ~v_876;
assign x_23741 = v_2129 | ~v_817;
assign x_23742 = v_2129 | ~v_820;
assign x_23743 = v_2129 | ~v_2093;
assign x_23744 = v_2129 | ~v_2094;
assign x_23745 = v_2129 | ~v_2095;
assign x_23746 = v_2129 | ~v_2096;
assign x_23747 = v_2129 | ~v_2125;
assign x_23748 = v_2129 | ~v_2126;
assign x_23749 = v_2129 | ~v_2127;
assign x_23750 = v_2129 | ~v_2128;
assign x_23751 = v_2129 | ~v_2075;
assign x_23752 = v_2129 | ~v_2078;
assign x_23753 = v_2129 | ~v_925;
assign x_23754 = v_2129 | ~v_926;
assign x_23755 = v_2129 | ~v_885;
assign x_23756 = v_2129 | ~v_886;
assign x_23757 = v_2129 | ~v_927;
assign x_23758 = v_2129 | ~v_928;
assign x_23759 = v_2129 | ~v_929;
assign x_23760 = v_2129 | ~v_930;
assign x_23761 = v_2129 | ~v_931;
assign x_23762 = v_2129 | ~v_932;
assign x_23763 = v_2129 | ~v_184;
assign x_23764 = v_2129 | ~v_181;
assign x_23765 = v_2129 | ~v_171;
assign x_23766 = v_2129 | ~v_169;
assign x_23767 = v_2129 | ~v_150;
assign x_23768 = v_2129 | ~v_149;
assign x_23769 = v_2129 | ~v_147;
assign x_23770 = v_2129 | ~v_103;
assign x_23771 = v_2129 | ~v_102;
assign x_23772 = v_2129 | ~v_101;
assign x_23773 = v_2129 | ~v_96;
assign x_23774 = v_2129 | ~v_94;
assign x_23775 = ~v_130 | ~v_141 | v_2128;
assign x_23776 = ~v_122 | ~v_141 | v_2127;
assign x_23777 = ~v_115 | v_141 | v_2126;
assign x_23778 = ~v_107 | v_141 | v_2125;
assign x_23779 = v_2124 | ~v_2052;
assign x_23780 = v_2124 | ~v_2053;
assign x_23781 = v_2124 | ~v_2054;
assign x_23782 = v_2124 | ~v_2055;
assign x_23783 = v_2124 | ~v_904;
assign x_23784 = v_2124 | ~v_905;
assign x_23785 = v_2124 | ~v_858;
assign x_23786 = v_2124 | ~v_859;
assign x_23787 = v_2124 | ~v_860;
assign x_23788 = v_2124 | ~v_861;
assign x_23789 = v_2124 | ~v_784;
assign x_23790 = v_2124 | ~v_787;
assign x_23791 = v_2124 | ~v_2088;
assign x_23792 = v_2124 | ~v_2089;
assign x_23793 = v_2124 | ~v_2090;
assign x_23794 = v_2124 | ~v_2091;
assign x_23795 = v_2124 | ~v_2120;
assign x_23796 = v_2124 | ~v_2121;
assign x_23797 = v_2124 | ~v_2122;
assign x_23798 = v_2124 | ~v_2123;
assign x_23799 = v_2124 | ~v_2060;
assign x_23800 = v_2124 | ~v_2063;
assign x_23801 = v_2124 | ~v_910;
assign x_23802 = v_2124 | ~v_911;
assign x_23803 = v_2124 | ~v_870;
assign x_23804 = v_2124 | ~v_871;
assign x_23805 = v_2124 | ~v_912;
assign x_23806 = v_2124 | ~v_913;
assign x_23807 = v_2124 | ~v_914;
assign x_23808 = v_2124 | ~v_915;
assign x_23809 = v_2124 | ~v_916;
assign x_23810 = v_2124 | ~v_917;
assign x_23811 = v_2124 | ~v_183;
assign x_23812 = v_2124 | ~v_180;
assign x_23813 = v_2124 | ~v_167;
assign x_23814 = v_2124 | ~v_165;
assign x_23815 = v_2124 | ~v_145;
assign x_23816 = v_2124 | ~v_144;
assign x_23817 = v_2124 | ~v_142;
assign x_23818 = v_2124 | ~v_61;
assign x_23819 = v_2124 | ~v_60;
assign x_23820 = v_2124 | ~v_59;
assign x_23821 = v_2124 | ~v_54;
assign x_23822 = v_2124 | ~v_52;
assign x_23823 = ~v_88 | ~v_141 | v_2123;
assign x_23824 = ~v_80 | ~v_141 | v_2122;
assign x_23825 = ~v_73 | v_141 | v_2121;
assign x_23826 = ~v_65 | v_141 | v_2120;
assign x_23827 = v_2119 | ~v_2037;
assign x_23828 = v_2119 | ~v_2038;
assign x_23829 = v_2119 | ~v_2039;
assign x_23830 = v_2119 | ~v_2040;
assign x_23831 = v_2119 | ~v_889;
assign x_23832 = v_2119 | ~v_890;
assign x_23833 = v_2119 | ~v_843;
assign x_23834 = v_2119 | ~v_844;
assign x_23835 = v_2119 | ~v_845;
assign x_23836 = v_2119 | ~v_846;
assign x_23837 = v_2119 | ~v_751;
assign x_23838 = v_2119 | ~v_754;
assign x_23839 = v_2119 | ~v_2083;
assign x_23840 = v_2119 | ~v_2084;
assign x_23841 = v_2119 | ~v_2085;
assign x_23842 = v_2119 | ~v_2086;
assign x_23843 = v_2119 | ~v_2115;
assign x_23844 = v_2119 | ~v_2116;
assign x_23845 = v_2119 | ~v_2117;
assign x_23846 = v_2119 | ~v_2118;
assign x_23847 = v_2119 | ~v_2045;
assign x_23848 = v_2119 | ~v_2048;
assign x_23849 = v_2119 | ~v_895;
assign x_23850 = v_2119 | ~v_896;
assign x_23851 = v_2119 | ~v_855;
assign x_23852 = v_2119 | ~v_856;
assign x_23853 = v_2119 | ~v_897;
assign x_23854 = v_2119 | ~v_898;
assign x_23855 = v_2119 | ~v_899;
assign x_23856 = v_2119 | ~v_900;
assign x_23857 = v_2119 | ~v_901;
assign x_23858 = v_2119 | ~v_902;
assign x_23859 = v_2119 | ~v_182;
assign x_23860 = v_2119 | ~v_179;
assign x_23861 = v_2119 | ~v_163;
assign x_23862 = v_2119 | ~v_161;
assign x_23863 = v_2119 | ~v_137;
assign x_23864 = v_2119 | ~v_136;
assign x_23865 = v_2119 | ~v_134;
assign x_23866 = v_2119 | ~v_18;
assign x_23867 = v_2119 | ~v_17;
assign x_23868 = v_2119 | ~v_16;
assign x_23869 = v_2119 | ~v_11;
assign x_23870 = v_2119 | ~v_9;
assign x_23871 = ~v_46 | ~v_141 | v_2118;
assign x_23872 = ~v_38 | ~v_141 | v_2117;
assign x_23873 = ~v_31 | v_141 | v_2116;
assign x_23874 = ~v_23 | v_141 | v_2115;
assign x_23875 = ~v_2113 | ~v_2108 | ~v_2103 | v_2114;
assign x_23876 = v_2113 | ~v_2067;
assign x_23877 = v_2113 | ~v_2068;
assign x_23878 = v_2113 | ~v_2069;
assign x_23879 = v_2113 | ~v_2070;
assign x_23880 = v_2113 | ~v_965;
assign x_23881 = v_2113 | ~v_966;
assign x_23882 = v_2113 | ~v_967;
assign x_23883 = v_2113 | ~v_968;
assign x_23884 = v_2113 | ~v_873;
assign x_23885 = v_2113 | ~v_874;
assign x_23886 = v_2113 | ~v_875;
assign x_23887 = v_2113 | ~v_876;
assign x_23888 = v_2113 | ~v_817;
assign x_23889 = v_2113 | ~v_820;
assign x_23890 = v_2113 | ~v_2093;
assign x_23891 = v_2113 | ~v_2094;
assign x_23892 = v_2113 | ~v_2095;
assign x_23893 = v_2113 | ~v_2096;
assign x_23894 = v_2113 | ~v_2109;
assign x_23895 = v_2113 | ~v_2110;
assign x_23896 = v_2113 | ~v_2111;
assign x_23897 = v_2113 | ~v_2112;
assign x_23898 = v_2113 | ~v_2075;
assign x_23899 = v_2113 | ~v_2078;
assign x_23900 = v_2113 | ~v_973;
assign x_23901 = v_2113 | ~v_974;
assign x_23902 = v_2113 | ~v_885;
assign x_23903 = v_2113 | ~v_886;
assign x_23904 = v_2113 | ~v_975;
assign x_23905 = v_2113 | ~v_976;
assign x_23906 = v_2113 | ~v_977;
assign x_23907 = v_2113 | ~v_978;
assign x_23908 = v_2113 | ~v_184;
assign x_23909 = v_2113 | ~v_181;
assign x_23910 = v_2113 | ~v_172;
assign x_23911 = v_2113 | ~v_171;
assign x_23912 = v_2113 | ~v_169;
assign x_23913 = v_2113 | ~v_150;
assign x_23914 = v_2113 | ~v_149;
assign x_23915 = v_2113 | ~v_148;
assign x_23916 = v_2113 | ~v_147;
assign x_23917 = v_2113 | ~v_102;
assign x_23918 = v_2113 | ~v_101;
assign x_23919 = v_2113 | ~v_94;
assign x_23920 = ~v_130 | ~v_174 | v_2112;
assign x_23921 = ~v_122 | ~v_173 | v_2111;
assign x_23922 = ~v_115 | v_174 | v_2110;
assign x_23923 = ~v_107 | v_173 | v_2109;
assign x_23924 = v_2108 | ~v_2052;
assign x_23925 = v_2108 | ~v_2053;
assign x_23926 = v_2108 | ~v_2054;
assign x_23927 = v_2108 | ~v_2055;
assign x_23928 = v_2108 | ~v_950;
assign x_23929 = v_2108 | ~v_951;
assign x_23930 = v_2108 | ~v_952;
assign x_23931 = v_2108 | ~v_953;
assign x_23932 = v_2108 | ~v_858;
assign x_23933 = v_2108 | ~v_859;
assign x_23934 = v_2108 | ~v_860;
assign x_23935 = v_2108 | ~v_861;
assign x_23936 = v_2108 | ~v_784;
assign x_23937 = v_2108 | ~v_787;
assign x_23938 = v_2108 | ~v_2088;
assign x_23939 = v_2108 | ~v_2089;
assign x_23940 = v_2108 | ~v_2090;
assign x_23941 = v_2108 | ~v_2091;
assign x_23942 = v_2108 | ~v_2104;
assign x_23943 = v_2108 | ~v_2105;
assign x_23944 = v_2108 | ~v_2106;
assign x_23945 = v_2108 | ~v_2107;
assign x_23946 = v_2108 | ~v_2060;
assign x_23947 = v_2108 | ~v_2063;
assign x_23948 = v_2108 | ~v_958;
assign x_23949 = v_2108 | ~v_959;
assign x_23950 = v_2108 | ~v_870;
assign x_23951 = v_2108 | ~v_871;
assign x_23952 = v_2108 | ~v_960;
assign x_23953 = v_2108 | ~v_961;
assign x_23954 = v_2108 | ~v_962;
assign x_23955 = v_2108 | ~v_963;
assign x_23956 = v_2108 | ~v_183;
assign x_23957 = v_2108 | ~v_180;
assign x_23958 = v_2108 | ~v_168;
assign x_23959 = v_2108 | ~v_167;
assign x_23960 = v_2108 | ~v_165;
assign x_23961 = v_2108 | ~v_145;
assign x_23962 = v_2108 | ~v_144;
assign x_23963 = v_2108 | ~v_143;
assign x_23964 = v_2108 | ~v_142;
assign x_23965 = v_2108 | ~v_60;
assign x_23966 = v_2108 | ~v_59;
assign x_23967 = v_2108 | ~v_52;
assign x_23968 = ~v_88 | ~v_174 | v_2107;
assign x_23969 = ~v_80 | ~v_173 | v_2106;
assign x_23970 = ~v_73 | v_174 | v_2105;
assign x_23971 = ~v_65 | v_173 | v_2104;
assign x_23972 = v_2103 | ~v_2037;
assign x_23973 = v_2103 | ~v_2038;
assign x_23974 = v_2103 | ~v_2039;
assign x_23975 = v_2103 | ~v_2040;
assign x_23976 = v_2103 | ~v_935;
assign x_23977 = v_2103 | ~v_936;
assign x_23978 = v_2103 | ~v_937;
assign x_23979 = v_2103 | ~v_938;
assign x_23980 = v_2103 | ~v_843;
assign x_23981 = v_2103 | ~v_844;
assign x_23982 = v_2103 | ~v_845;
assign x_23983 = v_2103 | ~v_846;
assign x_23984 = v_2103 | ~v_751;
assign x_23985 = v_2103 | ~v_754;
assign x_23986 = v_2103 | ~v_2083;
assign x_23987 = v_2103 | ~v_2084;
assign x_23988 = v_2103 | ~v_2085;
assign x_23989 = v_2103 | ~v_2086;
assign x_23990 = v_2103 | ~v_2099;
assign x_23991 = v_2103 | ~v_2100;
assign x_23992 = v_2103 | ~v_2101;
assign x_23993 = v_2103 | ~v_2102;
assign x_23994 = v_2103 | ~v_2045;
assign x_23995 = v_2103 | ~v_2048;
assign x_23996 = v_2103 | ~v_943;
assign x_23997 = v_2103 | ~v_944;
assign x_23998 = v_2103 | ~v_855;
assign x_23999 = v_2103 | ~v_856;
assign x_24000 = v_2103 | ~v_945;
assign x_24001 = v_2103 | ~v_946;
assign x_24002 = v_2103 | ~v_947;
assign x_24003 = v_2103 | ~v_948;
assign x_24004 = v_2103 | ~v_182;
assign x_24005 = v_2103 | ~v_179;
assign x_24006 = v_2103 | ~v_164;
assign x_24007 = v_2103 | ~v_163;
assign x_24008 = v_2103 | ~v_161;
assign x_24009 = v_2103 | ~v_137;
assign x_24010 = v_2103 | ~v_136;
assign x_24011 = v_2103 | ~v_135;
assign x_24012 = v_2103 | ~v_134;
assign x_24013 = v_2103 | ~v_17;
assign x_24014 = v_2103 | ~v_16;
assign x_24015 = v_2103 | ~v_9;
assign x_24016 = ~v_46 | ~v_174 | v_2102;
assign x_24017 = ~v_38 | ~v_173 | v_2101;
assign x_24018 = ~v_31 | v_174 | v_2100;
assign x_24019 = ~v_23 | v_173 | v_2099;
assign x_24020 = ~v_2097 | ~v_2092 | ~v_2087 | v_2098;
assign x_24021 = v_2097 | ~v_2067;
assign x_24022 = v_2097 | ~v_2068;
assign x_24023 = v_2097 | ~v_2069;
assign x_24024 = v_2097 | ~v_2070;
assign x_24025 = v_2097 | ~v_813;
assign x_24026 = v_2097 | ~v_814;
assign x_24027 = v_2097 | ~v_815;
assign x_24028 = v_2097 | ~v_816;
assign x_24029 = v_2097 | ~v_873;
assign x_24030 = v_2097 | ~v_874;
assign x_24031 = v_2097 | ~v_875;
assign x_24032 = v_2097 | ~v_876;
assign x_24033 = v_2097 | ~v_817;
assign x_24034 = v_2097 | ~v_820;
assign x_24035 = v_2097 | ~v_2093;
assign x_24036 = v_2097 | ~v_2094;
assign x_24037 = v_2097 | ~v_2095;
assign x_24038 = v_2097 | ~v_2096;
assign x_24039 = v_2097 | ~v_2071;
assign x_24040 = v_2097 | ~v_2072;
assign x_24041 = v_2097 | ~v_2073;
assign x_24042 = v_2097 | ~v_2074;
assign x_24043 = v_2097 | ~v_2075;
assign x_24044 = v_2097 | ~v_2078;
assign x_24045 = v_2097 | ~v_881;
assign x_24046 = v_2097 | ~v_882;
assign x_24047 = v_2097 | ~v_883;
assign x_24048 = v_2097 | ~v_884;
assign x_24049 = v_2097 | ~v_885;
assign x_24050 = v_2097 | ~v_886;
assign x_24051 = v_2097 | ~v_837;
assign x_24052 = v_2097 | ~v_838;
assign x_24053 = v_2097 | ~v_184;
assign x_24054 = v_2097 | ~v_181;
assign x_24055 = v_2097 | ~v_171;
assign x_24056 = v_2097 | ~v_169;
assign x_24057 = v_2097 | ~v_160;
assign x_24058 = v_2097 | ~v_150;
assign x_24059 = v_2097 | ~v_148;
assign x_24060 = v_2097 | ~v_103;
assign x_24061 = v_2097 | ~v_102;
assign x_24062 = v_2097 | ~v_97;
assign x_24063 = v_2097 | ~v_95;
assign x_24064 = v_2097 | ~v_94;
assign x_24065 = ~v_127 | ~v_176 | v_2096;
assign x_24066 = ~v_121 | ~v_175 | v_2095;
assign x_24067 = ~v_112 | v_176 | v_2094;
assign x_24068 = ~v_106 | v_175 | v_2093;
assign x_24069 = v_2092 | ~v_2052;
assign x_24070 = v_2092 | ~v_2053;
assign x_24071 = v_2092 | ~v_2054;
assign x_24072 = v_2092 | ~v_2055;
assign x_24073 = v_2092 | ~v_780;
assign x_24074 = v_2092 | ~v_781;
assign x_24075 = v_2092 | ~v_782;
assign x_24076 = v_2092 | ~v_783;
assign x_24077 = v_2092 | ~v_858;
assign x_24078 = v_2092 | ~v_859;
assign x_24079 = v_2092 | ~v_860;
assign x_24080 = v_2092 | ~v_861;
assign x_24081 = v_2092 | ~v_784;
assign x_24082 = v_2092 | ~v_787;
assign x_24083 = v_2092 | ~v_2088;
assign x_24084 = v_2092 | ~v_2089;
assign x_24085 = v_2092 | ~v_2090;
assign x_24086 = v_2092 | ~v_2091;
assign x_24087 = v_2092 | ~v_2056;
assign x_24088 = v_2092 | ~v_2057;
assign x_24089 = v_2092 | ~v_2058;
assign x_24090 = v_2092 | ~v_2059;
assign x_24091 = v_2092 | ~v_2060;
assign x_24092 = v_2092 | ~v_2063;
assign x_24093 = v_2092 | ~v_866;
assign x_24094 = v_2092 | ~v_867;
assign x_24095 = v_2092 | ~v_868;
assign x_24096 = v_2092 | ~v_869;
assign x_24097 = v_2092 | ~v_870;
assign x_24098 = v_2092 | ~v_871;
assign x_24099 = v_2092 | ~v_804;
assign x_24100 = v_2092 | ~v_805;
assign x_24101 = v_2092 | ~v_183;
assign x_24102 = v_2092 | ~v_180;
assign x_24103 = v_2092 | ~v_167;
assign x_24104 = v_2092 | ~v_165;
assign x_24105 = v_2092 | ~v_159;
assign x_24106 = v_2092 | ~v_145;
assign x_24107 = v_2092 | ~v_143;
assign x_24108 = v_2092 | ~v_61;
assign x_24109 = v_2092 | ~v_60;
assign x_24110 = v_2092 | ~v_55;
assign x_24111 = v_2092 | ~v_53;
assign x_24112 = v_2092 | ~v_52;
assign x_24113 = ~v_85 | ~v_176 | v_2091;
assign x_24114 = ~v_79 | ~v_175 | v_2090;
assign x_24115 = ~v_70 | v_176 | v_2089;
assign x_24116 = ~v_64 | v_175 | v_2088;
assign x_24117 = v_2087 | ~v_2037;
assign x_24118 = v_2087 | ~v_2038;
assign x_24119 = v_2087 | ~v_2039;
assign x_24120 = v_2087 | ~v_2040;
assign x_24121 = v_2087 | ~v_747;
assign x_24122 = v_2087 | ~v_748;
assign x_24123 = v_2087 | ~v_749;
assign x_24124 = v_2087 | ~v_750;
assign x_24125 = v_2087 | ~v_843;
assign x_24126 = v_2087 | ~v_844;
assign x_24127 = v_2087 | ~v_845;
assign x_24128 = v_2087 | ~v_846;
assign x_24129 = v_2087 | ~v_751;
assign x_24130 = v_2087 | ~v_754;
assign x_24131 = v_2087 | ~v_2083;
assign x_24132 = v_2087 | ~v_2084;
assign x_24133 = v_2087 | ~v_2085;
assign x_24134 = v_2087 | ~v_2086;
assign x_24135 = v_2087 | ~v_2041;
assign x_24136 = v_2087 | ~v_2042;
assign x_24137 = v_2087 | ~v_2043;
assign x_24138 = v_2087 | ~v_2044;
assign x_24139 = v_2087 | ~v_2045;
assign x_24140 = v_2087 | ~v_2048;
assign x_24141 = v_2087 | ~v_851;
assign x_24142 = v_2087 | ~v_852;
assign x_24143 = v_2087 | ~v_853;
assign x_24144 = v_2087 | ~v_854;
assign x_24145 = v_2087 | ~v_855;
assign x_24146 = v_2087 | ~v_856;
assign x_24147 = v_2087 | ~v_771;
assign x_24148 = v_2087 | ~v_772;
assign x_24149 = v_2087 | ~v_182;
assign x_24150 = v_2087 | ~v_179;
assign x_24151 = v_2087 | ~v_163;
assign x_24152 = v_2087 | ~v_161;
assign x_24153 = v_2087 | ~v_155;
assign x_24154 = v_2087 | ~v_137;
assign x_24155 = v_2087 | ~v_135;
assign x_24156 = v_2087 | ~v_18;
assign x_24157 = v_2087 | ~v_17;
assign x_24158 = v_2087 | ~v_12;
assign x_24159 = v_2087 | ~v_10;
assign x_24160 = v_2087 | ~v_9;
assign x_24161 = ~v_43 | ~v_176 | v_2086;
assign x_24162 = ~v_37 | ~v_175 | v_2085;
assign x_24163 = ~v_28 | v_176 | v_2084;
assign x_24164 = ~v_22 | v_175 | v_2083;
assign x_24165 = ~v_2081 | ~v_2066 | ~v_2051 | v_2082;
assign x_24166 = v_2081 | ~v_2067;
assign x_24167 = v_2081 | ~v_2068;
assign x_24168 = v_2081 | ~v_2069;
assign x_24169 = v_2081 | ~v_2070;
assign x_24170 = v_2081 | ~v_813;
assign x_24171 = v_2081 | ~v_814;
assign x_24172 = v_2081 | ~v_815;
assign x_24173 = v_2081 | ~v_816;
assign x_24174 = v_2081 | ~v_817;
assign x_24175 = v_2081 | ~v_818;
assign x_24176 = v_2081 | ~v_819;
assign x_24177 = v_2081 | ~v_820;
assign x_24178 = v_2081 | ~v_821;
assign x_24179 = v_2081 | ~v_822;
assign x_24180 = v_2081 | ~v_2071;
assign x_24181 = v_2081 | ~v_2072;
assign x_24182 = v_2081 | ~v_2073;
assign x_24183 = v_2081 | ~v_2074;
assign x_24184 = v_2081 | ~v_2075;
assign x_24185 = v_2081 | ~v_2076;
assign x_24186 = v_2081 | ~v_2077;
assign x_24187 = v_2081 | ~v_2078;
assign x_24188 = v_2081 | ~v_2079;
assign x_24189 = v_2081 | ~v_2080;
assign x_24190 = v_2081 | ~v_833;
assign x_24191 = v_2081 | ~v_834;
assign x_24192 = v_2081 | ~v_835;
assign x_24193 = v_2081 | ~v_836;
assign x_24194 = v_2081 | ~v_837;
assign x_24195 = v_2081 | ~v_838;
assign x_24196 = v_2081 | ~v_839;
assign x_24197 = v_2081 | ~v_840;
assign x_24198 = v_2081 | ~v_184;
assign x_24199 = v_2081 | ~v_170;
assign x_24200 = v_2081 | ~v_169;
assign x_24201 = v_2081 | ~v_160;
assign x_24202 = v_2081 | ~v_150;
assign x_24203 = v_2081 | ~v_148;
assign x_24204 = v_2081 | ~v_147;
assign x_24205 = v_2081 | ~v_103;
assign x_24206 = v_2081 | ~v_102;
assign x_24207 = v_2081 | ~v_100;
assign x_24208 = v_2081 | ~v_98;
assign x_24209 = v_2081 | ~v_97;
assign x_24210 = ~v_127 | ~v_139 | v_2080;
assign x_24211 = ~v_121 | ~v_140 | v_2079;
assign x_24212 = ~v_119 | ~v_141 | v_2078;
assign x_24213 = ~v_112 | v_139 | v_2077;
assign x_24214 = ~v_106 | v_140 | v_2076;
assign x_24215 = ~v_104 | v_141 | v_2075;
assign x_24216 = ~v_130 | ~v_176 | v_2074;
assign x_24217 = ~v_122 | ~v_175 | v_2073;
assign x_24218 = ~v_115 | v_176 | v_2072;
assign x_24219 = ~v_107 | v_175 | v_2071;
assign x_24220 = ~v_123 | ~v_176 | v_2070;
assign x_24221 = ~v_120 | ~v_175 | v_2069;
assign x_24222 = ~v_108 | v_176 | v_2068;
assign x_24223 = ~v_105 | v_175 | v_2067;
assign x_24224 = v_2066 | ~v_2052;
assign x_24225 = v_2066 | ~v_2053;
assign x_24226 = v_2066 | ~v_2054;
assign x_24227 = v_2066 | ~v_2055;
assign x_24228 = v_2066 | ~v_780;
assign x_24229 = v_2066 | ~v_781;
assign x_24230 = v_2066 | ~v_782;
assign x_24231 = v_2066 | ~v_783;
assign x_24232 = v_2066 | ~v_784;
assign x_24233 = v_2066 | ~v_785;
assign x_24234 = v_2066 | ~v_786;
assign x_24235 = v_2066 | ~v_787;
assign x_24236 = v_2066 | ~v_788;
assign x_24237 = v_2066 | ~v_789;
assign x_24238 = v_2066 | ~v_2056;
assign x_24239 = v_2066 | ~v_2057;
assign x_24240 = v_2066 | ~v_2058;
assign x_24241 = v_2066 | ~v_2059;
assign x_24242 = v_2066 | ~v_2060;
assign x_24243 = v_2066 | ~v_2061;
assign x_24244 = v_2066 | ~v_2062;
assign x_24245 = v_2066 | ~v_2063;
assign x_24246 = v_2066 | ~v_2064;
assign x_24247 = v_2066 | ~v_2065;
assign x_24248 = v_2066 | ~v_800;
assign x_24249 = v_2066 | ~v_801;
assign x_24250 = v_2066 | ~v_802;
assign x_24251 = v_2066 | ~v_803;
assign x_24252 = v_2066 | ~v_804;
assign x_24253 = v_2066 | ~v_805;
assign x_24254 = v_2066 | ~v_806;
assign x_24255 = v_2066 | ~v_807;
assign x_24256 = v_2066 | ~v_183;
assign x_24257 = v_2066 | ~v_166;
assign x_24258 = v_2066 | ~v_165;
assign x_24259 = v_2066 | ~v_159;
assign x_24260 = v_2066 | ~v_145;
assign x_24261 = v_2066 | ~v_143;
assign x_24262 = v_2066 | ~v_142;
assign x_24263 = v_2066 | ~v_61;
assign x_24264 = v_2066 | ~v_60;
assign x_24265 = v_2066 | ~v_58;
assign x_24266 = v_2066 | ~v_56;
assign x_24267 = v_2066 | ~v_55;
assign x_24268 = ~v_85 | ~v_139 | v_2065;
assign x_24269 = ~v_79 | ~v_140 | v_2064;
assign x_24270 = ~v_77 | ~v_141 | v_2063;
assign x_24271 = ~v_70 | v_139 | v_2062;
assign x_24272 = ~v_64 | v_140 | v_2061;
assign x_24273 = ~v_62 | v_141 | v_2060;
assign x_24274 = ~v_88 | ~v_176 | v_2059;
assign x_24275 = ~v_80 | ~v_175 | v_2058;
assign x_24276 = ~v_73 | v_176 | v_2057;
assign x_24277 = ~v_65 | v_175 | v_2056;
assign x_24278 = ~v_81 | ~v_176 | v_2055;
assign x_24279 = ~v_78 | ~v_175 | v_2054;
assign x_24280 = ~v_66 | v_176 | v_2053;
assign x_24281 = ~v_63 | v_175 | v_2052;
assign x_24282 = v_2051 | ~v_2037;
assign x_24283 = v_2051 | ~v_2038;
assign x_24284 = v_2051 | ~v_2039;
assign x_24285 = v_2051 | ~v_2040;
assign x_24286 = v_2051 | ~v_747;
assign x_24287 = v_2051 | ~v_748;
assign x_24288 = v_2051 | ~v_749;
assign x_24289 = v_2051 | ~v_750;
assign x_24290 = v_2051 | ~v_751;
assign x_24291 = v_2051 | ~v_752;
assign x_24292 = v_2051 | ~v_753;
assign x_24293 = v_2051 | ~v_754;
assign x_24294 = v_2051 | ~v_755;
assign x_24295 = v_2051 | ~v_756;
assign x_24296 = v_2051 | ~v_2041;
assign x_24297 = v_2051 | ~v_2042;
assign x_24298 = v_2051 | ~v_2043;
assign x_24299 = v_2051 | ~v_2044;
assign x_24300 = v_2051 | ~v_2045;
assign x_24301 = v_2051 | ~v_2046;
assign x_24302 = v_2051 | ~v_2047;
assign x_24303 = v_2051 | ~v_2048;
assign x_24304 = v_2051 | ~v_2049;
assign x_24305 = v_2051 | ~v_2050;
assign x_24306 = v_2051 | ~v_767;
assign x_24307 = v_2051 | ~v_768;
assign x_24308 = v_2051 | ~v_769;
assign x_24309 = v_2051 | ~v_770;
assign x_24310 = v_2051 | ~v_771;
assign x_24311 = v_2051 | ~v_772;
assign x_24312 = v_2051 | ~v_773;
assign x_24313 = v_2051 | ~v_774;
assign x_24314 = v_2051 | ~v_182;
assign x_24315 = v_2051 | ~v_162;
assign x_24316 = v_2051 | ~v_161;
assign x_24317 = v_2051 | ~v_155;
assign x_24318 = v_2051 | ~v_137;
assign x_24319 = v_2051 | ~v_135;
assign x_24320 = v_2051 | ~v_134;
assign x_24321 = v_2051 | ~v_18;
assign x_24322 = v_2051 | ~v_17;
assign x_24323 = v_2051 | ~v_15;
assign x_24324 = v_2051 | ~v_13;
assign x_24325 = v_2051 | ~v_12;
assign x_24326 = ~v_43 | ~v_139 | v_2050;
assign x_24327 = ~v_37 | ~v_140 | v_2049;
assign x_24328 = ~v_35 | ~v_141 | v_2048;
assign x_24329 = ~v_28 | v_139 | v_2047;
assign x_24330 = ~v_22 | v_140 | v_2046;
assign x_24331 = ~v_20 | v_141 | v_2045;
assign x_24332 = ~v_46 | ~v_176 | v_2044;
assign x_24333 = ~v_38 | ~v_175 | v_2043;
assign x_24334 = ~v_31 | v_176 | v_2042;
assign x_24335 = ~v_23 | v_175 | v_2041;
assign x_24336 = ~v_39 | ~v_176 | v_2040;
assign x_24337 = ~v_36 | ~v_175 | v_2039;
assign x_24338 = ~v_24 | v_176 | v_2038;
assign x_24339 = ~v_21 | v_175 | v_2037;
assign x_24340 = v_2036 | ~v_739;
assign x_24341 = v_2036 | ~v_728;
assign x_24342 = v_2035 | ~v_2034;
assign x_24343 = v_2035 | ~v_731;
assign x_24344 = v_177 | v_178 | ~v_742 | ~v_741 | v_2034;
assign x_24345 = ~v_725 | ~v_724 | ~v_723 | ~v_722 | ~v_2032 | ~v_2028 | ~v_2024 | ~v_2020 | ~v_2016 | ~v_2000 | ~v_1996 | ~v_1992 | ~v_1988 | ~v_1984 | ~v_1968 | ~v_1964 | ~v_1948 | ~v_1932 | ~v_1916 | ~v_1900 | ~v_1854 | v_2033;
assign x_24346 = v_2032 | ~v_2029;
assign x_24347 = v_2032 | ~v_2030;
assign x_24348 = v_2032 | ~v_2031;
assign x_24349 = v_98 | v_103 | v_101 | v_100 | v_95 | v_99 | v_102 | ~v_719 | ~v_718 | v_170 | v_169 | v_149 | v_148 | v_184 | ~v_483 | ~v_717 | ~v_299 | ~v_482 | ~v_716 | ~v_298 | ~v_1962 | ~v_1898 | ~v_1961 | ~v_1897 | ~v_1896 | ~v_1960 | ~v_1895 | ~v_1959 | ~v_1894 | ~v_1893 | ~v_473 | ~v_281 | ~v_472 | ~v_280 | ~v_279 | ~v_471 | ~v_278 | ~v_470 | ~v_277 | ~v_276 | ~v_1888 | ~v_1887 | ~v_1886 | ~v_1885 | v_2031;
assign x_24350 = v_53 | v_56 | v_61 | v_60 | v_59 | v_58 | v_57 | ~v_714 | ~v_713 | v_144 | v_143 | v_166 | v_165 | v_183 | ~v_266 | ~v_468 | ~v_712 | ~v_467 | ~v_711 | ~v_265 | ~v_1957 | ~v_1883 | ~v_1956 | ~v_1882 | ~v_1881 | ~v_1955 | ~v_1880 | ~v_1954 | ~v_1879 | ~v_1878 | ~v_458 | ~v_248 | ~v_457 | ~v_247 | ~v_246 | ~v_456 | ~v_245 | ~v_455 | ~v_244 | ~v_243 | ~v_1873 | ~v_1872 | ~v_1871 | ~v_1870 | v_2030;
assign x_24351 = v_13 | v_18 | v_17 | v_16 | v_15 | v_14 | v_10 | ~v_453 | ~v_709 | ~v_452 | ~v_708 | v_136 | v_135 | ~v_707 | ~v_706 | v_162 | v_161 | v_182 | ~v_233 | ~v_232 | ~v_1952 | ~v_1868 | ~v_1951 | ~v_1867 | ~v_1866 | ~v_1950 | ~v_1865 | ~v_1949 | ~v_1864 | ~v_1863 | ~v_443 | ~v_215 | ~v_442 | ~v_214 | ~v_213 | ~v_441 | ~v_212 | ~v_440 | ~v_211 | ~v_210 | ~v_1858 | ~v_1857 | ~v_1856 | ~v_1855 | v_2029;
assign x_24352 = v_2028 | ~v_2025;
assign x_24353 = v_2028 | ~v_2026;
assign x_24354 = v_2028 | ~v_2027;
assign x_24355 = v_101 | v_100 | v_99 | v_93 | v_102 | v_172 | v_171 | v_170 | v_149 | v_148 | v_147 | v_184 | ~v_483 | ~v_482 | ~v_593 | ~v_592 | ~v_545 | ~v_591 | ~v_590 | ~v_544 | ~v_1962 | ~v_1961 | ~v_1896 | ~v_1960 | ~v_1959 | ~v_1893 | ~v_2014 | ~v_2013 | ~v_2012 | ~v_2011 | ~v_473 | ~v_472 | ~v_279 | ~v_471 | ~v_470 | ~v_276 | ~v_535 | ~v_534 | ~v_533 | ~v_532 | ~v_1888 | ~v_1887 | ~v_1886 | ~v_1885 | v_2027;
assign x_24356 = v_51 | v_60 | v_59 | v_58 | v_57 | v_144 | v_143 | v_142 | v_168 | v_167 | v_166 | v_183 | ~v_468 | ~v_467 | ~v_588 | ~v_587 | ~v_530 | ~v_586 | ~v_585 | ~v_529 | ~v_1957 | ~v_1956 | ~v_1881 | ~v_1955 | ~v_1954 | ~v_1878 | ~v_2009 | ~v_2008 | ~v_2007 | ~v_2006 | ~v_458 | ~v_457 | ~v_246 | ~v_456 | ~v_455 | ~v_243 | ~v_520 | ~v_519 | ~v_518 | ~v_517 | ~v_1873 | ~v_1872 | ~v_1871 | ~v_1870 | v_2026;
assign x_24357 = v_17 | v_16 | v_8 | v_15 | v_14 | ~v_453 | ~v_452 | v_136 | v_135 | v_134 | v_164 | v_163 | v_162 | v_182 | ~v_583 | ~v_582 | ~v_515 | ~v_581 | ~v_580 | ~v_514 | ~v_1952 | ~v_1951 | ~v_1866 | ~v_1950 | ~v_1949 | ~v_1863 | ~v_2004 | ~v_2003 | ~v_2002 | ~v_2001 | ~v_443 | ~v_442 | ~v_213 | ~v_441 | ~v_440 | ~v_210 | ~v_505 | ~v_504 | ~v_503 | ~v_502 | ~v_1858 | ~v_1857 | ~v_1856 | ~v_1855 | v_2025;
assign x_24358 = v_2024 | ~v_2021;
assign x_24359 = v_2024 | ~v_2022;
assign x_24360 = v_2024 | ~v_2023;
assign x_24361 = v_103 | v_101 | v_96 | v_100 | v_95 | v_93 | v_102 | v_171 | v_170 | v_150 | v_149 | v_184 | ~v_389 | ~v_388 | ~v_545 | ~v_544 | ~v_561 | ~v_560 | ~v_559 | ~v_558 | ~v_387 | ~v_386 | ~v_1896 | ~v_1893 | ~v_2014 | ~v_2013 | ~v_2012 | ~v_2011 | ~v_1946 | ~v_1945 | ~v_1944 | ~v_1943 | ~v_279 | ~v_276 | ~v_379 | ~v_378 | ~v_535 | ~v_534 | ~v_533 | ~v_532 | ~v_1888 | ~v_1887 | ~v_1886 | ~v_1885 | v_2023;
assign x_24362 = v_54 | v_53 | v_61 | v_51 | v_60 | v_59 | v_58 | v_144 | v_145 | v_167 | v_166 | v_183 | ~v_374 | ~v_373 | ~v_530 | ~v_529 | ~v_556 | ~v_555 | ~v_554 | ~v_553 | ~v_372 | ~v_371 | ~v_1881 | ~v_1878 | ~v_2009 | ~v_2008 | ~v_2007 | ~v_2006 | ~v_1941 | ~v_1940 | ~v_1939 | ~v_1938 | ~v_246 | ~v_243 | ~v_364 | ~v_363 | ~v_520 | ~v_519 | ~v_518 | ~v_517 | ~v_1873 | ~v_1872 | ~v_1871 | ~v_1870 | v_2022;
assign x_24363 = v_18 | v_17 | v_16 | v_8 | v_15 | v_11 | v_10 | v_136 | v_137 | v_163 | v_162 | v_182 | ~v_359 | ~v_358 | ~v_515 | ~v_514 | ~v_551 | ~v_550 | ~v_549 | ~v_548 | ~v_357 | ~v_356 | ~v_1866 | ~v_1863 | ~v_2004 | ~v_2003 | ~v_2002 | ~v_2001 | ~v_1936 | ~v_1935 | ~v_1934 | ~v_1933 | ~v_213 | ~v_210 | ~v_349 | ~v_348 | ~v_505 | ~v_504 | ~v_503 | ~v_502 | ~v_1858 | ~v_1857 | ~v_1856 | ~v_1855 | v_2021;
assign x_24364 = v_2020 | ~v_2017;
assign x_24365 = v_2020 | ~v_2018;
assign x_24366 = v_2020 | ~v_2019;
assign x_24367 = v_103 | v_101 | v_100 | v_93 | v_151 | v_171 | v_170 | v_150 | v_149 | v_148 | v_147 | v_184 | ~v_577 | ~v_576 | ~v_545 | ~v_544 | ~v_575 | ~v_574 | ~v_435 | ~v_434 | ~v_1896 | ~v_1893 | ~v_2014 | ~v_2013 | ~v_2012 | ~v_2011 | ~v_1930 | ~v_1929 | ~v_1928 | ~v_1927 | ~v_279 | ~v_276 | ~v_427 | ~v_426 | ~v_425 | ~v_424 | ~v_535 | ~v_534 | ~v_533 | ~v_532 | ~v_1888 | ~v_1887 | ~v_1886 | ~v_1885 | v_2019;
assign x_24368 = v_61 | v_51 | v_59 | v_58 | v_144 | v_145 | v_143 | v_142 | v_167 | v_166 | v_146 | v_183 | ~v_572 | ~v_571 | ~v_530 | ~v_529 | ~v_570 | ~v_569 | ~v_420 | ~v_419 | ~v_1881 | ~v_1878 | ~v_2009 | ~v_2008 | ~v_2007 | ~v_2006 | ~v_1925 | ~v_1924 | ~v_1923 | ~v_1922 | ~v_246 | ~v_243 | ~v_412 | ~v_411 | ~v_410 | ~v_409 | ~v_520 | ~v_519 | ~v_518 | ~v_517 | ~v_1873 | ~v_1872 | ~v_1871 | ~v_1870 | v_2018;
assign x_24369 = v_18 | v_16 | v_8 | v_15 | v_136 | v_135 | v_134 | v_137 | v_138 | v_163 | v_162 | v_182 | ~v_567 | ~v_566 | ~v_515 | ~v_514 | ~v_565 | ~v_564 | ~v_405 | ~v_404 | ~v_1866 | ~v_1863 | ~v_2004 | ~v_2003 | ~v_2002 | ~v_2001 | ~v_1920 | ~v_1919 | ~v_1918 | ~v_1917 | ~v_213 | ~v_210 | ~v_397 | ~v_396 | ~v_395 | ~v_394 | ~v_505 | ~v_504 | ~v_503 | ~v_502 | ~v_1858 | ~v_1857 | ~v_1856 | ~v_1855 | v_2017;
assign x_24370 = v_2016 | ~v_2005;
assign x_24371 = v_2016 | ~v_2010;
assign x_24372 = v_2016 | ~v_2015;
assign x_24373 = v_103 | v_97 | v_100 | v_93 | v_102 | v_171 | v_170 | v_160 | v_150 | v_148 | v_147 | v_184 | ~v_545 | ~v_544 | ~v_543 | ~v_542 | ~v_541 | ~v_540 | ~v_297 | ~v_296 | ~v_1896 | ~v_1893 | ~v_2014 | ~v_2013 | ~v_2012 | ~v_2011 | ~v_1892 | ~v_1891 | ~v_1890 | ~v_1889 | ~v_279 | ~v_276 | ~v_275 | ~v_274 | ~v_273 | ~v_272 | ~v_535 | ~v_534 | ~v_533 | ~v_532 | ~v_1888 | ~v_1887 | ~v_1886 | ~v_1885 | v_2015;
assign x_24374 = v_2014 | v_141;
assign x_24375 = v_2014 | v_127;
assign x_24376 = v_2013 | v_141;
assign x_24377 = v_2013 | v_121;
assign x_24378 = v_2012 | ~v_141;
assign x_24379 = v_2012 | v_112;
assign x_24380 = v_2011 | ~v_141;
assign x_24381 = v_2011 | v_106;
assign x_24382 = v_55 | v_61 | v_51 | v_60 | v_58 | v_159 | v_145 | v_143 | v_142 | v_167 | v_166 | v_183 | ~v_530 | ~v_529 | ~v_528 | ~v_527 | ~v_526 | ~v_525 | ~v_264 | ~v_263 | ~v_1881 | ~v_1878 | ~v_2009 | ~v_2008 | ~v_2007 | ~v_2006 | ~v_1877 | ~v_1876 | ~v_1875 | ~v_1874 | ~v_246 | ~v_243 | ~v_242 | ~v_241 | ~v_240 | ~v_239 | ~v_520 | ~v_519 | ~v_518 | ~v_517 | ~v_1873 | ~v_1872 | ~v_1871 | ~v_1870 | v_2010;
assign x_24383 = v_2009 | v_141;
assign x_24384 = v_2009 | v_85;
assign x_24385 = v_2008 | v_141;
assign x_24386 = v_2008 | v_79;
assign x_24387 = v_2007 | ~v_141;
assign x_24388 = v_2007 | v_70;
assign x_24389 = v_2006 | ~v_141;
assign x_24390 = v_2006 | v_64;
assign x_24391 = v_18 | v_17 | v_8 | v_15 | v_12 | v_135 | v_134 | v_137 | v_163 | v_162 | v_155 | v_182 | ~v_515 | ~v_514 | ~v_513 | ~v_512 | ~v_511 | ~v_510 | ~v_231 | ~v_230 | ~v_1866 | ~v_1863 | ~v_2004 | ~v_2003 | ~v_2002 | ~v_2001 | ~v_1862 | ~v_1861 | ~v_1860 | ~v_1859 | ~v_213 | ~v_210 | ~v_209 | ~v_208 | ~v_207 | ~v_206 | ~v_505 | ~v_504 | ~v_503 | ~v_502 | ~v_1858 | ~v_1857 | ~v_1856 | ~v_1855 | v_2005;
assign x_24392 = v_2004 | v_141;
assign x_24393 = v_2004 | v_43;
assign x_24394 = v_2003 | v_141;
assign x_24395 = v_2003 | v_37;
assign x_24396 = v_2002 | ~v_141;
assign x_24397 = v_2002 | v_28;
assign x_24398 = v_2001 | ~v_141;
assign x_24399 = v_2001 | v_22;
assign x_24400 = v_2000 | ~v_1997;
assign x_24401 = v_2000 | ~v_1998;
assign x_24402 = v_2000 | ~v_1999;
assign x_24403 = v_98 | v_103 | v_101 | v_96 | v_100 | v_151 | v_170 | v_169 | v_150 | v_149 | v_147 | v_184 | ~v_389 | ~v_388 | ~v_299 | ~v_298 | ~v_387 | ~v_386 | ~v_499 | ~v_498 | ~v_497 | ~v_496 | ~v_1898 | ~v_1897 | ~v_1896 | ~v_1895 | ~v_1894 | ~v_1893 | ~v_1946 | ~v_1945 | ~v_1944 | ~v_1943 | ~v_281 | ~v_280 | ~v_279 | ~v_278 | ~v_277 | ~v_276 | ~v_379 | ~v_378 | ~v_1888 | ~v_1887 | ~v_1886 | ~v_1885 | v_1999;
assign x_24404 = v_54 | v_56 | v_61 | v_59 | v_58 | v_144 | v_145 | v_142 | v_166 | v_165 | v_146 | v_183 | ~v_374 | ~v_373 | ~v_266 | ~v_265 | ~v_372 | ~v_371 | ~v_494 | ~v_493 | ~v_492 | ~v_491 | ~v_1883 | ~v_1882 | ~v_1881 | ~v_1880 | ~v_1879 | ~v_1878 | ~v_1941 | ~v_1940 | ~v_1939 | ~v_1938 | ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_244 | ~v_243 | ~v_364 | ~v_363 | ~v_1873 | ~v_1872 | ~v_1871 | ~v_1870 | v_1998;
assign x_24405 = v_13 | v_18 | v_16 | v_15 | v_11 | v_136 | v_134 | v_137 | v_138 | v_162 | v_161 | v_182 | ~v_359 | ~v_358 | ~v_233 | ~v_232 | ~v_357 | ~v_356 | ~v_489 | ~v_488 | ~v_487 | ~v_486 | ~v_1868 | ~v_1867 | ~v_1866 | ~v_1865 | ~v_1864 | ~v_1863 | ~v_1936 | ~v_1935 | ~v_1934 | ~v_1933 | ~v_215 | ~v_214 | ~v_213 | ~v_212 | ~v_211 | ~v_210 | ~v_349 | ~v_348 | ~v_1858 | ~v_1857 | ~v_1856 | ~v_1855 | v_1997;
assign x_24406 = v_1996 | ~v_1993;
assign x_24407 = v_1996 | ~v_1994;
assign x_24408 = v_1996 | ~v_1995;
assign x_24409 = v_103 | v_101 | v_100 | v_99 | v_102 | v_171 | v_170 | v_169 | v_149 | v_148 | v_147 | v_184 | ~v_703 | ~v_702 | ~v_483 | ~v_482 | ~v_701 | ~v_653 | ~v_700 | ~v_652 | ~v_1962 | ~v_1961 | ~v_1896 | ~v_1960 | ~v_1959 | ~v_1893 | ~v_1982 | ~v_1981 | ~v_1980 | ~v_1979 | ~v_473 | ~v_472 | ~v_279 | ~v_471 | ~v_470 | ~v_276 | ~v_645 | ~v_644 | ~v_643 | ~v_642 | ~v_1888 | ~v_1887 | ~v_1886 | ~v_1885 | v_1995;
assign x_24410 = v_61 | v_60 | v_59 | v_58 | v_57 | v_144 | v_143 | v_142 | v_167 | v_166 | v_165 | v_183 | ~v_698 | ~v_697 | ~v_468 | ~v_467 | ~v_696 | ~v_638 | ~v_695 | ~v_637 | ~v_1957 | ~v_1956 | ~v_1881 | ~v_1955 | ~v_1954 | ~v_1878 | ~v_1977 | ~v_1976 | ~v_1975 | ~v_1974 | ~v_458 | ~v_457 | ~v_246 | ~v_456 | ~v_455 | ~v_243 | ~v_630 | ~v_629 | ~v_628 | ~v_627 | ~v_1873 | ~v_1872 | ~v_1871 | ~v_1870 | v_1994;
assign x_24411 = v_18 | v_17 | v_16 | v_15 | v_14 | ~v_453 | ~v_452 | v_136 | v_135 | v_134 | v_163 | v_162 | v_161 | v_182 | ~v_693 | ~v_692 | ~v_691 | ~v_623 | ~v_690 | ~v_622 | ~v_1952 | ~v_1951 | ~v_1866 | ~v_1950 | ~v_1949 | ~v_1863 | ~v_1972 | ~v_1971 | ~v_1970 | ~v_1969 | ~v_443 | ~v_442 | ~v_213 | ~v_441 | ~v_440 | ~v_210 | ~v_615 | ~v_614 | ~v_613 | ~v_612 | ~v_1858 | ~v_1857 | ~v_1856 | ~v_1855 | v_1993;
assign x_24412 = v_1992 | ~v_1989;
assign x_24413 = v_1992 | ~v_1990;
assign x_24414 = v_1992 | ~v_1991;
assign x_24415 = v_101 | v_96 | v_100 | v_102 | v_172 | v_171 | v_170 | v_169 | v_150 | v_149 | v_147 | v_184 | ~v_389 | ~v_388 | ~v_671 | ~v_670 | ~v_387 | ~v_386 | ~v_653 | ~v_652 | ~v_669 | ~v_668 | ~v_1896 | ~v_1893 | ~v_1946 | ~v_1945 | ~v_1944 | ~v_1943 | ~v_1982 | ~v_1981 | ~v_1980 | ~v_1979 | ~v_279 | ~v_276 | ~v_379 | ~v_378 | ~v_645 | ~v_644 | ~v_643 | ~v_642 | ~v_1888 | ~v_1887 | ~v_1886 | ~v_1885 | v_1991;
assign x_24416 = v_54 | v_60 | v_59 | v_58 | v_144 | v_145 | v_142 | v_168 | v_167 | v_166 | v_165 | v_183 | ~v_374 | ~v_373 | ~v_666 | ~v_665 | ~v_372 | ~v_371 | ~v_638 | ~v_637 | ~v_664 | ~v_663 | ~v_1881 | ~v_1878 | ~v_1941 | ~v_1940 | ~v_1939 | ~v_1938 | ~v_1977 | ~v_1976 | ~v_1975 | ~v_1974 | ~v_246 | ~v_243 | ~v_364 | ~v_363 | ~v_630 | ~v_629 | ~v_628 | ~v_627 | ~v_1873 | ~v_1872 | ~v_1871 | ~v_1870 | v_1990;
assign x_24417 = v_17 | v_16 | v_15 | v_11 | v_136 | v_134 | v_137 | v_164 | v_163 | v_162 | v_161 | v_182 | ~v_359 | ~v_358 | ~v_661 | ~v_660 | ~v_357 | ~v_356 | ~v_623 | ~v_622 | ~v_659 | ~v_658 | ~v_1866 | ~v_1863 | ~v_1936 | ~v_1935 | ~v_1934 | ~v_1933 | ~v_1972 | ~v_1971 | ~v_1970 | ~v_1969 | ~v_213 | ~v_210 | ~v_349 | ~v_348 | ~v_615 | ~v_614 | ~v_613 | ~v_612 | ~v_1858 | ~v_1857 | ~v_1856 | ~v_1855 | v_1989;
assign x_24418 = v_1988 | ~v_1985;
assign x_24419 = v_1988 | ~v_1986;
assign x_24420 = v_1988 | ~v_1987;
assign x_24421 = v_103 | v_101 | v_100 | v_95 | v_102 | v_171 | v_170 | v_169 | v_150 | v_149 | v_148 | v_184 | ~v_435 | ~v_434 | ~v_653 | ~v_652 | ~v_687 | ~v_686 | ~v_685 | ~v_684 | ~v_1896 | ~v_1893 | ~v_1930 | ~v_1929 | ~v_1928 | ~v_1927 | ~v_1982 | ~v_1981 | ~v_1980 | ~v_1979 | ~v_279 | ~v_276 | ~v_427 | ~v_426 | ~v_425 | ~v_424 | ~v_645 | ~v_644 | ~v_643 | ~v_642 | ~v_1888 | ~v_1887 | ~v_1886 | ~v_1885 | v_1987;
assign x_24422 = v_53 | v_61 | v_60 | v_59 | v_58 | v_144 | v_145 | v_143 | v_167 | v_166 | v_165 | v_183 | ~v_420 | ~v_419 | ~v_638 | ~v_637 | ~v_682 | ~v_681 | ~v_680 | ~v_679 | ~v_1881 | ~v_1878 | ~v_1925 | ~v_1924 | ~v_1923 | ~v_1922 | ~v_1977 | ~v_1976 | ~v_1975 | ~v_1974 | ~v_246 | ~v_243 | ~v_412 | ~v_411 | ~v_410 | ~v_409 | ~v_630 | ~v_629 | ~v_628 | ~v_627 | ~v_1873 | ~v_1872 | ~v_1871 | ~v_1870 | v_1986;
assign x_24423 = v_18 | v_17 | v_16 | v_15 | v_10 | v_136 | v_135 | v_137 | v_163 | v_162 | v_161 | v_182 | ~v_405 | ~v_404 | ~v_623 | ~v_622 | ~v_677 | ~v_676 | ~v_675 | ~v_674 | ~v_1866 | ~v_1863 | ~v_1920 | ~v_1919 | ~v_1918 | ~v_1917 | ~v_1972 | ~v_1971 | ~v_1970 | ~v_1969 | ~v_213 | ~v_210 | ~v_397 | ~v_396 | ~v_395 | ~v_394 | ~v_615 | ~v_614 | ~v_613 | ~v_612 | ~v_1858 | ~v_1857 | ~v_1856 | ~v_1855 | v_1985;
assign x_24424 = v_1984 | ~v_1973;
assign x_24425 = v_1984 | ~v_1978;
assign x_24426 = v_1984 | ~v_1983;
assign x_24427 = v_103 | v_97 | v_100 | v_151 | v_171 | v_170 | v_169 | v_160 | v_150 | v_148 | v_147 | v_184 | ~v_655 | ~v_654 | ~v_297 | ~v_296 | ~v_653 | ~v_652 | ~v_651 | ~v_650 | ~v_1896 | ~v_1893 | ~v_1892 | ~v_1891 | ~v_1890 | ~v_1889 | ~v_1982 | ~v_1981 | ~v_1980 | ~v_1979 | ~v_279 | ~v_276 | ~v_275 | ~v_274 | ~v_273 | ~v_272 | ~v_645 | ~v_644 | ~v_643 | ~v_642 | ~v_1888 | ~v_1887 | ~v_1886 | ~v_1885 | v_1983;
assign x_24428 = v_1982 | v_174;
assign x_24429 = v_1982 | v_127;
assign x_24430 = v_1981 | v_173;
assign x_24431 = v_1981 | v_121;
assign x_24432 = v_1980 | ~v_174;
assign x_24433 = v_1980 | v_112;
assign x_24434 = v_1979 | ~v_173;
assign x_24435 = v_1979 | v_106;
assign x_24436 = v_55 | v_61 | v_58 | v_159 | v_145 | v_143 | v_142 | v_167 | v_166 | v_165 | v_146 | v_183 | ~v_640 | ~v_639 | ~v_264 | ~v_263 | ~v_638 | ~v_637 | ~v_636 | ~v_635 | ~v_1881 | ~v_1878 | ~v_1877 | ~v_1876 | ~v_1875 | ~v_1874 | ~v_1977 | ~v_1976 | ~v_1975 | ~v_1974 | ~v_246 | ~v_243 | ~v_242 | ~v_241 | ~v_240 | ~v_239 | ~v_630 | ~v_629 | ~v_628 | ~v_627 | ~v_1873 | ~v_1872 | ~v_1871 | ~v_1870 | v_1978;
assign x_24437 = v_1977 | v_174;
assign x_24438 = v_1977 | v_85;
assign x_24439 = v_1976 | v_173;
assign x_24440 = v_1976 | v_79;
assign x_24441 = v_1975 | ~v_174;
assign x_24442 = v_1975 | v_70;
assign x_24443 = v_1974 | ~v_173;
assign x_24444 = v_1974 | v_64;
assign x_24445 = v_18 | v_15 | v_12 | v_135 | v_134 | v_137 | v_138 | v_163 | v_162 | v_161 | v_155 | v_182 | ~v_625 | ~v_624 | ~v_231 | ~v_230 | ~v_623 | ~v_622 | ~v_621 | ~v_620 | ~v_1866 | ~v_1863 | ~v_1862 | ~v_1861 | ~v_1860 | ~v_1859 | ~v_1972 | ~v_1971 | ~v_1970 | ~v_1969 | ~v_213 | ~v_210 | ~v_209 | ~v_208 | ~v_207 | ~v_206 | ~v_615 | ~v_614 | ~v_613 | ~v_612 | ~v_1858 | ~v_1857 | ~v_1856 | ~v_1855 | v_1973;
assign x_24446 = v_1972 | v_174;
assign x_24447 = v_1972 | v_43;
assign x_24448 = v_1971 | v_173;
assign x_24449 = v_1971 | v_37;
assign x_24450 = v_1970 | ~v_174;
assign x_24451 = v_1970 | v_28;
assign x_24452 = v_1969 | ~v_173;
assign x_24453 = v_1969 | v_22;
assign x_24454 = v_1968 | ~v_1965;
assign x_24455 = v_1968 | ~v_1966;
assign x_24456 = v_1968 | ~v_1967;
assign x_24457 = v_98 | v_103 | v_101 | v_100 | v_102 | v_170 | v_169 | v_150 | v_149 | v_148 | v_147 | v_184 | ~v_609 | ~v_608 | ~v_299 | ~v_298 | ~v_435 | ~v_434 | ~v_607 | ~v_606 | ~v_1898 | ~v_1897 | ~v_1896 | ~v_1895 | ~v_1894 | ~v_1893 | ~v_1930 | ~v_1929 | ~v_1928 | ~v_1927 | ~v_281 | ~v_280 | ~v_279 | ~v_278 | ~v_277 | ~v_276 | ~v_427 | ~v_426 | ~v_425 | ~v_424 | ~v_1888 | ~v_1887 | ~v_1886 | ~v_1885 | v_1967;
assign x_24458 = v_56 | v_61 | v_60 | v_59 | v_58 | v_144 | v_145 | v_143 | v_142 | v_166 | v_165 | v_183 | ~v_604 | ~v_603 | ~v_266 | ~v_265 | ~v_420 | ~v_419 | ~v_602 | ~v_601 | ~v_1883 | ~v_1882 | ~v_1881 | ~v_1880 | ~v_1879 | ~v_1878 | ~v_1925 | ~v_1924 | ~v_1923 | ~v_1922 | ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_244 | ~v_243 | ~v_412 | ~v_411 | ~v_410 | ~v_409 | ~v_1873 | ~v_1872 | ~v_1871 | ~v_1870 | v_1966;
assign x_24459 = v_13 | v_18 | v_17 | v_16 | v_15 | v_136 | v_135 | v_134 | v_137 | v_162 | v_161 | v_182 | ~v_599 | ~v_598 | ~v_233 | ~v_232 | ~v_405 | ~v_404 | ~v_597 | ~v_596 | ~v_1868 | ~v_1867 | ~v_1866 | ~v_1865 | ~v_1864 | ~v_1863 | ~v_1920 | ~v_1919 | ~v_1918 | ~v_1917 | ~v_215 | ~v_214 | ~v_213 | ~v_212 | ~v_211 | ~v_210 | ~v_397 | ~v_396 | ~v_395 | ~v_394 | ~v_1858 | ~v_1857 | ~v_1856 | ~v_1855 | v_1965;
assign x_24460 = v_1964 | ~v_1953;
assign x_24461 = v_1964 | ~v_1958;
assign x_24462 = v_1964 | ~v_1963;
assign x_24463 = v_103 | v_101 | v_94 | v_99 | v_102 | v_171 | v_169 | v_149 | v_148 | v_147 | v_184 | v_181 | ~v_483 | ~v_482 | ~v_481 | ~v_480 | ~v_345 | ~v_479 | ~v_478 | ~v_344 | ~v_1962 | ~v_1961 | ~v_1896 | ~v_1960 | ~v_1959 | ~v_1893 | ~v_1914 | ~v_1913 | ~v_1912 | ~v_1911 | ~v_473 | ~v_472 | ~v_279 | ~v_471 | ~v_470 | ~v_276 | ~v_335 | ~v_334 | ~v_333 | ~v_332 | ~v_1888 | ~v_1887 | ~v_1886 | ~v_1885 | v_1963;
assign x_24464 = v_1962 | v_139;
assign x_24465 = v_1962 | v_130;
assign x_24466 = v_1961 | v_140;
assign x_24467 = v_1961 | v_122;
assign x_24468 = v_1960 | ~v_139;
assign x_24469 = v_1960 | v_115;
assign x_24470 = v_1959 | ~v_140;
assign x_24471 = v_1959 | v_107;
assign x_24472 = v_61 | v_52 | v_60 | v_59 | v_57 | v_144 | v_180 | v_143 | v_142 | v_167 | v_165 | v_183 | ~v_468 | ~v_467 | ~v_466 | ~v_465 | ~v_330 | ~v_464 | ~v_463 | ~v_329 | ~v_1957 | ~v_1956 | ~v_1881 | ~v_1955 | ~v_1954 | ~v_1878 | ~v_1909 | ~v_1908 | ~v_1907 | ~v_1906 | ~v_458 | ~v_457 | ~v_246 | ~v_456 | ~v_455 | ~v_243 | ~v_320 | ~v_319 | ~v_318 | ~v_317 | ~v_1873 | ~v_1872 | ~v_1871 | ~v_1870 | v_1958;
assign x_24473 = v_1957 | v_139;
assign x_24474 = v_1957 | v_88;
assign x_24475 = v_1956 | v_140;
assign x_24476 = v_1956 | v_80;
assign x_24477 = v_1955 | ~v_139;
assign x_24478 = v_1955 | v_73;
assign x_24479 = v_1954 | ~v_140;
assign x_24480 = v_1954 | v_65;
assign x_24481 = v_9 | v_18 | v_17 | v_16 | v_14 | ~v_453 | ~v_452 | v_136 | v_135 | v_134 | v_179 | v_163 | v_161 | v_182 | ~v_451 | ~v_450 | ~v_315 | ~v_449 | ~v_448 | ~v_314 | ~v_1952 | ~v_1951 | ~v_1866 | ~v_1950 | ~v_1949 | ~v_1863 | ~v_1904 | ~v_1903 | ~v_1902 | ~v_1901 | ~v_443 | ~v_442 | ~v_213 | ~v_441 | ~v_440 | ~v_210 | ~v_305 | ~v_304 | ~v_303 | ~v_302 | ~v_1858 | ~v_1857 | ~v_1856 | ~v_1855 | v_1953;
assign x_24482 = v_1952 | v_139;
assign x_24483 = v_1952 | v_46;
assign x_24484 = v_1951 | v_140;
assign x_24485 = v_1951 | v_38;
assign x_24486 = v_1950 | ~v_139;
assign x_24487 = v_1950 | v_31;
assign x_24488 = v_1949 | ~v_140;
assign x_24489 = v_1949 | v_23;
assign x_24490 = v_1948 | ~v_1937;
assign x_24491 = v_1948 | ~v_1942;
assign x_24492 = v_1948 | ~v_1947;
assign x_24493 = v_103 | v_101 | v_96 | v_94 | v_102 | v_171 | v_169 | v_150 | v_149 | v_147 | v_184 | v_181 | ~v_391 | ~v_390 | ~v_389 | ~v_388 | ~v_387 | ~v_386 | ~v_345 | ~v_344 | ~v_385 | ~v_384 | ~v_1896 | ~v_1893 | ~v_1946 | ~v_1945 | ~v_1944 | ~v_1943 | ~v_1914 | ~v_1913 | ~v_1912 | ~v_1911 | ~v_279 | ~v_276 | ~v_335 | ~v_334 | ~v_333 | ~v_332 | ~v_379 | ~v_378 | ~v_1888 | ~v_1887 | ~v_1886 | ~v_1885 | v_1947;
assign x_24494 = v_1946 | v_141;
assign x_24495 = v_1946 | v_130;
assign x_24496 = v_1945 | v_141;
assign x_24497 = v_1945 | v_122;
assign x_24498 = v_1944 | ~v_141;
assign x_24499 = v_1944 | v_115;
assign x_24500 = v_1943 | ~v_141;
assign x_24501 = v_1943 | v_107;
assign x_24502 = v_54 | v_61 | v_52 | v_60 | v_59 | v_144 | v_180 | v_145 | v_142 | v_167 | v_165 | v_183 | ~v_376 | ~v_375 | ~v_374 | ~v_373 | ~v_372 | ~v_371 | ~v_330 | ~v_329 | ~v_370 | ~v_369 | ~v_1881 | ~v_1878 | ~v_1941 | ~v_1940 | ~v_1939 | ~v_1938 | ~v_1909 | ~v_1908 | ~v_1907 | ~v_1906 | ~v_246 | ~v_243 | ~v_320 | ~v_319 | ~v_318 | ~v_317 | ~v_364 | ~v_363 | ~v_1873 | ~v_1872 | ~v_1871 | ~v_1870 | v_1942;
assign x_24503 = v_1941 | v_141;
assign x_24504 = v_1941 | v_88;
assign x_24505 = v_1940 | v_141;
assign x_24506 = v_1940 | v_80;
assign x_24507 = v_1939 | ~v_141;
assign x_24508 = v_1939 | v_73;
assign x_24509 = v_1938 | ~v_141;
assign x_24510 = v_1938 | v_65;
assign x_24511 = v_9 | v_18 | v_17 | v_16 | v_11 | v_136 | v_134 | v_137 | v_179 | v_163 | v_161 | v_182 | ~v_361 | ~v_360 | ~v_359 | ~v_358 | ~v_357 | ~v_356 | ~v_315 | ~v_314 | ~v_355 | ~v_354 | ~v_1866 | ~v_1863 | ~v_1936 | ~v_1935 | ~v_1934 | ~v_1933 | ~v_1904 | ~v_1903 | ~v_1902 | ~v_1901 | ~v_213 | ~v_210 | ~v_305 | ~v_304 | ~v_303 | ~v_302 | ~v_349 | ~v_348 | ~v_1858 | ~v_1857 | ~v_1856 | ~v_1855 | v_1937;
assign x_24512 = v_1936 | v_141;
assign x_24513 = v_1936 | v_46;
assign x_24514 = v_1935 | v_141;
assign x_24515 = v_1935 | v_38;
assign x_24516 = v_1934 | ~v_141;
assign x_24517 = v_1934 | v_31;
assign x_24518 = v_1933 | ~v_141;
assign x_24519 = v_1933 | v_23;
assign x_24520 = v_1932 | ~v_1921;
assign x_24521 = v_1932 | ~v_1926;
assign x_24522 = v_1932 | ~v_1931;
assign x_24523 = v_101 | v_94 | v_102 | v_172 | v_171 | v_169 | v_150 | v_149 | v_148 | v_147 | v_184 | v_181 | ~v_437 | ~v_436 | ~v_435 | ~v_434 | ~v_345 | ~v_344 | ~v_433 | ~v_432 | ~v_1896 | ~v_1893 | ~v_1930 | ~v_1929 | ~v_1928 | ~v_1927 | ~v_1914 | ~v_1913 | ~v_1912 | ~v_1911 | ~v_279 | ~v_276 | ~v_335 | ~v_334 | ~v_333 | ~v_332 | ~v_427 | ~v_426 | ~v_425 | ~v_424 | ~v_1888 | ~v_1887 | ~v_1886 | ~v_1885 | v_1931;
assign x_24524 = v_1930 | v_174;
assign x_24525 = v_1930 | v_130;
assign x_24526 = v_1929 | v_173;
assign x_24527 = v_1929 | v_122;
assign x_24528 = v_1928 | ~v_174;
assign x_24529 = v_1928 | v_115;
assign x_24530 = v_1927 | ~v_173;
assign x_24531 = v_1927 | v_107;
assign x_24532 = v_52 | v_60 | v_59 | v_144 | v_180 | v_145 | v_143 | v_142 | v_168 | v_167 | v_165 | v_183 | ~v_422 | ~v_421 | ~v_420 | ~v_419 | ~v_330 | ~v_329 | ~v_418 | ~v_417 | ~v_1881 | ~v_1878 | ~v_1925 | ~v_1924 | ~v_1923 | ~v_1922 | ~v_1909 | ~v_1908 | ~v_1907 | ~v_1906 | ~v_246 | ~v_243 | ~v_320 | ~v_319 | ~v_318 | ~v_317 | ~v_412 | ~v_411 | ~v_410 | ~v_409 | ~v_1873 | ~v_1872 | ~v_1871 | ~v_1870 | v_1926;
assign x_24533 = v_1925 | v_174;
assign x_24534 = v_1925 | v_88;
assign x_24535 = v_1924 | v_173;
assign x_24536 = v_1924 | v_80;
assign x_24537 = v_1923 | ~v_174;
assign x_24538 = v_1923 | v_73;
assign x_24539 = v_1922 | ~v_173;
assign x_24540 = v_1922 | v_65;
assign x_24541 = v_9 | v_17 | v_16 | v_136 | v_135 | v_134 | v_137 | v_179 | v_164 | v_163 | v_161 | v_182 | ~v_407 | ~v_406 | ~v_405 | ~v_404 | ~v_315 | ~v_314 | ~v_403 | ~v_402 | ~v_1866 | ~v_1863 | ~v_1920 | ~v_1919 | ~v_1918 | ~v_1917 | ~v_1904 | ~v_1903 | ~v_1902 | ~v_1901 | ~v_213 | ~v_210 | ~v_305 | ~v_304 | ~v_303 | ~v_302 | ~v_397 | ~v_396 | ~v_395 | ~v_394 | ~v_1858 | ~v_1857 | ~v_1856 | ~v_1855 | v_1921;
assign x_24542 = v_1920 | v_174;
assign x_24543 = v_1920 | v_46;
assign x_24544 = v_1919 | v_173;
assign x_24545 = v_1919 | v_38;
assign x_24546 = v_1918 | ~v_174;
assign x_24547 = v_1918 | v_31;
assign x_24548 = v_1917 | ~v_173;
assign x_24549 = v_1917 | v_23;
assign x_24550 = v_1916 | ~v_1905;
assign x_24551 = v_1916 | ~v_1910;
assign x_24552 = v_1916 | ~v_1915;
assign x_24553 = v_103 | v_97 | v_95 | v_94 | v_102 | v_171 | v_169 | v_160 | v_150 | v_148 | v_184 | v_181 | ~v_297 | ~v_296 | ~v_345 | ~v_344 | ~v_343 | ~v_342 | ~v_341 | ~v_340 | ~v_1896 | ~v_1893 | ~v_1892 | ~v_1891 | ~v_1890 | ~v_1889 | ~v_1914 | ~v_1913 | ~v_1912 | ~v_1911 | ~v_279 | ~v_276 | ~v_335 | ~v_334 | ~v_333 | ~v_332 | ~v_275 | ~v_274 | ~v_273 | ~v_272 | ~v_1888 | ~v_1887 | ~v_1886 | ~v_1885 | v_1915;
assign x_24554 = v_1914 | v_176;
assign x_24555 = v_1914 | v_127;
assign x_24556 = v_1913 | v_175;
assign x_24557 = v_1913 | v_121;
assign x_24558 = v_1912 | ~v_176;
assign x_24559 = v_1912 | v_112;
assign x_24560 = v_1911 | ~v_175;
assign x_24561 = v_1911 | v_106;
assign x_24562 = v_53 | v_55 | v_61 | v_52 | v_60 | v_180 | v_159 | v_145 | v_143 | v_167 | v_165 | v_183 | ~v_264 | ~v_263 | ~v_330 | ~v_329 | ~v_328 | ~v_327 | ~v_326 | ~v_325 | ~v_1881 | ~v_1878 | ~v_1877 | ~v_1876 | ~v_1875 | ~v_1874 | ~v_1909 | ~v_1908 | ~v_1907 | ~v_1906 | ~v_246 | ~v_243 | ~v_320 | ~v_319 | ~v_318 | ~v_317 | ~v_242 | ~v_241 | ~v_240 | ~v_239 | ~v_1873 | ~v_1872 | ~v_1871 | ~v_1870 | v_1910;
assign x_24563 = v_1909 | v_176;
assign x_24564 = v_1909 | v_85;
assign x_24565 = v_1908 | v_175;
assign x_24566 = v_1908 | v_79;
assign x_24567 = v_1907 | ~v_176;
assign x_24568 = v_1907 | v_70;
assign x_24569 = v_1906 | ~v_175;
assign x_24570 = v_1906 | v_64;
assign x_24571 = v_9 | v_18 | v_17 | v_12 | v_10 | v_135 | v_137 | v_179 | v_163 | v_161 | v_155 | v_182 | ~v_231 | ~v_230 | ~v_315 | ~v_314 | ~v_313 | ~v_312 | ~v_311 | ~v_310 | ~v_1866 | ~v_1863 | ~v_1862 | ~v_1861 | ~v_1860 | ~v_1859 | ~v_1904 | ~v_1903 | ~v_1902 | ~v_1901 | ~v_213 | ~v_210 | ~v_305 | ~v_304 | ~v_303 | ~v_302 | ~v_209 | ~v_208 | ~v_207 | ~v_206 | ~v_1858 | ~v_1857 | ~v_1856 | ~v_1855 | v_1905;
assign x_24572 = v_1904 | v_176;
assign x_24573 = v_1904 | v_43;
assign x_24574 = v_1903 | v_175;
assign x_24575 = v_1903 | v_37;
assign x_24576 = v_1902 | ~v_176;
assign x_24577 = v_1902 | v_28;
assign x_24578 = v_1901 | ~v_175;
assign x_24579 = v_1901 | v_22;
assign x_24580 = v_1900 | ~v_1869;
assign x_24581 = v_1900 | ~v_1884;
assign x_24582 = v_1900 | ~v_1899;
assign x_24583 = v_98 | v_103 | v_97 | v_100 | v_102 | v_170 | v_169 | v_160 | v_150 | v_148 | v_147 | v_184 | ~v_299 | ~v_298 | ~v_297 | ~v_296 | ~v_295 | ~v_294 | ~v_293 | ~v_292 | ~v_1898 | ~v_1897 | ~v_1896 | ~v_1895 | ~v_1894 | ~v_1893 | ~v_1892 | ~v_1891 | ~v_1890 | ~v_1889 | ~v_281 | ~v_280 | ~v_279 | ~v_278 | ~v_277 | ~v_276 | ~v_275 | ~v_274 | ~v_273 | ~v_272 | ~v_1888 | ~v_1887 | ~v_1886 | ~v_1885 | v_1899;
assign x_24584 = v_1898 | v_139;
assign x_24585 = v_1898 | v_127;
assign x_24586 = v_1897 | v_140;
assign x_24587 = v_1897 | v_121;
assign x_24588 = v_1896 | v_141;
assign x_24589 = v_1896 | v_119;
assign x_24590 = v_1895 | ~v_139;
assign x_24591 = v_1895 | v_112;
assign x_24592 = v_1894 | ~v_140;
assign x_24593 = v_1894 | v_106;
assign x_24594 = v_1893 | ~v_141;
assign x_24595 = v_1893 | v_104;
assign x_24596 = v_1892 | v_176;
assign x_24597 = v_1892 | v_130;
assign x_24598 = v_1891 | v_175;
assign x_24599 = v_1891 | v_122;
assign x_24600 = v_1890 | ~v_176;
assign x_24601 = v_1890 | v_115;
assign x_24602 = v_1889 | ~v_175;
assign x_24603 = v_1889 | v_107;
assign x_24604 = v_1888 | v_176;
assign x_24605 = v_1888 | v_123;
assign x_24606 = v_1887 | v_175;
assign x_24607 = v_1887 | v_120;
assign x_24608 = v_1886 | ~v_176;
assign x_24609 = v_1886 | v_108;
assign x_24610 = v_1885 | ~v_175;
assign x_24611 = v_1885 | v_105;
assign x_24612 = v_56 | v_55 | v_61 | v_60 | v_58 | v_159 | v_145 | v_143 | v_142 | v_166 | v_165 | v_183 | ~v_266 | ~v_265 | ~v_264 | ~v_263 | ~v_262 | ~v_261 | ~v_260 | ~v_259 | ~v_1883 | ~v_1882 | ~v_1881 | ~v_1880 | ~v_1879 | ~v_1878 | ~v_1877 | ~v_1876 | ~v_1875 | ~v_1874 | ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_244 | ~v_243 | ~v_242 | ~v_241 | ~v_240 | ~v_239 | ~v_1873 | ~v_1872 | ~v_1871 | ~v_1870 | v_1884;
assign x_24613 = v_1883 | v_139;
assign x_24614 = v_1883 | v_85;
assign x_24615 = v_1882 | v_140;
assign x_24616 = v_1882 | v_79;
assign x_24617 = v_1881 | v_141;
assign x_24618 = v_1881 | v_77;
assign x_24619 = v_1880 | ~v_139;
assign x_24620 = v_1880 | v_70;
assign x_24621 = v_1879 | ~v_140;
assign x_24622 = v_1879 | v_64;
assign x_24623 = v_1878 | ~v_141;
assign x_24624 = v_1878 | v_62;
assign x_24625 = v_1877 | v_176;
assign x_24626 = v_1877 | v_88;
assign x_24627 = v_1876 | v_175;
assign x_24628 = v_1876 | v_80;
assign x_24629 = v_1875 | ~v_176;
assign x_24630 = v_1875 | v_73;
assign x_24631 = v_1874 | ~v_175;
assign x_24632 = v_1874 | v_65;
assign x_24633 = v_1873 | v_176;
assign x_24634 = v_1873 | v_81;
assign x_24635 = v_1872 | v_175;
assign x_24636 = v_1872 | v_78;
assign x_24637 = v_1871 | ~v_176;
assign x_24638 = v_1871 | v_66;
assign x_24639 = v_1870 | ~v_175;
assign x_24640 = v_1870 | v_63;
assign x_24641 = v_13 | v_18 | v_17 | v_15 | v_12 | v_135 | v_134 | v_137 | v_162 | v_161 | v_155 | v_182 | ~v_233 | ~v_232 | ~v_231 | ~v_230 | ~v_229 | ~v_228 | ~v_227 | ~v_226 | ~v_1868 | ~v_1867 | ~v_1866 | ~v_1865 | ~v_1864 | ~v_1863 | ~v_1862 | ~v_1861 | ~v_1860 | ~v_1859 | ~v_215 | ~v_214 | ~v_213 | ~v_212 | ~v_211 | ~v_210 | ~v_209 | ~v_208 | ~v_207 | ~v_206 | ~v_1858 | ~v_1857 | ~v_1856 | ~v_1855 | v_1869;
assign x_24642 = v_1868 | v_139;
assign x_24643 = v_1868 | v_43;
assign x_24644 = v_1867 | v_140;
assign x_24645 = v_1867 | v_37;
assign x_24646 = v_1866 | v_141;
assign x_24647 = v_1866 | v_35;
assign x_24648 = v_1865 | ~v_139;
assign x_24649 = v_1865 | v_28;
assign x_24650 = v_1864 | ~v_140;
assign x_24651 = v_1864 | v_22;
assign x_24652 = v_1863 | ~v_141;
assign x_24653 = v_1863 | v_20;
assign x_24654 = v_1862 | v_176;
assign x_24655 = v_1862 | v_46;
assign x_24656 = v_1861 | v_175;
assign x_24657 = v_1861 | v_38;
assign x_24658 = v_1860 | ~v_176;
assign x_24659 = v_1860 | v_31;
assign x_24660 = v_1859 | ~v_175;
assign x_24661 = v_1859 | v_23;
assign x_24662 = v_1858 | v_176;
assign x_24663 = v_1858 | v_39;
assign x_24664 = v_1857 | v_175;
assign x_24665 = v_1857 | v_36;
assign x_24666 = v_1856 | ~v_176;
assign x_24667 = v_1856 | v_24;
assign x_24668 = v_1855 | ~v_175;
assign x_24669 = v_1855 | v_21;
assign x_24670 = v_1854 | ~v_1852;
assign x_24671 = v_1854 | ~v_1853;
assign x_24672 = v_1854 | ~v_187;
assign x_24673 = v_1854 | ~v_190;
assign x_24674 = v_1854 | ~v_176;
assign x_24675 = v_1854 | ~v_175;
assign x_24676 = ~v_186 | ~v_197 | v_1853;
assign x_24677 = ~v_189 | ~v_1851 | v_1852;
assign x_24678 = v_1851 | ~v_199;
assign x_24679 = v_1851 | ~v_200;
assign x_24680 = v_1851 | ~v_178;
assign x_24681 = v_1851 | ~v_177;
assign x_24682 = v_1850 | ~v_1559;
assign x_24683 = v_1850 | ~v_1849;
assign x_24684 = v_177 | v_178 | ~v_1848 | ~v_742 | ~v_741 | ~v_1567 | ~v_1563 | v_1849;
assign x_24685 = v_1848 | ~v_1643;
assign x_24686 = v_1848 | ~v_1671;
assign x_24687 = v_1848 | ~v_1699;
assign x_24688 = v_1848 | ~v_1727;
assign x_24689 = v_1848 | ~v_1755;
assign x_24690 = v_1848 | ~v_1759;
assign x_24691 = v_1848 | ~v_1787;
assign x_24692 = v_1848 | ~v_1791;
assign x_24693 = v_1848 | ~v_1795;
assign x_24694 = v_1848 | ~v_1799;
assign x_24695 = v_1848 | ~v_1803;
assign x_24696 = v_1848 | ~v_1831;
assign x_24697 = v_1848 | ~v_1835;
assign x_24698 = v_1848 | ~v_1839;
assign x_24699 = v_1848 | ~v_1843;
assign x_24700 = v_1848 | ~v_1847;
assign x_24701 = v_1848 | ~v_1263;
assign x_24702 = v_1848 | ~v_1264;
assign x_24703 = v_1848 | ~v_1265;
assign x_24704 = v_1848 | ~v_1266;
assign x_24705 = ~v_1846 | ~v_1845 | ~v_1844 | v_1847;
assign x_24706 = v_1846 | ~v_1618;
assign x_24707 = v_1846 | ~v_1619;
assign x_24708 = v_1846 | ~v_1620;
assign x_24709 = v_1846 | ~v_1621;
assign x_24710 = v_1846 | ~v_1626;
assign x_24711 = v_1846 | ~v_1627;
assign x_24712 = v_1846 | ~v_1746;
assign x_24713 = v_1846 | ~v_1628;
assign x_24714 = v_1846 | ~v_1747;
assign x_24715 = v_1846 | ~v_1629;
assign x_24716 = v_1846 | ~v_1630;
assign x_24717 = v_1846 | ~v_1748;
assign x_24718 = v_1846 | ~v_1631;
assign x_24719 = v_1846 | ~v_1749;
assign x_24720 = v_1846 | ~v_1636;
assign x_24721 = v_1846 | ~v_1637;
assign x_24722 = v_1846 | ~v_1750;
assign x_24723 = v_1846 | ~v_1638;
assign x_24724 = v_1846 | ~v_1751;
assign x_24725 = v_1846 | ~v_1639;
assign x_24726 = v_1846 | ~v_1640;
assign x_24727 = v_1846 | ~v_1752;
assign x_24728 = v_1846 | ~v_1641;
assign x_24729 = v_1846 | ~v_1753;
assign x_24730 = v_1846 | ~v_839;
assign x_24731 = v_1846 | ~v_1257;
assign x_24732 = v_1846 | ~v_1023;
assign x_24733 = v_1846 | ~v_840;
assign x_24734 = v_1846 | ~v_1258;
assign x_24735 = v_1846 | ~v_1024;
assign x_24736 = v_1846 | ~v_184;
assign x_24737 = v_1846 | ~v_170;
assign x_24738 = v_1846 | ~v_169;
assign x_24739 = v_1846 | ~v_149;
assign x_24740 = v_1846 | ~v_148;
assign x_24741 = v_1846 | ~v_1259;
assign x_24742 = v_1846 | ~v_1260;
assign x_24743 = v_1846 | ~v_103;
assign x_24744 = v_1846 | ~v_102;
assign x_24745 = v_1846 | ~v_101;
assign x_24746 = v_1846 | ~v_100;
assign x_24747 = v_1846 | ~v_99;
assign x_24748 = v_1846 | ~v_98;
assign x_24749 = v_1846 | ~v_95;
assign x_24750 = v_1845 | ~v_1593;
assign x_24751 = v_1845 | ~v_1594;
assign x_24752 = v_1845 | ~v_1595;
assign x_24753 = v_1845 | ~v_1596;
assign x_24754 = v_1845 | ~v_1601;
assign x_24755 = v_1845 | ~v_1602;
assign x_24756 = v_1845 | ~v_1737;
assign x_24757 = v_1845 | ~v_1603;
assign x_24758 = v_1845 | ~v_1738;
assign x_24759 = v_1845 | ~v_1604;
assign x_24760 = v_1845 | ~v_1605;
assign x_24761 = v_1845 | ~v_1739;
assign x_24762 = v_1845 | ~v_1606;
assign x_24763 = v_1845 | ~v_1740;
assign x_24764 = v_1845 | ~v_1611;
assign x_24765 = v_1845 | ~v_1612;
assign x_24766 = v_1845 | ~v_1741;
assign x_24767 = v_1845 | ~v_1613;
assign x_24768 = v_1845 | ~v_1742;
assign x_24769 = v_1845 | ~v_1614;
assign x_24770 = v_1845 | ~v_1615;
assign x_24771 = v_1845 | ~v_1743;
assign x_24772 = v_1845 | ~v_1616;
assign x_24773 = v_1845 | ~v_1744;
assign x_24774 = v_1845 | ~v_806;
assign x_24775 = v_1845 | ~v_1252;
assign x_24776 = v_1845 | ~v_1008;
assign x_24777 = v_1845 | ~v_1253;
assign x_24778 = v_1845 | ~v_1009;
assign x_24779 = v_1845 | ~v_807;
assign x_24780 = v_1845 | ~v_183;
assign x_24781 = v_1845 | ~v_166;
assign x_24782 = v_1845 | ~v_165;
assign x_24783 = v_1845 | ~v_144;
assign x_24784 = v_1845 | ~v_143;
assign x_24785 = v_1845 | ~v_1254;
assign x_24786 = v_1845 | ~v_1255;
assign x_24787 = v_1845 | ~v_61;
assign x_24788 = v_1845 | ~v_60;
assign x_24789 = v_1845 | ~v_59;
assign x_24790 = v_1845 | ~v_58;
assign x_24791 = v_1845 | ~v_57;
assign x_24792 = v_1845 | ~v_56;
assign x_24793 = v_1845 | ~v_53;
assign x_24794 = v_1844 | ~v_1568;
assign x_24795 = v_1844 | ~v_1569;
assign x_24796 = v_1844 | ~v_1570;
assign x_24797 = v_1844 | ~v_1571;
assign x_24798 = v_1844 | ~v_1576;
assign x_24799 = v_1844 | ~v_1577;
assign x_24800 = v_1844 | ~v_1728;
assign x_24801 = v_1844 | ~v_1578;
assign x_24802 = v_1844 | ~v_1729;
assign x_24803 = v_1844 | ~v_1579;
assign x_24804 = v_1844 | ~v_1580;
assign x_24805 = v_1844 | ~v_1730;
assign x_24806 = v_1844 | ~v_1581;
assign x_24807 = v_1844 | ~v_1731;
assign x_24808 = v_1844 | ~v_1586;
assign x_24809 = v_1844 | ~v_1587;
assign x_24810 = v_1844 | ~v_1732;
assign x_24811 = v_1844 | ~v_1588;
assign x_24812 = v_1844 | ~v_1733;
assign x_24813 = v_1844 | ~v_1589;
assign x_24814 = v_1844 | ~v_1590;
assign x_24815 = v_1844 | ~v_1734;
assign x_24816 = v_1844 | ~v_1591;
assign x_24817 = v_1844 | ~v_1735;
assign x_24818 = v_1844 | ~v_773;
assign x_24819 = v_1844 | ~v_774;
assign x_24820 = v_1844 | ~v_182;
assign x_24821 = v_1844 | ~v_162;
assign x_24822 = v_1844 | ~v_161;
assign x_24823 = v_1844 | ~v_1247;
assign x_24824 = v_1844 | ~v_1248;
assign x_24825 = v_1844 | ~v_136;
assign x_24826 = v_1844 | ~v_135;
assign x_24827 = v_1844 | ~v_1249;
assign x_24828 = v_1844 | ~v_993;
assign x_24829 = v_1844 | ~v_1250;
assign x_24830 = v_1844 | ~v_994;
assign x_24831 = v_1844 | ~v_18;
assign x_24832 = v_1844 | ~v_17;
assign x_24833 = v_1844 | ~v_16;
assign x_24834 = v_1844 | ~v_15;
assign x_24835 = v_1844 | ~v_14;
assign x_24836 = v_1844 | ~v_13;
assign x_24837 = v_1844 | ~v_10;
assign x_24838 = ~v_1842 | ~v_1841 | ~v_1840 | v_1843;
assign x_24839 = v_1842 | ~v_1618;
assign x_24840 = v_1842 | ~v_1619;
assign x_24841 = v_1842 | ~v_1620;
assign x_24842 = v_1842 | ~v_1621;
assign x_24843 = v_1842 | ~v_1822;
assign x_24844 = v_1842 | ~v_1823;
assign x_24845 = v_1842 | ~v_1824;
assign x_24846 = v_1842 | ~v_1825;
assign x_24847 = v_1842 | ~v_1626;
assign x_24848 = v_1842 | ~v_1746;
assign x_24849 = v_1842 | ~v_1747;
assign x_24850 = v_1842 | ~v_1629;
assign x_24851 = v_1842 | ~v_1748;
assign x_24852 = v_1842 | ~v_1749;
assign x_24853 = v_1842 | ~v_1826;
assign x_24854 = v_1842 | ~v_1827;
assign x_24855 = v_1842 | ~v_1828;
assign x_24856 = v_1842 | ~v_1829;
assign x_24857 = v_1842 | ~v_1636;
assign x_24858 = v_1842 | ~v_1750;
assign x_24859 = v_1842 | ~v_1751;
assign x_24860 = v_1842 | ~v_1639;
assign x_24861 = v_1842 | ~v_1752;
assign x_24862 = v_1842 | ~v_1753;
assign x_24863 = v_1842 | ~v_885;
assign x_24864 = v_1842 | ~v_1019;
assign x_24865 = v_1842 | ~v_1020;
assign x_24866 = v_1842 | ~v_886;
assign x_24867 = v_1842 | ~v_1021;
assign x_24868 = v_1842 | ~v_1022;
assign x_24869 = v_1842 | ~v_1023;
assign x_24870 = v_1842 | ~v_1024;
assign x_24871 = v_1842 | ~v_184;
assign x_24872 = v_1842 | ~v_181;
assign x_24873 = v_1842 | ~v_171;
assign x_24874 = v_1842 | ~v_170;
assign x_24875 = v_1842 | ~v_149;
assign x_24876 = v_1842 | ~v_148;
assign x_24877 = v_1842 | ~v_147;
assign x_24878 = v_1842 | ~v_103;
assign x_24879 = v_1842 | ~v_102;
assign x_24880 = v_1842 | ~v_101;
assign x_24881 = v_1842 | ~v_99;
assign x_24882 = v_1842 | ~v_93;
assign x_24883 = v_1841 | ~v_1593;
assign x_24884 = v_1841 | ~v_1594;
assign x_24885 = v_1841 | ~v_1595;
assign x_24886 = v_1841 | ~v_1596;
assign x_24887 = v_1841 | ~v_1813;
assign x_24888 = v_1841 | ~v_1814;
assign x_24889 = v_1841 | ~v_1815;
assign x_24890 = v_1841 | ~v_1816;
assign x_24891 = v_1841 | ~v_1601;
assign x_24892 = v_1841 | ~v_1737;
assign x_24893 = v_1841 | ~v_1738;
assign x_24894 = v_1841 | ~v_1604;
assign x_24895 = v_1841 | ~v_1739;
assign x_24896 = v_1841 | ~v_1740;
assign x_24897 = v_1841 | ~v_1817;
assign x_24898 = v_1841 | ~v_1818;
assign x_24899 = v_1841 | ~v_1819;
assign x_24900 = v_1841 | ~v_1820;
assign x_24901 = v_1841 | ~v_1611;
assign x_24902 = v_1841 | ~v_1741;
assign x_24903 = v_1841 | ~v_1742;
assign x_24904 = v_1841 | ~v_1614;
assign x_24905 = v_1841 | ~v_1743;
assign x_24906 = v_1841 | ~v_1744;
assign x_24907 = v_1841 | ~v_870;
assign x_24908 = v_1841 | ~v_1004;
assign x_24909 = v_1841 | ~v_1005;
assign x_24910 = v_1841 | ~v_871;
assign x_24911 = v_1841 | ~v_1006;
assign x_24912 = v_1841 | ~v_1007;
assign x_24913 = v_1841 | ~v_1008;
assign x_24914 = v_1841 | ~v_1009;
assign x_24915 = v_1841 | ~v_183;
assign x_24916 = v_1841 | ~v_180;
assign x_24917 = v_1841 | ~v_167;
assign x_24918 = v_1841 | ~v_166;
assign x_24919 = v_1841 | ~v_144;
assign x_24920 = v_1841 | ~v_143;
assign x_24921 = v_1841 | ~v_142;
assign x_24922 = v_1841 | ~v_61;
assign x_24923 = v_1841 | ~v_60;
assign x_24924 = v_1841 | ~v_59;
assign x_24925 = v_1841 | ~v_57;
assign x_24926 = v_1841 | ~v_51;
assign x_24927 = v_1840 | ~v_1568;
assign x_24928 = v_1840 | ~v_1569;
assign x_24929 = v_1840 | ~v_1570;
assign x_24930 = v_1840 | ~v_1571;
assign x_24931 = v_1840 | ~v_1804;
assign x_24932 = v_1840 | ~v_1805;
assign x_24933 = v_1840 | ~v_1806;
assign x_24934 = v_1840 | ~v_1807;
assign x_24935 = v_1840 | ~v_1576;
assign x_24936 = v_1840 | ~v_1728;
assign x_24937 = v_1840 | ~v_1729;
assign x_24938 = v_1840 | ~v_1579;
assign x_24939 = v_1840 | ~v_1730;
assign x_24940 = v_1840 | ~v_1731;
assign x_24941 = v_1840 | ~v_1808;
assign x_24942 = v_1840 | ~v_1809;
assign x_24943 = v_1840 | ~v_1810;
assign x_24944 = v_1840 | ~v_1811;
assign x_24945 = v_1840 | ~v_1586;
assign x_24946 = v_1840 | ~v_1732;
assign x_24947 = v_1840 | ~v_1733;
assign x_24948 = v_1840 | ~v_1589;
assign x_24949 = v_1840 | ~v_1734;
assign x_24950 = v_1840 | ~v_1735;
assign x_24951 = v_1840 | ~v_855;
assign x_24952 = v_1840 | ~v_989;
assign x_24953 = v_1840 | ~v_990;
assign x_24954 = v_1840 | ~v_856;
assign x_24955 = v_1840 | ~v_991;
assign x_24956 = v_1840 | ~v_992;
assign x_24957 = v_1840 | ~v_182;
assign x_24958 = v_1840 | ~v_179;
assign x_24959 = v_1840 | ~v_163;
assign x_24960 = v_1840 | ~v_162;
assign x_24961 = v_1840 | ~v_136;
assign x_24962 = v_1840 | ~v_135;
assign x_24963 = v_1840 | ~v_134;
assign x_24964 = v_1840 | ~v_993;
assign x_24965 = v_1840 | ~v_994;
assign x_24966 = v_1840 | ~v_18;
assign x_24967 = v_1840 | ~v_17;
assign x_24968 = v_1840 | ~v_16;
assign x_24969 = v_1840 | ~v_14;
assign x_24970 = v_1840 | ~v_8;
assign x_24971 = ~v_1838 | ~v_1837 | ~v_1836 | v_1839;
assign x_24972 = v_1838 | ~v_1618;
assign x_24973 = v_1838 | ~v_1619;
assign x_24974 = v_1838 | ~v_1620;
assign x_24975 = v_1838 | ~v_1621;
assign x_24976 = v_1838 | ~v_1718;
assign x_24977 = v_1838 | ~v_1719;
assign x_24978 = v_1838 | ~v_1720;
assign x_24979 = v_1838 | ~v_1721;
assign x_24980 = v_1838 | ~v_1822;
assign x_24981 = v_1838 | ~v_1823;
assign x_24982 = v_1838 | ~v_1824;
assign x_24983 = v_1838 | ~v_1825;
assign x_24984 = v_1838 | ~v_1626;
assign x_24985 = v_1838 | ~v_1629;
assign x_24986 = v_1838 | ~v_1826;
assign x_24987 = v_1838 | ~v_1827;
assign x_24988 = v_1838 | ~v_1828;
assign x_24989 = v_1838 | ~v_1829;
assign x_24990 = v_1838 | ~v_1722;
assign x_24991 = v_1838 | ~v_1723;
assign x_24992 = v_1838 | ~v_1724;
assign x_24993 = v_1838 | ~v_1725;
assign x_24994 = v_1838 | ~v_1636;
assign x_24995 = v_1838 | ~v_1639;
assign x_24996 = v_1838 | ~v_881;
assign x_24997 = v_1838 | ~v_882;
assign x_24998 = v_1838 | ~v_883;
assign x_24999 = v_1838 | ~v_884;
assign x_25000 = v_1838 | ~v_885;
assign x_25001 = v_1838 | ~v_886;
assign x_25002 = v_1838 | ~v_837;
assign x_25003 = v_1838 | ~v_838;
assign x_25004 = v_1838 | ~v_184;
assign x_25005 = v_1838 | ~v_181;
assign x_25006 = v_1838 | ~v_171;
assign x_25007 = v_1838 | ~v_170;
assign x_25008 = v_1838 | ~v_160;
assign x_25009 = v_1838 | ~v_150;
assign x_25010 = v_1838 | ~v_149;
assign x_25011 = v_1838 | ~v_103;
assign x_25012 = v_1838 | ~v_102;
assign x_25013 = v_1838 | ~v_96;
assign x_25014 = v_1838 | ~v_95;
assign x_25015 = v_1838 | ~v_93;
assign x_25016 = v_1837 | ~v_1593;
assign x_25017 = v_1837 | ~v_1594;
assign x_25018 = v_1837 | ~v_1595;
assign x_25019 = v_1837 | ~v_1596;
assign x_25020 = v_1837 | ~v_1709;
assign x_25021 = v_1837 | ~v_1710;
assign x_25022 = v_1837 | ~v_1711;
assign x_25023 = v_1837 | ~v_1712;
assign x_25024 = v_1837 | ~v_1813;
assign x_25025 = v_1837 | ~v_1814;
assign x_25026 = v_1837 | ~v_1815;
assign x_25027 = v_1837 | ~v_1816;
assign x_25028 = v_1837 | ~v_1601;
assign x_25029 = v_1837 | ~v_1604;
assign x_25030 = v_1837 | ~v_1817;
assign x_25031 = v_1837 | ~v_1818;
assign x_25032 = v_1837 | ~v_1819;
assign x_25033 = v_1837 | ~v_1820;
assign x_25034 = v_1837 | ~v_1713;
assign x_25035 = v_1837 | ~v_1714;
assign x_25036 = v_1837 | ~v_1715;
assign x_25037 = v_1837 | ~v_1716;
assign x_25038 = v_1837 | ~v_1611;
assign x_25039 = v_1837 | ~v_1614;
assign x_25040 = v_1837 | ~v_866;
assign x_25041 = v_1837 | ~v_867;
assign x_25042 = v_1837 | ~v_868;
assign x_25043 = v_1837 | ~v_869;
assign x_25044 = v_1837 | ~v_870;
assign x_25045 = v_1837 | ~v_871;
assign x_25046 = v_1837 | ~v_804;
assign x_25047 = v_1837 | ~v_805;
assign x_25048 = v_1837 | ~v_183;
assign x_25049 = v_1837 | ~v_180;
assign x_25050 = v_1837 | ~v_167;
assign x_25051 = v_1837 | ~v_166;
assign x_25052 = v_1837 | ~v_159;
assign x_25053 = v_1837 | ~v_145;
assign x_25054 = v_1837 | ~v_144;
assign x_25055 = v_1837 | ~v_61;
assign x_25056 = v_1837 | ~v_60;
assign x_25057 = v_1837 | ~v_54;
assign x_25058 = v_1837 | ~v_53;
assign x_25059 = v_1837 | ~v_51;
assign x_25060 = v_1836 | ~v_1568;
assign x_25061 = v_1836 | ~v_1569;
assign x_25062 = v_1836 | ~v_1570;
assign x_25063 = v_1836 | ~v_1571;
assign x_25064 = v_1836 | ~v_1700;
assign x_25065 = v_1836 | ~v_1701;
assign x_25066 = v_1836 | ~v_1702;
assign x_25067 = v_1836 | ~v_1703;
assign x_25068 = v_1836 | ~v_1804;
assign x_25069 = v_1836 | ~v_1805;
assign x_25070 = v_1836 | ~v_1806;
assign x_25071 = v_1836 | ~v_1807;
assign x_25072 = v_1836 | ~v_1576;
assign x_25073 = v_1836 | ~v_1579;
assign x_25074 = v_1836 | ~v_1808;
assign x_25075 = v_1836 | ~v_1809;
assign x_25076 = v_1836 | ~v_1810;
assign x_25077 = v_1836 | ~v_1811;
assign x_25078 = v_1836 | ~v_1704;
assign x_25079 = v_1836 | ~v_1705;
assign x_25080 = v_1836 | ~v_1706;
assign x_25081 = v_1836 | ~v_1707;
assign x_25082 = v_1836 | ~v_1586;
assign x_25083 = v_1836 | ~v_1589;
assign x_25084 = v_1836 | ~v_851;
assign x_25085 = v_1836 | ~v_852;
assign x_25086 = v_1836 | ~v_853;
assign x_25087 = v_1836 | ~v_854;
assign x_25088 = v_1836 | ~v_855;
assign x_25089 = v_1836 | ~v_856;
assign x_25090 = v_1836 | ~v_771;
assign x_25091 = v_1836 | ~v_772;
assign x_25092 = v_1836 | ~v_182;
assign x_25093 = v_1836 | ~v_179;
assign x_25094 = v_1836 | ~v_163;
assign x_25095 = v_1836 | ~v_162;
assign x_25096 = v_1836 | ~v_155;
assign x_25097 = v_1836 | ~v_137;
assign x_25098 = v_1836 | ~v_136;
assign x_25099 = v_1836 | ~v_18;
assign x_25100 = v_1836 | ~v_17;
assign x_25101 = v_1836 | ~v_11;
assign x_25102 = v_1836 | ~v_10;
assign x_25103 = v_1836 | ~v_8;
assign x_25104 = ~v_1834 | ~v_1833 | ~v_1832 | v_1835;
assign x_25105 = v_1834 | ~v_1618;
assign x_25106 = v_1834 | ~v_1619;
assign x_25107 = v_1834 | ~v_1620;
assign x_25108 = v_1834 | ~v_1621;
assign x_25109 = v_1834 | ~v_1690;
assign x_25110 = v_1834 | ~v_1691;
assign x_25111 = v_1834 | ~v_1692;
assign x_25112 = v_1834 | ~v_1693;
assign x_25113 = v_1834 | ~v_1822;
assign x_25114 = v_1834 | ~v_1823;
assign x_25115 = v_1834 | ~v_1824;
assign x_25116 = v_1834 | ~v_1825;
assign x_25117 = v_1834 | ~v_1626;
assign x_25118 = v_1834 | ~v_1629;
assign x_25119 = v_1834 | ~v_1826;
assign x_25120 = v_1834 | ~v_1827;
assign x_25121 = v_1834 | ~v_1828;
assign x_25122 = v_1834 | ~v_1829;
assign x_25123 = v_1834 | ~v_1694;
assign x_25124 = v_1834 | ~v_1695;
assign x_25125 = v_1834 | ~v_1696;
assign x_25126 = v_1834 | ~v_1697;
assign x_25127 = v_1834 | ~v_1636;
assign x_25128 = v_1834 | ~v_1639;
assign x_25129 = v_1834 | ~v_925;
assign x_25130 = v_1834 | ~v_926;
assign x_25131 = v_1834 | ~v_885;
assign x_25132 = v_1834 | ~v_886;
assign x_25133 = v_1834 | ~v_927;
assign x_25134 = v_1834 | ~v_928;
assign x_25135 = v_1834 | ~v_929;
assign x_25136 = v_1834 | ~v_930;
assign x_25137 = v_1834 | ~v_184;
assign x_25138 = v_1834 | ~v_181;
assign x_25139 = v_1834 | ~v_171;
assign x_25140 = v_1834 | ~v_170;
assign x_25141 = v_1834 | ~v_150;
assign x_25142 = v_1834 | ~v_149;
assign x_25143 = v_1834 | ~v_148;
assign x_25144 = v_1834 | ~v_147;
assign x_25145 = v_1834 | ~v_103;
assign x_25146 = v_1834 | ~v_102;
assign x_25147 = v_1834 | ~v_101;
assign x_25148 = v_1834 | ~v_93;
assign x_25149 = v_1833 | ~v_1593;
assign x_25150 = v_1833 | ~v_1594;
assign x_25151 = v_1833 | ~v_1595;
assign x_25152 = v_1833 | ~v_1596;
assign x_25153 = v_1833 | ~v_1681;
assign x_25154 = v_1833 | ~v_1682;
assign x_25155 = v_1833 | ~v_1683;
assign x_25156 = v_1833 | ~v_1684;
assign x_25157 = v_1833 | ~v_1813;
assign x_25158 = v_1833 | ~v_1814;
assign x_25159 = v_1833 | ~v_1815;
assign x_25160 = v_1833 | ~v_1816;
assign x_25161 = v_1833 | ~v_1601;
assign x_25162 = v_1833 | ~v_1604;
assign x_25163 = v_1833 | ~v_1817;
assign x_25164 = v_1833 | ~v_1818;
assign x_25165 = v_1833 | ~v_1819;
assign x_25166 = v_1833 | ~v_1820;
assign x_25167 = v_1833 | ~v_1685;
assign x_25168 = v_1833 | ~v_1686;
assign x_25169 = v_1833 | ~v_1687;
assign x_25170 = v_1833 | ~v_1688;
assign x_25171 = v_1833 | ~v_1611;
assign x_25172 = v_1833 | ~v_1614;
assign x_25173 = v_1833 | ~v_910;
assign x_25174 = v_1833 | ~v_911;
assign x_25175 = v_1833 | ~v_870;
assign x_25176 = v_1833 | ~v_871;
assign x_25177 = v_1833 | ~v_912;
assign x_25178 = v_1833 | ~v_913;
assign x_25179 = v_1833 | ~v_914;
assign x_25180 = v_1833 | ~v_915;
assign x_25181 = v_1833 | ~v_183;
assign x_25182 = v_1833 | ~v_180;
assign x_25183 = v_1833 | ~v_167;
assign x_25184 = v_1833 | ~v_166;
assign x_25185 = v_1833 | ~v_145;
assign x_25186 = v_1833 | ~v_144;
assign x_25187 = v_1833 | ~v_143;
assign x_25188 = v_1833 | ~v_142;
assign x_25189 = v_1833 | ~v_61;
assign x_25190 = v_1833 | ~v_60;
assign x_25191 = v_1833 | ~v_59;
assign x_25192 = v_1833 | ~v_51;
assign x_25193 = v_1832 | ~v_1568;
assign x_25194 = v_1832 | ~v_1569;
assign x_25195 = v_1832 | ~v_1570;
assign x_25196 = v_1832 | ~v_1571;
assign x_25197 = v_1832 | ~v_1672;
assign x_25198 = v_1832 | ~v_1673;
assign x_25199 = v_1832 | ~v_1674;
assign x_25200 = v_1832 | ~v_1675;
assign x_25201 = v_1832 | ~v_1804;
assign x_25202 = v_1832 | ~v_1805;
assign x_25203 = v_1832 | ~v_1806;
assign x_25204 = v_1832 | ~v_1807;
assign x_25205 = v_1832 | ~v_1576;
assign x_25206 = v_1832 | ~v_1579;
assign x_25207 = v_1832 | ~v_1808;
assign x_25208 = v_1832 | ~v_1809;
assign x_25209 = v_1832 | ~v_1810;
assign x_25210 = v_1832 | ~v_1811;
assign x_25211 = v_1832 | ~v_1676;
assign x_25212 = v_1832 | ~v_1677;
assign x_25213 = v_1832 | ~v_1678;
assign x_25214 = v_1832 | ~v_1679;
assign x_25215 = v_1832 | ~v_1586;
assign x_25216 = v_1832 | ~v_1589;
assign x_25217 = v_1832 | ~v_895;
assign x_25218 = v_1832 | ~v_896;
assign x_25219 = v_1832 | ~v_855;
assign x_25220 = v_1832 | ~v_856;
assign x_25221 = v_1832 | ~v_897;
assign x_25222 = v_1832 | ~v_898;
assign x_25223 = v_1832 | ~v_899;
assign x_25224 = v_1832 | ~v_900;
assign x_25225 = v_1832 | ~v_182;
assign x_25226 = v_1832 | ~v_179;
assign x_25227 = v_1832 | ~v_163;
assign x_25228 = v_1832 | ~v_162;
assign x_25229 = v_1832 | ~v_137;
assign x_25230 = v_1832 | ~v_136;
assign x_25231 = v_1832 | ~v_135;
assign x_25232 = v_1832 | ~v_134;
assign x_25233 = v_1832 | ~v_18;
assign x_25234 = v_1832 | ~v_17;
assign x_25235 = v_1832 | ~v_16;
assign x_25236 = v_1832 | ~v_8;
assign x_25237 = ~v_1830 | ~v_1821 | ~v_1812 | v_1831;
assign x_25238 = v_1830 | ~v_1618;
assign x_25239 = v_1830 | ~v_1619;
assign x_25240 = v_1830 | ~v_1620;
assign x_25241 = v_1830 | ~v_1621;
assign x_25242 = v_1830 | ~v_1622;
assign x_25243 = v_1830 | ~v_1623;
assign x_25244 = v_1830 | ~v_1624;
assign x_25245 = v_1830 | ~v_1625;
assign x_25246 = v_1830 | ~v_1822;
assign x_25247 = v_1830 | ~v_1823;
assign x_25248 = v_1830 | ~v_1824;
assign x_25249 = v_1830 | ~v_1825;
assign x_25250 = v_1830 | ~v_1626;
assign x_25251 = v_1830 | ~v_1629;
assign x_25252 = v_1830 | ~v_1826;
assign x_25253 = v_1830 | ~v_1827;
assign x_25254 = v_1830 | ~v_1828;
assign x_25255 = v_1830 | ~v_1829;
assign x_25256 = v_1830 | ~v_1632;
assign x_25257 = v_1830 | ~v_1633;
assign x_25258 = v_1830 | ~v_1634;
assign x_25259 = v_1830 | ~v_1635;
assign x_25260 = v_1830 | ~v_1636;
assign x_25261 = v_1830 | ~v_1639;
assign x_25262 = v_1830 | ~v_973;
assign x_25263 = v_1830 | ~v_974;
assign x_25264 = v_1830 | ~v_885;
assign x_25265 = v_1830 | ~v_886;
assign x_25266 = v_1830 | ~v_975;
assign x_25267 = v_1830 | ~v_976;
assign x_25268 = v_1830 | ~v_977;
assign x_25269 = v_1830 | ~v_978;
assign x_25270 = v_1830 | ~v_184;
assign x_25271 = v_1830 | ~v_181;
assign x_25272 = v_1830 | ~v_172;
assign x_25273 = v_1830 | ~v_171;
assign x_25274 = v_1830 | ~v_170;
assign x_25275 = v_1830 | ~v_150;
assign x_25276 = v_1830 | ~v_148;
assign x_25277 = v_1830 | ~v_147;
assign x_25278 = v_1830 | ~v_102;
assign x_25279 = v_1830 | ~v_101;
assign x_25280 = v_1830 | ~v_97;
assign x_25281 = v_1830 | ~v_93;
assign x_25282 = ~v_128 | ~v_178 | v_1829;
assign x_25283 = ~v_125 | ~v_177 | v_1828;
assign x_25284 = ~v_113 | v_178 | v_1827;
assign x_25285 = ~v_110 | v_177 | v_1826;
assign x_25286 = ~v_127 | ~v_158 | v_1825;
assign x_25287 = ~v_121 | ~v_158 | v_1824;
assign x_25288 = ~v_112 | v_158 | v_1823;
assign x_25289 = ~v_106 | v_158 | v_1822;
assign x_25290 = v_1821 | ~v_1593;
assign x_25291 = v_1821 | ~v_1594;
assign x_25292 = v_1821 | ~v_1595;
assign x_25293 = v_1821 | ~v_1596;
assign x_25294 = v_1821 | ~v_1597;
assign x_25295 = v_1821 | ~v_1598;
assign x_25296 = v_1821 | ~v_1599;
assign x_25297 = v_1821 | ~v_1600;
assign x_25298 = v_1821 | ~v_1813;
assign x_25299 = v_1821 | ~v_1814;
assign x_25300 = v_1821 | ~v_1815;
assign x_25301 = v_1821 | ~v_1816;
assign x_25302 = v_1821 | ~v_1601;
assign x_25303 = v_1821 | ~v_1604;
assign x_25304 = v_1821 | ~v_1817;
assign x_25305 = v_1821 | ~v_1818;
assign x_25306 = v_1821 | ~v_1819;
assign x_25307 = v_1821 | ~v_1820;
assign x_25308 = v_1821 | ~v_1607;
assign x_25309 = v_1821 | ~v_1608;
assign x_25310 = v_1821 | ~v_1609;
assign x_25311 = v_1821 | ~v_1610;
assign x_25312 = v_1821 | ~v_1611;
assign x_25313 = v_1821 | ~v_1614;
assign x_25314 = v_1821 | ~v_958;
assign x_25315 = v_1821 | ~v_959;
assign x_25316 = v_1821 | ~v_870;
assign x_25317 = v_1821 | ~v_871;
assign x_25318 = v_1821 | ~v_960;
assign x_25319 = v_1821 | ~v_961;
assign x_25320 = v_1821 | ~v_962;
assign x_25321 = v_1821 | ~v_963;
assign x_25322 = v_1821 | ~v_183;
assign x_25323 = v_1821 | ~v_180;
assign x_25324 = v_1821 | ~v_168;
assign x_25325 = v_1821 | ~v_167;
assign x_25326 = v_1821 | ~v_166;
assign x_25327 = v_1821 | ~v_145;
assign x_25328 = v_1821 | ~v_143;
assign x_25329 = v_1821 | ~v_142;
assign x_25330 = v_1821 | ~v_60;
assign x_25331 = v_1821 | ~v_59;
assign x_25332 = v_1821 | ~v_55;
assign x_25333 = v_1821 | ~v_51;
assign x_25334 = ~v_86 | ~v_178 | v_1820;
assign x_25335 = ~v_83 | ~v_177 | v_1819;
assign x_25336 = ~v_71 | v_178 | v_1818;
assign x_25337 = ~v_68 | v_177 | v_1817;
assign x_25338 = ~v_85 | ~v_158 | v_1816;
assign x_25339 = ~v_79 | ~v_158 | v_1815;
assign x_25340 = ~v_70 | v_158 | v_1814;
assign x_25341 = ~v_64 | v_158 | v_1813;
assign x_25342 = v_1812 | ~v_1568;
assign x_25343 = v_1812 | ~v_1569;
assign x_25344 = v_1812 | ~v_1570;
assign x_25345 = v_1812 | ~v_1571;
assign x_25346 = v_1812 | ~v_1572;
assign x_25347 = v_1812 | ~v_1573;
assign x_25348 = v_1812 | ~v_1574;
assign x_25349 = v_1812 | ~v_1575;
assign x_25350 = v_1812 | ~v_1804;
assign x_25351 = v_1812 | ~v_1805;
assign x_25352 = v_1812 | ~v_1806;
assign x_25353 = v_1812 | ~v_1807;
assign x_25354 = v_1812 | ~v_1576;
assign x_25355 = v_1812 | ~v_1579;
assign x_25356 = v_1812 | ~v_1808;
assign x_25357 = v_1812 | ~v_1809;
assign x_25358 = v_1812 | ~v_1810;
assign x_25359 = v_1812 | ~v_1811;
assign x_25360 = v_1812 | ~v_1582;
assign x_25361 = v_1812 | ~v_1583;
assign x_25362 = v_1812 | ~v_1584;
assign x_25363 = v_1812 | ~v_1585;
assign x_25364 = v_1812 | ~v_1586;
assign x_25365 = v_1812 | ~v_1589;
assign x_25366 = v_1812 | ~v_943;
assign x_25367 = v_1812 | ~v_944;
assign x_25368 = v_1812 | ~v_855;
assign x_25369 = v_1812 | ~v_856;
assign x_25370 = v_1812 | ~v_945;
assign x_25371 = v_1812 | ~v_946;
assign x_25372 = v_1812 | ~v_947;
assign x_25373 = v_1812 | ~v_948;
assign x_25374 = v_1812 | ~v_182;
assign x_25375 = v_1812 | ~v_179;
assign x_25376 = v_1812 | ~v_164;
assign x_25377 = v_1812 | ~v_163;
assign x_25378 = v_1812 | ~v_162;
assign x_25379 = v_1812 | ~v_137;
assign x_25380 = v_1812 | ~v_135;
assign x_25381 = v_1812 | ~v_134;
assign x_25382 = v_1812 | ~v_17;
assign x_25383 = v_1812 | ~v_16;
assign x_25384 = v_1812 | ~v_12;
assign x_25385 = v_1812 | ~v_8;
assign x_25386 = ~v_44 | ~v_178 | v_1811;
assign x_25387 = ~v_41 | ~v_177 | v_1810;
assign x_25388 = ~v_29 | v_178 | v_1809;
assign x_25389 = ~v_26 | v_177 | v_1808;
assign x_25390 = ~v_43 | ~v_158 | v_1807;
assign x_25391 = ~v_37 | ~v_158 | v_1806;
assign x_25392 = ~v_28 | v_158 | v_1805;
assign x_25393 = ~v_22 | v_158 | v_1804;
assign x_25394 = ~v_1802 | ~v_1801 | ~v_1800 | v_1803;
assign x_25395 = v_1802 | ~v_1618;
assign x_25396 = v_1802 | ~v_1619;
assign x_25397 = v_1802 | ~v_1620;
assign x_25398 = v_1802 | ~v_1621;
assign x_25399 = v_1802 | ~v_1718;
assign x_25400 = v_1802 | ~v_1719;
assign x_25401 = v_1802 | ~v_1720;
assign x_25402 = v_1802 | ~v_1721;
assign x_25403 = v_1802 | ~v_1626;
assign x_25404 = v_1802 | ~v_1627;
assign x_25405 = v_1802 | ~v_1628;
assign x_25406 = v_1802 | ~v_1629;
assign x_25407 = v_1802 | ~v_1630;
assign x_25408 = v_1802 | ~v_1631;
assign x_25409 = v_1802 | ~v_1722;
assign x_25410 = v_1802 | ~v_1723;
assign x_25411 = v_1802 | ~v_1724;
assign x_25412 = v_1802 | ~v_1725;
assign x_25413 = v_1802 | ~v_1636;
assign x_25414 = v_1802 | ~v_1637;
assign x_25415 = v_1802 | ~v_1638;
assign x_25416 = v_1802 | ~v_1639;
assign x_25417 = v_1802 | ~v_1640;
assign x_25418 = v_1802 | ~v_1641;
assign x_25419 = v_1802 | ~v_833;
assign x_25420 = v_1802 | ~v_834;
assign x_25421 = v_1802 | ~v_835;
assign x_25422 = v_1802 | ~v_836;
assign x_25423 = v_1802 | ~v_837;
assign x_25424 = v_1802 | ~v_838;
assign x_25425 = v_1802 | ~v_839;
assign x_25426 = v_1802 | ~v_840;
assign x_25427 = v_1802 | ~v_184;
assign x_25428 = v_1802 | ~v_170;
assign x_25429 = v_1802 | ~v_169;
assign x_25430 = v_1802 | ~v_160;
assign x_25431 = v_1802 | ~v_150;
assign x_25432 = v_1802 | ~v_149;
assign x_25433 = v_1802 | ~v_147;
assign x_25434 = v_1802 | ~v_103;
assign x_25435 = v_1802 | ~v_102;
assign x_25436 = v_1802 | ~v_100;
assign x_25437 = v_1802 | ~v_98;
assign x_25438 = v_1802 | ~v_96;
assign x_25439 = v_1801 | ~v_1593;
assign x_25440 = v_1801 | ~v_1594;
assign x_25441 = v_1801 | ~v_1595;
assign x_25442 = v_1801 | ~v_1596;
assign x_25443 = v_1801 | ~v_1709;
assign x_25444 = v_1801 | ~v_1710;
assign x_25445 = v_1801 | ~v_1711;
assign x_25446 = v_1801 | ~v_1712;
assign x_25447 = v_1801 | ~v_1601;
assign x_25448 = v_1801 | ~v_1602;
assign x_25449 = v_1801 | ~v_1603;
assign x_25450 = v_1801 | ~v_1604;
assign x_25451 = v_1801 | ~v_1605;
assign x_25452 = v_1801 | ~v_1606;
assign x_25453 = v_1801 | ~v_1713;
assign x_25454 = v_1801 | ~v_1714;
assign x_25455 = v_1801 | ~v_1715;
assign x_25456 = v_1801 | ~v_1716;
assign x_25457 = v_1801 | ~v_1611;
assign x_25458 = v_1801 | ~v_1612;
assign x_25459 = v_1801 | ~v_1613;
assign x_25460 = v_1801 | ~v_1614;
assign x_25461 = v_1801 | ~v_1615;
assign x_25462 = v_1801 | ~v_1616;
assign x_25463 = v_1801 | ~v_800;
assign x_25464 = v_1801 | ~v_801;
assign x_25465 = v_1801 | ~v_802;
assign x_25466 = v_1801 | ~v_803;
assign x_25467 = v_1801 | ~v_804;
assign x_25468 = v_1801 | ~v_805;
assign x_25469 = v_1801 | ~v_806;
assign x_25470 = v_1801 | ~v_807;
assign x_25471 = v_1801 | ~v_183;
assign x_25472 = v_1801 | ~v_166;
assign x_25473 = v_1801 | ~v_165;
assign x_25474 = v_1801 | ~v_159;
assign x_25475 = v_1801 | ~v_145;
assign x_25476 = v_1801 | ~v_144;
assign x_25477 = v_1801 | ~v_142;
assign x_25478 = v_1801 | ~v_61;
assign x_25479 = v_1801 | ~v_60;
assign x_25480 = v_1801 | ~v_58;
assign x_25481 = v_1801 | ~v_56;
assign x_25482 = v_1801 | ~v_54;
assign x_25483 = v_1800 | ~v_1568;
assign x_25484 = v_1800 | ~v_1569;
assign x_25485 = v_1800 | ~v_1570;
assign x_25486 = v_1800 | ~v_1571;
assign x_25487 = v_1800 | ~v_1700;
assign x_25488 = v_1800 | ~v_1701;
assign x_25489 = v_1800 | ~v_1702;
assign x_25490 = v_1800 | ~v_1703;
assign x_25491 = v_1800 | ~v_1576;
assign x_25492 = v_1800 | ~v_1577;
assign x_25493 = v_1800 | ~v_1578;
assign x_25494 = v_1800 | ~v_1579;
assign x_25495 = v_1800 | ~v_1580;
assign x_25496 = v_1800 | ~v_1581;
assign x_25497 = v_1800 | ~v_1704;
assign x_25498 = v_1800 | ~v_1705;
assign x_25499 = v_1800 | ~v_1706;
assign x_25500 = v_1800 | ~v_1707;
assign x_25501 = v_1800 | ~v_1586;
assign x_25502 = v_1800 | ~v_1587;
assign x_25503 = v_1800 | ~v_1588;
assign x_25504 = v_1800 | ~v_1589;
assign x_25505 = v_1800 | ~v_1590;
assign x_25506 = v_1800 | ~v_1591;
assign x_25507 = v_1800 | ~v_767;
assign x_25508 = v_1800 | ~v_768;
assign x_25509 = v_1800 | ~v_769;
assign x_25510 = v_1800 | ~v_770;
assign x_25511 = v_1800 | ~v_771;
assign x_25512 = v_1800 | ~v_772;
assign x_25513 = v_1800 | ~v_773;
assign x_25514 = v_1800 | ~v_774;
assign x_25515 = v_1800 | ~v_182;
assign x_25516 = v_1800 | ~v_162;
assign x_25517 = v_1800 | ~v_161;
assign x_25518 = v_1800 | ~v_155;
assign x_25519 = v_1800 | ~v_137;
assign x_25520 = v_1800 | ~v_136;
assign x_25521 = v_1800 | ~v_134;
assign x_25522 = v_1800 | ~v_18;
assign x_25523 = v_1800 | ~v_17;
assign x_25524 = v_1800 | ~v_15;
assign x_25525 = v_1800 | ~v_13;
assign x_25526 = v_1800 | ~v_11;
assign x_25527 = ~v_1798 | ~v_1797 | ~v_1796 | v_1799;
assign x_25528 = v_1798 | ~v_1618;
assign x_25529 = v_1798 | ~v_1619;
assign x_25530 = v_1798 | ~v_1620;
assign x_25531 = v_1798 | ~v_1621;
assign x_25532 = v_1798 | ~v_1778;
assign x_25533 = v_1798 | ~v_1779;
assign x_25534 = v_1798 | ~v_1780;
assign x_25535 = v_1798 | ~v_1781;
assign x_25536 = v_1798 | ~v_1626;
assign x_25537 = v_1798 | ~v_1746;
assign x_25538 = v_1798 | ~v_1747;
assign x_25539 = v_1798 | ~v_1629;
assign x_25540 = v_1798 | ~v_1748;
assign x_25541 = v_1798 | ~v_1749;
assign x_25542 = v_1798 | ~v_1782;
assign x_25543 = v_1798 | ~v_1783;
assign x_25544 = v_1798 | ~v_1784;
assign x_25545 = v_1798 | ~v_1785;
assign x_25546 = v_1798 | ~v_1636;
assign x_25547 = v_1798 | ~v_1750;
assign x_25548 = v_1798 | ~v_1751;
assign x_25549 = v_1798 | ~v_1639;
assign x_25550 = v_1798 | ~v_1752;
assign x_25551 = v_1798 | ~v_1753;
assign x_25552 = v_1798 | ~v_1085;
assign x_25553 = v_1798 | ~v_1131;
assign x_25554 = v_1798 | ~v_1132;
assign x_25555 = v_1798 | ~v_1086;
assign x_25556 = v_1798 | ~v_1133;
assign x_25557 = v_1798 | ~v_1134;
assign x_25558 = v_1798 | ~v_1023;
assign x_25559 = v_1798 | ~v_1024;
assign x_25560 = v_1798 | ~v_184;
assign x_25561 = v_1798 | ~v_172;
assign x_25562 = v_1798 | ~v_171;
assign x_25563 = v_1798 | ~v_170;
assign x_25564 = v_1798 | ~v_169;
assign x_25565 = v_1798 | ~v_149;
assign x_25566 = v_1798 | ~v_148;
assign x_25567 = v_1798 | ~v_147;
assign x_25568 = v_1798 | ~v_102;
assign x_25569 = v_1798 | ~v_101;
assign x_25570 = v_1798 | ~v_100;
assign x_25571 = v_1798 | ~v_99;
assign x_25572 = v_1797 | ~v_1593;
assign x_25573 = v_1797 | ~v_1594;
assign x_25574 = v_1797 | ~v_1595;
assign x_25575 = v_1797 | ~v_1596;
assign x_25576 = v_1797 | ~v_1769;
assign x_25577 = v_1797 | ~v_1770;
assign x_25578 = v_1797 | ~v_1771;
assign x_25579 = v_1797 | ~v_1772;
assign x_25580 = v_1797 | ~v_1601;
assign x_25581 = v_1797 | ~v_1737;
assign x_25582 = v_1797 | ~v_1738;
assign x_25583 = v_1797 | ~v_1604;
assign x_25584 = v_1797 | ~v_1739;
assign x_25585 = v_1797 | ~v_1740;
assign x_25586 = v_1797 | ~v_1773;
assign x_25587 = v_1797 | ~v_1774;
assign x_25588 = v_1797 | ~v_1775;
assign x_25589 = v_1797 | ~v_1776;
assign x_25590 = v_1797 | ~v_1611;
assign x_25591 = v_1797 | ~v_1741;
assign x_25592 = v_1797 | ~v_1742;
assign x_25593 = v_1797 | ~v_1614;
assign x_25594 = v_1797 | ~v_1743;
assign x_25595 = v_1797 | ~v_1744;
assign x_25596 = v_1797 | ~v_1070;
assign x_25597 = v_1797 | ~v_1126;
assign x_25598 = v_1797 | ~v_1127;
assign x_25599 = v_1797 | ~v_1071;
assign x_25600 = v_1797 | ~v_1128;
assign x_25601 = v_1797 | ~v_1129;
assign x_25602 = v_1797 | ~v_1008;
assign x_25603 = v_1797 | ~v_1009;
assign x_25604 = v_1797 | ~v_183;
assign x_25605 = v_1797 | ~v_168;
assign x_25606 = v_1797 | ~v_167;
assign x_25607 = v_1797 | ~v_166;
assign x_25608 = v_1797 | ~v_165;
assign x_25609 = v_1797 | ~v_144;
assign x_25610 = v_1797 | ~v_143;
assign x_25611 = v_1797 | ~v_142;
assign x_25612 = v_1797 | ~v_60;
assign x_25613 = v_1797 | ~v_59;
assign x_25614 = v_1797 | ~v_58;
assign x_25615 = v_1797 | ~v_57;
assign x_25616 = v_1796 | ~v_1568;
assign x_25617 = v_1796 | ~v_1569;
assign x_25618 = v_1796 | ~v_1570;
assign x_25619 = v_1796 | ~v_1571;
assign x_25620 = v_1796 | ~v_1760;
assign x_25621 = v_1796 | ~v_1761;
assign x_25622 = v_1796 | ~v_1762;
assign x_25623 = v_1796 | ~v_1763;
assign x_25624 = v_1796 | ~v_1576;
assign x_25625 = v_1796 | ~v_1728;
assign x_25626 = v_1796 | ~v_1729;
assign x_25627 = v_1796 | ~v_1579;
assign x_25628 = v_1796 | ~v_1730;
assign x_25629 = v_1796 | ~v_1731;
assign x_25630 = v_1796 | ~v_1764;
assign x_25631 = v_1796 | ~v_1765;
assign x_25632 = v_1796 | ~v_1766;
assign x_25633 = v_1796 | ~v_1767;
assign x_25634 = v_1796 | ~v_1586;
assign x_25635 = v_1796 | ~v_1732;
assign x_25636 = v_1796 | ~v_1733;
assign x_25637 = v_1796 | ~v_1589;
assign x_25638 = v_1796 | ~v_1734;
assign x_25639 = v_1796 | ~v_1735;
assign x_25640 = v_1796 | ~v_1055;
assign x_25641 = v_1796 | ~v_1121;
assign x_25642 = v_1796 | ~v_1122;
assign x_25643 = v_1796 | ~v_1056;
assign x_25644 = v_1796 | ~v_1123;
assign x_25645 = v_1796 | ~v_1124;
assign x_25646 = v_1796 | ~v_182;
assign x_25647 = v_1796 | ~v_164;
assign x_25648 = v_1796 | ~v_163;
assign x_25649 = v_1796 | ~v_162;
assign x_25650 = v_1796 | ~v_161;
assign x_25651 = v_1796 | ~v_136;
assign x_25652 = v_1796 | ~v_135;
assign x_25653 = v_1796 | ~v_134;
assign x_25654 = v_1796 | ~v_993;
assign x_25655 = v_1796 | ~v_994;
assign x_25656 = v_1796 | ~v_17;
assign x_25657 = v_1796 | ~v_16;
assign x_25658 = v_1796 | ~v_15;
assign x_25659 = v_1796 | ~v_14;
assign x_25660 = ~v_1794 | ~v_1793 | ~v_1792 | v_1795;
assign x_25661 = v_1794 | ~v_1618;
assign x_25662 = v_1794 | ~v_1619;
assign x_25663 = v_1794 | ~v_1620;
assign x_25664 = v_1794 | ~v_1621;
assign x_25665 = v_1794 | ~v_1778;
assign x_25666 = v_1794 | ~v_1779;
assign x_25667 = v_1794 | ~v_1780;
assign x_25668 = v_1794 | ~v_1781;
assign x_25669 = v_1794 | ~v_1718;
assign x_25670 = v_1794 | ~v_1719;
assign x_25671 = v_1794 | ~v_1720;
assign x_25672 = v_1794 | ~v_1721;
assign x_25673 = v_1794 | ~v_1626;
assign x_25674 = v_1794 | ~v_1629;
assign x_25675 = v_1794 | ~v_1782;
assign x_25676 = v_1794 | ~v_1783;
assign x_25677 = v_1794 | ~v_1784;
assign x_25678 = v_1794 | ~v_1785;
assign x_25679 = v_1794 | ~v_1722;
assign x_25680 = v_1794 | ~v_1723;
assign x_25681 = v_1794 | ~v_1724;
assign x_25682 = v_1794 | ~v_1725;
assign x_25683 = v_1794 | ~v_1636;
assign x_25684 = v_1794 | ~v_1639;
assign x_25685 = v_1794 | ~v_837;
assign x_25686 = v_1794 | ~v_838;
assign x_25687 = v_1794 | ~v_1081;
assign x_25688 = v_1794 | ~v_1082;
assign x_25689 = v_1794 | ~v_1083;
assign x_25690 = v_1794 | ~v_1084;
assign x_25691 = v_1794 | ~v_1085;
assign x_25692 = v_1794 | ~v_1086;
assign x_25693 = v_1794 | ~v_184;
assign x_25694 = v_1794 | ~v_171;
assign x_25695 = v_1794 | ~v_170;
assign x_25696 = v_1794 | ~v_169;
assign x_25697 = v_1794 | ~v_160;
assign x_25698 = v_1794 | ~v_150;
assign x_25699 = v_1794 | ~v_149;
assign x_25700 = v_1794 | ~v_147;
assign x_25701 = v_1794 | ~v_103;
assign x_25702 = v_1794 | ~v_102;
assign x_25703 = v_1794 | ~v_100;
assign x_25704 = v_1794 | ~v_96;
assign x_25705 = v_1793 | ~v_1593;
assign x_25706 = v_1793 | ~v_1594;
assign x_25707 = v_1793 | ~v_1595;
assign x_25708 = v_1793 | ~v_1596;
assign x_25709 = v_1793 | ~v_1769;
assign x_25710 = v_1793 | ~v_1770;
assign x_25711 = v_1793 | ~v_1771;
assign x_25712 = v_1793 | ~v_1772;
assign x_25713 = v_1793 | ~v_1709;
assign x_25714 = v_1793 | ~v_1710;
assign x_25715 = v_1793 | ~v_1711;
assign x_25716 = v_1793 | ~v_1712;
assign x_25717 = v_1793 | ~v_1601;
assign x_25718 = v_1793 | ~v_1604;
assign x_25719 = v_1793 | ~v_1773;
assign x_25720 = v_1793 | ~v_1774;
assign x_25721 = v_1793 | ~v_1775;
assign x_25722 = v_1793 | ~v_1776;
assign x_25723 = v_1793 | ~v_1713;
assign x_25724 = v_1793 | ~v_1714;
assign x_25725 = v_1793 | ~v_1715;
assign x_25726 = v_1793 | ~v_1716;
assign x_25727 = v_1793 | ~v_1611;
assign x_25728 = v_1793 | ~v_1614;
assign x_25729 = v_1793 | ~v_804;
assign x_25730 = v_1793 | ~v_805;
assign x_25731 = v_1793 | ~v_1066;
assign x_25732 = v_1793 | ~v_1067;
assign x_25733 = v_1793 | ~v_1068;
assign x_25734 = v_1793 | ~v_1069;
assign x_25735 = v_1793 | ~v_1070;
assign x_25736 = v_1793 | ~v_1071;
assign x_25737 = v_1793 | ~v_183;
assign x_25738 = v_1793 | ~v_167;
assign x_25739 = v_1793 | ~v_166;
assign x_25740 = v_1793 | ~v_165;
assign x_25741 = v_1793 | ~v_159;
assign x_25742 = v_1793 | ~v_145;
assign x_25743 = v_1793 | ~v_144;
assign x_25744 = v_1793 | ~v_142;
assign x_25745 = v_1793 | ~v_61;
assign x_25746 = v_1793 | ~v_60;
assign x_25747 = v_1793 | ~v_58;
assign x_25748 = v_1793 | ~v_54;
assign x_25749 = v_1792 | ~v_1568;
assign x_25750 = v_1792 | ~v_1569;
assign x_25751 = v_1792 | ~v_1570;
assign x_25752 = v_1792 | ~v_1571;
assign x_25753 = v_1792 | ~v_1760;
assign x_25754 = v_1792 | ~v_1761;
assign x_25755 = v_1792 | ~v_1762;
assign x_25756 = v_1792 | ~v_1763;
assign x_25757 = v_1792 | ~v_1700;
assign x_25758 = v_1792 | ~v_1701;
assign x_25759 = v_1792 | ~v_1702;
assign x_25760 = v_1792 | ~v_1703;
assign x_25761 = v_1792 | ~v_1576;
assign x_25762 = v_1792 | ~v_1579;
assign x_25763 = v_1792 | ~v_1764;
assign x_25764 = v_1792 | ~v_1765;
assign x_25765 = v_1792 | ~v_1766;
assign x_25766 = v_1792 | ~v_1767;
assign x_25767 = v_1792 | ~v_1704;
assign x_25768 = v_1792 | ~v_1705;
assign x_25769 = v_1792 | ~v_1706;
assign x_25770 = v_1792 | ~v_1707;
assign x_25771 = v_1792 | ~v_1586;
assign x_25772 = v_1792 | ~v_1589;
assign x_25773 = v_1792 | ~v_771;
assign x_25774 = v_1792 | ~v_772;
assign x_25775 = v_1792 | ~v_1051;
assign x_25776 = v_1792 | ~v_1052;
assign x_25777 = v_1792 | ~v_1053;
assign x_25778 = v_1792 | ~v_1054;
assign x_25779 = v_1792 | ~v_1055;
assign x_25780 = v_1792 | ~v_1056;
assign x_25781 = v_1792 | ~v_182;
assign x_25782 = v_1792 | ~v_163;
assign x_25783 = v_1792 | ~v_162;
assign x_25784 = v_1792 | ~v_161;
assign x_25785 = v_1792 | ~v_155;
assign x_25786 = v_1792 | ~v_137;
assign x_25787 = v_1792 | ~v_136;
assign x_25788 = v_1792 | ~v_134;
assign x_25789 = v_1792 | ~v_18;
assign x_25790 = v_1792 | ~v_17;
assign x_25791 = v_1792 | ~v_15;
assign x_25792 = v_1792 | ~v_11;
assign x_25793 = ~v_1790 | ~v_1789 | ~v_1788 | v_1791;
assign x_25794 = v_1790 | ~v_1618;
assign x_25795 = v_1790 | ~v_1619;
assign x_25796 = v_1790 | ~v_1620;
assign x_25797 = v_1790 | ~v_1621;
assign x_25798 = v_1790 | ~v_1778;
assign x_25799 = v_1790 | ~v_1779;
assign x_25800 = v_1790 | ~v_1780;
assign x_25801 = v_1790 | ~v_1781;
assign x_25802 = v_1790 | ~v_1690;
assign x_25803 = v_1790 | ~v_1691;
assign x_25804 = v_1790 | ~v_1692;
assign x_25805 = v_1790 | ~v_1693;
assign x_25806 = v_1790 | ~v_1626;
assign x_25807 = v_1790 | ~v_1629;
assign x_25808 = v_1790 | ~v_1782;
assign x_25809 = v_1790 | ~v_1783;
assign x_25810 = v_1790 | ~v_1784;
assign x_25811 = v_1790 | ~v_1785;
assign x_25812 = v_1790 | ~v_1694;
assign x_25813 = v_1790 | ~v_1695;
assign x_25814 = v_1790 | ~v_1696;
assign x_25815 = v_1790 | ~v_1697;
assign x_25816 = v_1790 | ~v_1636;
assign x_25817 = v_1790 | ~v_1639;
assign x_25818 = v_1790 | ~v_927;
assign x_25819 = v_1790 | ~v_928;
assign x_25820 = v_1790 | ~v_1099;
assign x_25821 = v_1790 | ~v_1100;
assign x_25822 = v_1790 | ~v_1101;
assign x_25823 = v_1790 | ~v_1102;
assign x_25824 = v_1790 | ~v_1085;
assign x_25825 = v_1790 | ~v_1086;
assign x_25826 = v_1790 | ~v_184;
assign x_25827 = v_1790 | ~v_171;
assign x_25828 = v_1790 | ~v_170;
assign x_25829 = v_1790 | ~v_169;
assign x_25830 = v_1790 | ~v_150;
assign x_25831 = v_1790 | ~v_149;
assign x_25832 = v_1790 | ~v_148;
assign x_25833 = v_1790 | ~v_103;
assign x_25834 = v_1790 | ~v_102;
assign x_25835 = v_1790 | ~v_101;
assign x_25836 = v_1790 | ~v_100;
assign x_25837 = v_1790 | ~v_95;
assign x_25838 = v_1789 | ~v_1593;
assign x_25839 = v_1789 | ~v_1594;
assign x_25840 = v_1789 | ~v_1595;
assign x_25841 = v_1789 | ~v_1596;
assign x_25842 = v_1789 | ~v_1769;
assign x_25843 = v_1789 | ~v_1770;
assign x_25844 = v_1789 | ~v_1771;
assign x_25845 = v_1789 | ~v_1772;
assign x_25846 = v_1789 | ~v_1681;
assign x_25847 = v_1789 | ~v_1682;
assign x_25848 = v_1789 | ~v_1683;
assign x_25849 = v_1789 | ~v_1684;
assign x_25850 = v_1789 | ~v_1601;
assign x_25851 = v_1789 | ~v_1604;
assign x_25852 = v_1789 | ~v_1773;
assign x_25853 = v_1789 | ~v_1774;
assign x_25854 = v_1789 | ~v_1775;
assign x_25855 = v_1789 | ~v_1776;
assign x_25856 = v_1789 | ~v_1685;
assign x_25857 = v_1789 | ~v_1686;
assign x_25858 = v_1789 | ~v_1687;
assign x_25859 = v_1789 | ~v_1688;
assign x_25860 = v_1789 | ~v_1611;
assign x_25861 = v_1789 | ~v_1614;
assign x_25862 = v_1789 | ~v_912;
assign x_25863 = v_1789 | ~v_913;
assign x_25864 = v_1789 | ~v_1094;
assign x_25865 = v_1789 | ~v_1095;
assign x_25866 = v_1789 | ~v_1096;
assign x_25867 = v_1789 | ~v_1097;
assign x_25868 = v_1789 | ~v_1070;
assign x_25869 = v_1789 | ~v_1071;
assign x_25870 = v_1789 | ~v_183;
assign x_25871 = v_1789 | ~v_167;
assign x_25872 = v_1789 | ~v_166;
assign x_25873 = v_1789 | ~v_165;
assign x_25874 = v_1789 | ~v_145;
assign x_25875 = v_1789 | ~v_144;
assign x_25876 = v_1789 | ~v_143;
assign x_25877 = v_1789 | ~v_61;
assign x_25878 = v_1789 | ~v_60;
assign x_25879 = v_1789 | ~v_59;
assign x_25880 = v_1789 | ~v_58;
assign x_25881 = v_1789 | ~v_53;
assign x_25882 = v_1788 | ~v_1568;
assign x_25883 = v_1788 | ~v_1569;
assign x_25884 = v_1788 | ~v_1570;
assign x_25885 = v_1788 | ~v_1571;
assign x_25886 = v_1788 | ~v_1760;
assign x_25887 = v_1788 | ~v_1761;
assign x_25888 = v_1788 | ~v_1762;
assign x_25889 = v_1788 | ~v_1763;
assign x_25890 = v_1788 | ~v_1672;
assign x_25891 = v_1788 | ~v_1673;
assign x_25892 = v_1788 | ~v_1674;
assign x_25893 = v_1788 | ~v_1675;
assign x_25894 = v_1788 | ~v_1576;
assign x_25895 = v_1788 | ~v_1579;
assign x_25896 = v_1788 | ~v_1764;
assign x_25897 = v_1788 | ~v_1765;
assign x_25898 = v_1788 | ~v_1766;
assign x_25899 = v_1788 | ~v_1767;
assign x_25900 = v_1788 | ~v_1676;
assign x_25901 = v_1788 | ~v_1677;
assign x_25902 = v_1788 | ~v_1678;
assign x_25903 = v_1788 | ~v_1679;
assign x_25904 = v_1788 | ~v_1586;
assign x_25905 = v_1788 | ~v_1589;
assign x_25906 = v_1788 | ~v_897;
assign x_25907 = v_1788 | ~v_898;
assign x_25908 = v_1788 | ~v_1089;
assign x_25909 = v_1788 | ~v_1090;
assign x_25910 = v_1788 | ~v_1091;
assign x_25911 = v_1788 | ~v_1092;
assign x_25912 = v_1788 | ~v_1055;
assign x_25913 = v_1788 | ~v_1056;
assign x_25914 = v_1788 | ~v_182;
assign x_25915 = v_1788 | ~v_163;
assign x_25916 = v_1788 | ~v_162;
assign x_25917 = v_1788 | ~v_161;
assign x_25918 = v_1788 | ~v_137;
assign x_25919 = v_1788 | ~v_136;
assign x_25920 = v_1788 | ~v_135;
assign x_25921 = v_1788 | ~v_18;
assign x_25922 = v_1788 | ~v_17;
assign x_25923 = v_1788 | ~v_16;
assign x_25924 = v_1788 | ~v_15;
assign x_25925 = v_1788 | ~v_10;
assign x_25926 = ~v_1786 | ~v_1777 | ~v_1768 | v_1787;
assign x_25927 = v_1786 | ~v_1618;
assign x_25928 = v_1786 | ~v_1619;
assign x_25929 = v_1786 | ~v_1620;
assign x_25930 = v_1786 | ~v_1621;
assign x_25931 = v_1786 | ~v_1778;
assign x_25932 = v_1786 | ~v_1779;
assign x_25933 = v_1786 | ~v_1780;
assign x_25934 = v_1786 | ~v_1781;
assign x_25935 = v_1786 | ~v_1622;
assign x_25936 = v_1786 | ~v_1623;
assign x_25937 = v_1786 | ~v_1624;
assign x_25938 = v_1786 | ~v_1625;
assign x_25939 = v_1786 | ~v_1626;
assign x_25940 = v_1786 | ~v_1629;
assign x_25941 = v_1786 | ~v_1782;
assign x_25942 = v_1786 | ~v_1783;
assign x_25943 = v_1786 | ~v_1784;
assign x_25944 = v_1786 | ~v_1785;
assign x_25945 = v_1786 | ~v_1632;
assign x_25946 = v_1786 | ~v_1633;
assign x_25947 = v_1786 | ~v_1634;
assign x_25948 = v_1786 | ~v_1635;
assign x_25949 = v_1786 | ~v_1636;
assign x_25950 = v_1786 | ~v_1639;
assign x_25951 = v_1786 | ~v_975;
assign x_25952 = v_1786 | ~v_976;
assign x_25953 = v_1786 | ~v_1115;
assign x_25954 = v_1786 | ~v_1116;
assign x_25955 = v_1786 | ~v_1085;
assign x_25956 = v_1786 | ~v_1086;
assign x_25957 = v_1786 | ~v_1117;
assign x_25958 = v_1786 | ~v_1118;
assign x_25959 = v_1786 | ~v_184;
assign x_25960 = v_1786 | ~v_171;
assign x_25961 = v_1786 | ~v_170;
assign x_25962 = v_1786 | ~v_169;
assign x_25963 = v_1786 | ~v_151;
assign x_25964 = v_1786 | ~v_150;
assign x_25965 = v_1786 | ~v_148;
assign x_25966 = v_1786 | ~v_147;
assign x_25967 = v_1786 | ~v_103;
assign x_25968 = v_1786 | ~v_101;
assign x_25969 = v_1786 | ~v_100;
assign x_25970 = v_1786 | ~v_97;
assign x_25971 = ~v_128 | ~v_173 | v_1785;
assign x_25972 = ~v_125 | ~v_174 | v_1784;
assign x_25973 = ~v_113 | v_173 | v_1783;
assign x_25974 = ~v_110 | v_174 | v_1782;
assign x_25975 = ~v_127 | ~v_175 | v_1781;
assign x_25976 = ~v_121 | ~v_176 | v_1780;
assign x_25977 = ~v_112 | v_175 | v_1779;
assign x_25978 = ~v_106 | v_176 | v_1778;
assign x_25979 = v_1777 | ~v_1593;
assign x_25980 = v_1777 | ~v_1594;
assign x_25981 = v_1777 | ~v_1595;
assign x_25982 = v_1777 | ~v_1596;
assign x_25983 = v_1777 | ~v_1769;
assign x_25984 = v_1777 | ~v_1770;
assign x_25985 = v_1777 | ~v_1771;
assign x_25986 = v_1777 | ~v_1772;
assign x_25987 = v_1777 | ~v_1597;
assign x_25988 = v_1777 | ~v_1598;
assign x_25989 = v_1777 | ~v_1599;
assign x_25990 = v_1777 | ~v_1600;
assign x_25991 = v_1777 | ~v_1601;
assign x_25992 = v_1777 | ~v_1604;
assign x_25993 = v_1777 | ~v_1773;
assign x_25994 = v_1777 | ~v_1774;
assign x_25995 = v_1777 | ~v_1775;
assign x_25996 = v_1777 | ~v_1776;
assign x_25997 = v_1777 | ~v_1607;
assign x_25998 = v_1777 | ~v_1608;
assign x_25999 = v_1777 | ~v_1609;
assign x_26000 = v_1777 | ~v_1610;
assign x_26001 = v_1777 | ~v_1611;
assign x_26002 = v_1777 | ~v_1614;
assign x_26003 = v_1777 | ~v_960;
assign x_26004 = v_1777 | ~v_961;
assign x_26005 = v_1777 | ~v_1110;
assign x_26006 = v_1777 | ~v_1111;
assign x_26007 = v_1777 | ~v_1070;
assign x_26008 = v_1777 | ~v_1071;
assign x_26009 = v_1777 | ~v_1112;
assign x_26010 = v_1777 | ~v_1113;
assign x_26011 = v_1777 | ~v_183;
assign x_26012 = v_1777 | ~v_167;
assign x_26013 = v_1777 | ~v_166;
assign x_26014 = v_1777 | ~v_165;
assign x_26015 = v_1777 | ~v_146;
assign x_26016 = v_1777 | ~v_145;
assign x_26017 = v_1777 | ~v_143;
assign x_26018 = v_1777 | ~v_142;
assign x_26019 = v_1777 | ~v_61;
assign x_26020 = v_1777 | ~v_59;
assign x_26021 = v_1777 | ~v_58;
assign x_26022 = v_1777 | ~v_55;
assign x_26023 = ~v_86 | ~v_173 | v_1776;
assign x_26024 = ~v_83 | ~v_174 | v_1775;
assign x_26025 = ~v_71 | v_173 | v_1774;
assign x_26026 = ~v_68 | v_174 | v_1773;
assign x_26027 = ~v_85 | ~v_175 | v_1772;
assign x_26028 = ~v_79 | ~v_176 | v_1771;
assign x_26029 = ~v_70 | v_175 | v_1770;
assign x_26030 = ~v_64 | v_176 | v_1769;
assign x_26031 = v_1768 | ~v_1568;
assign x_26032 = v_1768 | ~v_1569;
assign x_26033 = v_1768 | ~v_1570;
assign x_26034 = v_1768 | ~v_1571;
assign x_26035 = v_1768 | ~v_1760;
assign x_26036 = v_1768 | ~v_1761;
assign x_26037 = v_1768 | ~v_1762;
assign x_26038 = v_1768 | ~v_1763;
assign x_26039 = v_1768 | ~v_1572;
assign x_26040 = v_1768 | ~v_1573;
assign x_26041 = v_1768 | ~v_1574;
assign x_26042 = v_1768 | ~v_1575;
assign x_26043 = v_1768 | ~v_1576;
assign x_26044 = v_1768 | ~v_1579;
assign x_26045 = v_1768 | ~v_1764;
assign x_26046 = v_1768 | ~v_1765;
assign x_26047 = v_1768 | ~v_1766;
assign x_26048 = v_1768 | ~v_1767;
assign x_26049 = v_1768 | ~v_1582;
assign x_26050 = v_1768 | ~v_1583;
assign x_26051 = v_1768 | ~v_1584;
assign x_26052 = v_1768 | ~v_1585;
assign x_26053 = v_1768 | ~v_1586;
assign x_26054 = v_1768 | ~v_1589;
assign x_26055 = v_1768 | ~v_945;
assign x_26056 = v_1768 | ~v_946;
assign x_26057 = v_1768 | ~v_1105;
assign x_26058 = v_1768 | ~v_1106;
assign x_26059 = v_1768 | ~v_1055;
assign x_26060 = v_1768 | ~v_1056;
assign x_26061 = v_1768 | ~v_1107;
assign x_26062 = v_1768 | ~v_1108;
assign x_26063 = v_1768 | ~v_182;
assign x_26064 = v_1768 | ~v_163;
assign x_26065 = v_1768 | ~v_162;
assign x_26066 = v_1768 | ~v_161;
assign x_26067 = v_1768 | ~v_138;
assign x_26068 = v_1768 | ~v_137;
assign x_26069 = v_1768 | ~v_135;
assign x_26070 = v_1768 | ~v_134;
assign x_26071 = v_1768 | ~v_18;
assign x_26072 = v_1768 | ~v_16;
assign x_26073 = v_1768 | ~v_15;
assign x_26074 = v_1768 | ~v_12;
assign x_26075 = ~v_44 | ~v_173 | v_1767;
assign x_26076 = ~v_41 | ~v_174 | v_1766;
assign x_26077 = ~v_29 | v_173 | v_1765;
assign x_26078 = ~v_26 | v_174 | v_1764;
assign x_26079 = ~v_43 | ~v_175 | v_1763;
assign x_26080 = ~v_37 | ~v_176 | v_1762;
assign x_26081 = ~v_28 | v_175 | v_1761;
assign x_26082 = ~v_22 | v_176 | v_1760;
assign x_26083 = ~v_1758 | ~v_1757 | ~v_1756 | v_1759;
assign x_26084 = v_1758 | ~v_1618;
assign x_26085 = v_1758 | ~v_1619;
assign x_26086 = v_1758 | ~v_1620;
assign x_26087 = v_1758 | ~v_1621;
assign x_26088 = v_1758 | ~v_1690;
assign x_26089 = v_1758 | ~v_1691;
assign x_26090 = v_1758 | ~v_1692;
assign x_26091 = v_1758 | ~v_1693;
assign x_26092 = v_1758 | ~v_1626;
assign x_26093 = v_1758 | ~v_1627;
assign x_26094 = v_1758 | ~v_1628;
assign x_26095 = v_1758 | ~v_1629;
assign x_26096 = v_1758 | ~v_1630;
assign x_26097 = v_1758 | ~v_1631;
assign x_26098 = v_1758 | ~v_1694;
assign x_26099 = v_1758 | ~v_1695;
assign x_26100 = v_1758 | ~v_1696;
assign x_26101 = v_1758 | ~v_1697;
assign x_26102 = v_1758 | ~v_1636;
assign x_26103 = v_1758 | ~v_1637;
assign x_26104 = v_1758 | ~v_1638;
assign x_26105 = v_1758 | ~v_1639;
assign x_26106 = v_1758 | ~v_1640;
assign x_26107 = v_1758 | ~v_1641;
assign x_26108 = v_1758 | ~v_1037;
assign x_26109 = v_1758 | ~v_1038;
assign x_26110 = v_1758 | ~v_1039;
assign x_26111 = v_1758 | ~v_1040;
assign x_26112 = v_1758 | ~v_927;
assign x_26113 = v_1758 | ~v_928;
assign x_26114 = v_1758 | ~v_839;
assign x_26115 = v_1758 | ~v_840;
assign x_26116 = v_1758 | ~v_184;
assign x_26117 = v_1758 | ~v_170;
assign x_26118 = v_1758 | ~v_169;
assign x_26119 = v_1758 | ~v_151;
assign x_26120 = v_1758 | ~v_150;
assign x_26121 = v_1758 | ~v_149;
assign x_26122 = v_1758 | ~v_148;
assign x_26123 = v_1758 | ~v_147;
assign x_26124 = v_1758 | ~v_103;
assign x_26125 = v_1758 | ~v_101;
assign x_26126 = v_1758 | ~v_100;
assign x_26127 = v_1758 | ~v_98;
assign x_26128 = v_1757 | ~v_1593;
assign x_26129 = v_1757 | ~v_1594;
assign x_26130 = v_1757 | ~v_1595;
assign x_26131 = v_1757 | ~v_1596;
assign x_26132 = v_1757 | ~v_1681;
assign x_26133 = v_1757 | ~v_1682;
assign x_26134 = v_1757 | ~v_1683;
assign x_26135 = v_1757 | ~v_1684;
assign x_26136 = v_1757 | ~v_1601;
assign x_26137 = v_1757 | ~v_1602;
assign x_26138 = v_1757 | ~v_1603;
assign x_26139 = v_1757 | ~v_1604;
assign x_26140 = v_1757 | ~v_1605;
assign x_26141 = v_1757 | ~v_1606;
assign x_26142 = v_1757 | ~v_1685;
assign x_26143 = v_1757 | ~v_1686;
assign x_26144 = v_1757 | ~v_1687;
assign x_26145 = v_1757 | ~v_1688;
assign x_26146 = v_1757 | ~v_1611;
assign x_26147 = v_1757 | ~v_1612;
assign x_26148 = v_1757 | ~v_1613;
assign x_26149 = v_1757 | ~v_1614;
assign x_26150 = v_1757 | ~v_1615;
assign x_26151 = v_1757 | ~v_1616;
assign x_26152 = v_1757 | ~v_1032;
assign x_26153 = v_1757 | ~v_1033;
assign x_26154 = v_1757 | ~v_1034;
assign x_26155 = v_1757 | ~v_1035;
assign x_26156 = v_1757 | ~v_912;
assign x_26157 = v_1757 | ~v_913;
assign x_26158 = v_1757 | ~v_806;
assign x_26159 = v_1757 | ~v_807;
assign x_26160 = v_1757 | ~v_183;
assign x_26161 = v_1757 | ~v_166;
assign x_26162 = v_1757 | ~v_165;
assign x_26163 = v_1757 | ~v_146;
assign x_26164 = v_1757 | ~v_145;
assign x_26165 = v_1757 | ~v_144;
assign x_26166 = v_1757 | ~v_143;
assign x_26167 = v_1757 | ~v_142;
assign x_26168 = v_1757 | ~v_61;
assign x_26169 = v_1757 | ~v_59;
assign x_26170 = v_1757 | ~v_58;
assign x_26171 = v_1757 | ~v_56;
assign x_26172 = v_1756 | ~v_1568;
assign x_26173 = v_1756 | ~v_1569;
assign x_26174 = v_1756 | ~v_1570;
assign x_26175 = v_1756 | ~v_1571;
assign x_26176 = v_1756 | ~v_1672;
assign x_26177 = v_1756 | ~v_1673;
assign x_26178 = v_1756 | ~v_1674;
assign x_26179 = v_1756 | ~v_1675;
assign x_26180 = v_1756 | ~v_1576;
assign x_26181 = v_1756 | ~v_1577;
assign x_26182 = v_1756 | ~v_1578;
assign x_26183 = v_1756 | ~v_1579;
assign x_26184 = v_1756 | ~v_1580;
assign x_26185 = v_1756 | ~v_1581;
assign x_26186 = v_1756 | ~v_1676;
assign x_26187 = v_1756 | ~v_1677;
assign x_26188 = v_1756 | ~v_1678;
assign x_26189 = v_1756 | ~v_1679;
assign x_26190 = v_1756 | ~v_1586;
assign x_26191 = v_1756 | ~v_1587;
assign x_26192 = v_1756 | ~v_1588;
assign x_26193 = v_1756 | ~v_1589;
assign x_26194 = v_1756 | ~v_1590;
assign x_26195 = v_1756 | ~v_1591;
assign x_26196 = v_1756 | ~v_1027;
assign x_26197 = v_1756 | ~v_1028;
assign x_26198 = v_1756 | ~v_1029;
assign x_26199 = v_1756 | ~v_1030;
assign x_26200 = v_1756 | ~v_897;
assign x_26201 = v_1756 | ~v_898;
assign x_26202 = v_1756 | ~v_773;
assign x_26203 = v_1756 | ~v_774;
assign x_26204 = v_1756 | ~v_182;
assign x_26205 = v_1756 | ~v_162;
assign x_26206 = v_1756 | ~v_161;
assign x_26207 = v_1756 | ~v_138;
assign x_26208 = v_1756 | ~v_137;
assign x_26209 = v_1756 | ~v_136;
assign x_26210 = v_1756 | ~v_135;
assign x_26211 = v_1756 | ~v_134;
assign x_26212 = v_1756 | ~v_18;
assign x_26213 = v_1756 | ~v_16;
assign x_26214 = v_1756 | ~v_15;
assign x_26215 = v_1756 | ~v_13;
assign x_26216 = ~v_1754 | ~v_1745 | ~v_1736 | v_1755;
assign x_26217 = v_1754 | ~v_1618;
assign x_26218 = v_1754 | ~v_1619;
assign x_26219 = v_1754 | ~v_1620;
assign x_26220 = v_1754 | ~v_1621;
assign x_26221 = v_1754 | ~v_1662;
assign x_26222 = v_1754 | ~v_1663;
assign x_26223 = v_1754 | ~v_1664;
assign x_26224 = v_1754 | ~v_1665;
assign x_26225 = v_1754 | ~v_1626;
assign x_26226 = v_1754 | ~v_1746;
assign x_26227 = v_1754 | ~v_1747;
assign x_26228 = v_1754 | ~v_1629;
assign x_26229 = v_1754 | ~v_1748;
assign x_26230 = v_1754 | ~v_1749;
assign x_26231 = v_1754 | ~v_1666;
assign x_26232 = v_1754 | ~v_1667;
assign x_26233 = v_1754 | ~v_1668;
assign x_26234 = v_1754 | ~v_1669;
assign x_26235 = v_1754 | ~v_1636;
assign x_26236 = v_1754 | ~v_1750;
assign x_26237 = v_1754 | ~v_1751;
assign x_26238 = v_1754 | ~v_1639;
assign x_26239 = v_1754 | ~v_1752;
assign x_26240 = v_1754 | ~v_1753;
assign x_26241 = v_1754 | ~v_1193;
assign x_26242 = v_1754 | ~v_1241;
assign x_26243 = v_1754 | ~v_1194;
assign x_26244 = v_1754 | ~v_1242;
assign x_26245 = v_1754 | ~v_1023;
assign x_26246 = v_1754 | ~v_1024;
assign x_26247 = v_1754 | ~v_1243;
assign x_26248 = v_1754 | ~v_1244;
assign x_26249 = v_1754 | ~v_184;
assign x_26250 = v_1754 | ~v_171;
assign x_26251 = v_1754 | ~v_169;
assign x_26252 = v_1754 | ~v_149;
assign x_26253 = v_1754 | ~v_148;
assign x_26254 = v_1754 | ~v_147;
assign x_26255 = v_1754 | ~v_103;
assign x_26256 = v_1754 | ~v_102;
assign x_26257 = v_1754 | ~v_101;
assign x_26258 = v_1754 | ~v_100;
assign x_26259 = v_1754 | ~v_99;
assign x_26260 = v_1754 | ~v_94;
assign x_26261 = ~v_131 | ~v_152 | v_1753;
assign x_26262 = ~v_126 | ~v_153 | v_1752;
assign x_26263 = ~v_116 | v_152 | v_1751;
assign x_26264 = ~v_111 | v_153 | v_1750;
assign x_26265 = ~v_130 | ~v_156 | v_1749;
assign x_26266 = ~v_122 | ~v_157 | v_1748;
assign x_26267 = ~v_115 | v_156 | v_1747;
assign x_26268 = ~v_107 | v_157 | v_1746;
assign x_26269 = v_1745 | ~v_1593;
assign x_26270 = v_1745 | ~v_1594;
assign x_26271 = v_1745 | ~v_1595;
assign x_26272 = v_1745 | ~v_1596;
assign x_26273 = v_1745 | ~v_1653;
assign x_26274 = v_1745 | ~v_1654;
assign x_26275 = v_1745 | ~v_1655;
assign x_26276 = v_1745 | ~v_1656;
assign x_26277 = v_1745 | ~v_1601;
assign x_26278 = v_1745 | ~v_1737;
assign x_26279 = v_1745 | ~v_1738;
assign x_26280 = v_1745 | ~v_1604;
assign x_26281 = v_1745 | ~v_1739;
assign x_26282 = v_1745 | ~v_1740;
assign x_26283 = v_1745 | ~v_1657;
assign x_26284 = v_1745 | ~v_1658;
assign x_26285 = v_1745 | ~v_1659;
assign x_26286 = v_1745 | ~v_1660;
assign x_26287 = v_1745 | ~v_1611;
assign x_26288 = v_1745 | ~v_1741;
assign x_26289 = v_1745 | ~v_1742;
assign x_26290 = v_1745 | ~v_1614;
assign x_26291 = v_1745 | ~v_1743;
assign x_26292 = v_1745 | ~v_1744;
assign x_26293 = v_1745 | ~v_1178;
assign x_26294 = v_1745 | ~v_1236;
assign x_26295 = v_1745 | ~v_1179;
assign x_26296 = v_1745 | ~v_1237;
assign x_26297 = v_1745 | ~v_1008;
assign x_26298 = v_1745 | ~v_1009;
assign x_26299 = v_1745 | ~v_1238;
assign x_26300 = v_1745 | ~v_1239;
assign x_26301 = v_1745 | ~v_183;
assign x_26302 = v_1745 | ~v_167;
assign x_26303 = v_1745 | ~v_165;
assign x_26304 = v_1745 | ~v_144;
assign x_26305 = v_1745 | ~v_143;
assign x_26306 = v_1745 | ~v_142;
assign x_26307 = v_1745 | ~v_61;
assign x_26308 = v_1745 | ~v_60;
assign x_26309 = v_1745 | ~v_59;
assign x_26310 = v_1745 | ~v_58;
assign x_26311 = v_1745 | ~v_57;
assign x_26312 = v_1745 | ~v_52;
assign x_26313 = ~v_89 | ~v_152 | v_1744;
assign x_26314 = ~v_84 | ~v_153 | v_1743;
assign x_26315 = ~v_74 | v_152 | v_1742;
assign x_26316 = ~v_69 | v_153 | v_1741;
assign x_26317 = ~v_88 | ~v_156 | v_1740;
assign x_26318 = ~v_80 | ~v_157 | v_1739;
assign x_26319 = ~v_73 | v_156 | v_1738;
assign x_26320 = ~v_65 | v_157 | v_1737;
assign x_26321 = v_1736 | ~v_1568;
assign x_26322 = v_1736 | ~v_1569;
assign x_26323 = v_1736 | ~v_1570;
assign x_26324 = v_1736 | ~v_1571;
assign x_26325 = v_1736 | ~v_1644;
assign x_26326 = v_1736 | ~v_1645;
assign x_26327 = v_1736 | ~v_1646;
assign x_26328 = v_1736 | ~v_1647;
assign x_26329 = v_1736 | ~v_1576;
assign x_26330 = v_1736 | ~v_1728;
assign x_26331 = v_1736 | ~v_1729;
assign x_26332 = v_1736 | ~v_1579;
assign x_26333 = v_1736 | ~v_1730;
assign x_26334 = v_1736 | ~v_1731;
assign x_26335 = v_1736 | ~v_1648;
assign x_26336 = v_1736 | ~v_1649;
assign x_26337 = v_1736 | ~v_1650;
assign x_26338 = v_1736 | ~v_1651;
assign x_26339 = v_1736 | ~v_1586;
assign x_26340 = v_1736 | ~v_1732;
assign x_26341 = v_1736 | ~v_1733;
assign x_26342 = v_1736 | ~v_1589;
assign x_26343 = v_1736 | ~v_1734;
assign x_26344 = v_1736 | ~v_1735;
assign x_26345 = v_1736 | ~v_1163;
assign x_26346 = v_1736 | ~v_1231;
assign x_26347 = v_1736 | ~v_1164;
assign x_26348 = v_1736 | ~v_1232;
assign x_26349 = v_1736 | ~v_1233;
assign x_26350 = v_1736 | ~v_1234;
assign x_26351 = v_1736 | ~v_182;
assign x_26352 = v_1736 | ~v_163;
assign x_26353 = v_1736 | ~v_161;
assign x_26354 = v_1736 | ~v_136;
assign x_26355 = v_1736 | ~v_135;
assign x_26356 = v_1736 | ~v_134;
assign x_26357 = v_1736 | ~v_993;
assign x_26358 = v_1736 | ~v_994;
assign x_26359 = v_1736 | ~v_18;
assign x_26360 = v_1736 | ~v_17;
assign x_26361 = v_1736 | ~v_16;
assign x_26362 = v_1736 | ~v_15;
assign x_26363 = v_1736 | ~v_14;
assign x_26364 = v_1736 | ~v_9;
assign x_26365 = ~v_47 | ~v_152 | v_1735;
assign x_26366 = ~v_42 | ~v_153 | v_1734;
assign x_26367 = ~v_32 | v_152 | v_1733;
assign x_26368 = ~v_27 | v_153 | v_1732;
assign x_26369 = ~v_46 | ~v_156 | v_1731;
assign x_26370 = ~v_38 | ~v_157 | v_1730;
assign x_26371 = ~v_31 | v_156 | v_1729;
assign x_26372 = ~v_23 | v_157 | v_1728;
assign x_26373 = ~v_1726 | ~v_1717 | ~v_1708 | v_1727;
assign x_26374 = v_1726 | ~v_1618;
assign x_26375 = v_1726 | ~v_1619;
assign x_26376 = v_1726 | ~v_1620;
assign x_26377 = v_1726 | ~v_1621;
assign x_26378 = v_1726 | ~v_1662;
assign x_26379 = v_1726 | ~v_1663;
assign x_26380 = v_1726 | ~v_1664;
assign x_26381 = v_1726 | ~v_1665;
assign x_26382 = v_1726 | ~v_1718;
assign x_26383 = v_1726 | ~v_1719;
assign x_26384 = v_1726 | ~v_1720;
assign x_26385 = v_1726 | ~v_1721;
assign x_26386 = v_1726 | ~v_1626;
assign x_26387 = v_1726 | ~v_1629;
assign x_26388 = v_1726 | ~v_1722;
assign x_26389 = v_1726 | ~v_1723;
assign x_26390 = v_1726 | ~v_1724;
assign x_26391 = v_1726 | ~v_1725;
assign x_26392 = v_1726 | ~v_1666;
assign x_26393 = v_1726 | ~v_1667;
assign x_26394 = v_1726 | ~v_1668;
assign x_26395 = v_1726 | ~v_1669;
assign x_26396 = v_1726 | ~v_1636;
assign x_26397 = v_1726 | ~v_1639;
assign x_26398 = v_1726 | ~v_1191;
assign x_26399 = v_1726 | ~v_1192;
assign x_26400 = v_1726 | ~v_1193;
assign x_26401 = v_1726 | ~v_1194;
assign x_26402 = v_1726 | ~v_837;
assign x_26403 = v_1726 | ~v_838;
assign x_26404 = v_1726 | ~v_1195;
assign x_26405 = v_1726 | ~v_1196;
assign x_26406 = v_1726 | ~v_184;
assign x_26407 = v_1726 | ~v_171;
assign x_26408 = v_1726 | ~v_169;
assign x_26409 = v_1726 | ~v_160;
assign x_26410 = v_1726 | ~v_151;
assign x_26411 = v_1726 | ~v_150;
assign x_26412 = v_1726 | ~v_149;
assign x_26413 = v_1726 | ~v_147;
assign x_26414 = v_1726 | ~v_103;
assign x_26415 = v_1726 | ~v_100;
assign x_26416 = v_1726 | ~v_96;
assign x_26417 = v_1726 | ~v_94;
assign x_26418 = ~v_131 | ~v_178 | v_1725;
assign x_26419 = ~v_126 | ~v_177 | v_1724;
assign x_26420 = ~v_116 | v_178 | v_1723;
assign x_26421 = ~v_111 | v_177 | v_1722;
assign x_26422 = ~v_130 | ~v_158 | v_1721;
assign x_26423 = ~v_122 | ~v_158 | v_1720;
assign x_26424 = ~v_115 | v_158 | v_1719;
assign x_26425 = ~v_107 | v_158 | v_1718;
assign x_26426 = v_1717 | ~v_1593;
assign x_26427 = v_1717 | ~v_1594;
assign x_26428 = v_1717 | ~v_1595;
assign x_26429 = v_1717 | ~v_1596;
assign x_26430 = v_1717 | ~v_1653;
assign x_26431 = v_1717 | ~v_1654;
assign x_26432 = v_1717 | ~v_1655;
assign x_26433 = v_1717 | ~v_1656;
assign x_26434 = v_1717 | ~v_1709;
assign x_26435 = v_1717 | ~v_1710;
assign x_26436 = v_1717 | ~v_1711;
assign x_26437 = v_1717 | ~v_1712;
assign x_26438 = v_1717 | ~v_1601;
assign x_26439 = v_1717 | ~v_1604;
assign x_26440 = v_1717 | ~v_1713;
assign x_26441 = v_1717 | ~v_1714;
assign x_26442 = v_1717 | ~v_1715;
assign x_26443 = v_1717 | ~v_1716;
assign x_26444 = v_1717 | ~v_1657;
assign x_26445 = v_1717 | ~v_1658;
assign x_26446 = v_1717 | ~v_1659;
assign x_26447 = v_1717 | ~v_1660;
assign x_26448 = v_1717 | ~v_1611;
assign x_26449 = v_1717 | ~v_1614;
assign x_26450 = v_1717 | ~v_1176;
assign x_26451 = v_1717 | ~v_1177;
assign x_26452 = v_1717 | ~v_1178;
assign x_26453 = v_1717 | ~v_1179;
assign x_26454 = v_1717 | ~v_804;
assign x_26455 = v_1717 | ~v_805;
assign x_26456 = v_1717 | ~v_1180;
assign x_26457 = v_1717 | ~v_1181;
assign x_26458 = v_1717 | ~v_183;
assign x_26459 = v_1717 | ~v_167;
assign x_26460 = v_1717 | ~v_165;
assign x_26461 = v_1717 | ~v_159;
assign x_26462 = v_1717 | ~v_146;
assign x_26463 = v_1717 | ~v_145;
assign x_26464 = v_1717 | ~v_144;
assign x_26465 = v_1717 | ~v_142;
assign x_26466 = v_1717 | ~v_61;
assign x_26467 = v_1717 | ~v_58;
assign x_26468 = v_1717 | ~v_54;
assign x_26469 = v_1717 | ~v_52;
assign x_26470 = ~v_89 | ~v_178 | v_1716;
assign x_26471 = ~v_84 | ~v_177 | v_1715;
assign x_26472 = ~v_74 | v_178 | v_1714;
assign x_26473 = ~v_69 | v_177 | v_1713;
assign x_26474 = ~v_88 | ~v_158 | v_1712;
assign x_26475 = ~v_80 | ~v_158 | v_1711;
assign x_26476 = ~v_73 | v_158 | v_1710;
assign x_26477 = ~v_65 | v_158 | v_1709;
assign x_26478 = v_1708 | ~v_1568;
assign x_26479 = v_1708 | ~v_1569;
assign x_26480 = v_1708 | ~v_1570;
assign x_26481 = v_1708 | ~v_1571;
assign x_26482 = v_1708 | ~v_1644;
assign x_26483 = v_1708 | ~v_1645;
assign x_26484 = v_1708 | ~v_1646;
assign x_26485 = v_1708 | ~v_1647;
assign x_26486 = v_1708 | ~v_1700;
assign x_26487 = v_1708 | ~v_1701;
assign x_26488 = v_1708 | ~v_1702;
assign x_26489 = v_1708 | ~v_1703;
assign x_26490 = v_1708 | ~v_1576;
assign x_26491 = v_1708 | ~v_1579;
assign x_26492 = v_1708 | ~v_1704;
assign x_26493 = v_1708 | ~v_1705;
assign x_26494 = v_1708 | ~v_1706;
assign x_26495 = v_1708 | ~v_1707;
assign x_26496 = v_1708 | ~v_1648;
assign x_26497 = v_1708 | ~v_1649;
assign x_26498 = v_1708 | ~v_1650;
assign x_26499 = v_1708 | ~v_1651;
assign x_26500 = v_1708 | ~v_1586;
assign x_26501 = v_1708 | ~v_1589;
assign x_26502 = v_1708 | ~v_1161;
assign x_26503 = v_1708 | ~v_1162;
assign x_26504 = v_1708 | ~v_1163;
assign x_26505 = v_1708 | ~v_1164;
assign x_26506 = v_1708 | ~v_771;
assign x_26507 = v_1708 | ~v_772;
assign x_26508 = v_1708 | ~v_1165;
assign x_26509 = v_1708 | ~v_1166;
assign x_26510 = v_1708 | ~v_182;
assign x_26511 = v_1708 | ~v_163;
assign x_26512 = v_1708 | ~v_161;
assign x_26513 = v_1708 | ~v_155;
assign x_26514 = v_1708 | ~v_138;
assign x_26515 = v_1708 | ~v_137;
assign x_26516 = v_1708 | ~v_136;
assign x_26517 = v_1708 | ~v_134;
assign x_26518 = v_1708 | ~v_18;
assign x_26519 = v_1708 | ~v_15;
assign x_26520 = v_1708 | ~v_11;
assign x_26521 = v_1708 | ~v_9;
assign x_26522 = ~v_47 | ~v_178 | v_1707;
assign x_26523 = ~v_42 | ~v_177 | v_1706;
assign x_26524 = ~v_32 | v_178 | v_1705;
assign x_26525 = ~v_27 | v_177 | v_1704;
assign x_26526 = ~v_46 | ~v_158 | v_1703;
assign x_26527 = ~v_38 | ~v_158 | v_1702;
assign x_26528 = ~v_31 | v_158 | v_1701;
assign x_26529 = ~v_23 | v_158 | v_1700;
assign x_26530 = ~v_1698 | ~v_1689 | ~v_1680 | v_1699;
assign x_26531 = v_1698 | ~v_1618;
assign x_26532 = v_1698 | ~v_1619;
assign x_26533 = v_1698 | ~v_1620;
assign x_26534 = v_1698 | ~v_1621;
assign x_26535 = v_1698 | ~v_1662;
assign x_26536 = v_1698 | ~v_1663;
assign x_26537 = v_1698 | ~v_1664;
assign x_26538 = v_1698 | ~v_1665;
assign x_26539 = v_1698 | ~v_1690;
assign x_26540 = v_1698 | ~v_1691;
assign x_26541 = v_1698 | ~v_1692;
assign x_26542 = v_1698 | ~v_1693;
assign x_26543 = v_1698 | ~v_1626;
assign x_26544 = v_1698 | ~v_1629;
assign x_26545 = v_1698 | ~v_1694;
assign x_26546 = v_1698 | ~v_1695;
assign x_26547 = v_1698 | ~v_1696;
assign x_26548 = v_1698 | ~v_1697;
assign x_26549 = v_1698 | ~v_1666;
assign x_26550 = v_1698 | ~v_1667;
assign x_26551 = v_1698 | ~v_1668;
assign x_26552 = v_1698 | ~v_1669;
assign x_26553 = v_1698 | ~v_1636;
assign x_26554 = v_1698 | ~v_1639;
assign x_26555 = v_1698 | ~v_1209;
assign x_26556 = v_1698 | ~v_1210;
assign x_26557 = v_1698 | ~v_1193;
assign x_26558 = v_1698 | ~v_1194;
assign x_26559 = v_1698 | ~v_927;
assign x_26560 = v_1698 | ~v_928;
assign x_26561 = v_1698 | ~v_1211;
assign x_26562 = v_1698 | ~v_1212;
assign x_26563 = v_1698 | ~v_184;
assign x_26564 = v_1698 | ~v_172;
assign x_26565 = v_1698 | ~v_171;
assign x_26566 = v_1698 | ~v_169;
assign x_26567 = v_1698 | ~v_150;
assign x_26568 = v_1698 | ~v_149;
assign x_26569 = v_1698 | ~v_148;
assign x_26570 = v_1698 | ~v_147;
assign x_26571 = v_1698 | ~v_102;
assign x_26572 = v_1698 | ~v_101;
assign x_26573 = v_1698 | ~v_100;
assign x_26574 = v_1698 | ~v_94;
assign x_26575 = ~v_131 | ~v_173 | v_1697;
assign x_26576 = ~v_126 | ~v_174 | v_1696;
assign x_26577 = ~v_116 | v_173 | v_1695;
assign x_26578 = ~v_111 | v_174 | v_1694;
assign x_26579 = ~v_130 | ~v_175 | v_1693;
assign x_26580 = ~v_122 | ~v_176 | v_1692;
assign x_26581 = ~v_115 | v_175 | v_1691;
assign x_26582 = ~v_107 | v_176 | v_1690;
assign x_26583 = v_1689 | ~v_1593;
assign x_26584 = v_1689 | ~v_1594;
assign x_26585 = v_1689 | ~v_1595;
assign x_26586 = v_1689 | ~v_1596;
assign x_26587 = v_1689 | ~v_1653;
assign x_26588 = v_1689 | ~v_1654;
assign x_26589 = v_1689 | ~v_1655;
assign x_26590 = v_1689 | ~v_1656;
assign x_26591 = v_1689 | ~v_1681;
assign x_26592 = v_1689 | ~v_1682;
assign x_26593 = v_1689 | ~v_1683;
assign x_26594 = v_1689 | ~v_1684;
assign x_26595 = v_1689 | ~v_1601;
assign x_26596 = v_1689 | ~v_1604;
assign x_26597 = v_1689 | ~v_1685;
assign x_26598 = v_1689 | ~v_1686;
assign x_26599 = v_1689 | ~v_1687;
assign x_26600 = v_1689 | ~v_1688;
assign x_26601 = v_1689 | ~v_1657;
assign x_26602 = v_1689 | ~v_1658;
assign x_26603 = v_1689 | ~v_1659;
assign x_26604 = v_1689 | ~v_1660;
assign x_26605 = v_1689 | ~v_1611;
assign x_26606 = v_1689 | ~v_1614;
assign x_26607 = v_1689 | ~v_1204;
assign x_26608 = v_1689 | ~v_1205;
assign x_26609 = v_1689 | ~v_1178;
assign x_26610 = v_1689 | ~v_1179;
assign x_26611 = v_1689 | ~v_912;
assign x_26612 = v_1689 | ~v_913;
assign x_26613 = v_1689 | ~v_1206;
assign x_26614 = v_1689 | ~v_1207;
assign x_26615 = v_1689 | ~v_183;
assign x_26616 = v_1689 | ~v_168;
assign x_26617 = v_1689 | ~v_167;
assign x_26618 = v_1689 | ~v_165;
assign x_26619 = v_1689 | ~v_145;
assign x_26620 = v_1689 | ~v_144;
assign x_26621 = v_1689 | ~v_143;
assign x_26622 = v_1689 | ~v_142;
assign x_26623 = v_1689 | ~v_60;
assign x_26624 = v_1689 | ~v_59;
assign x_26625 = v_1689 | ~v_58;
assign x_26626 = v_1689 | ~v_52;
assign x_26627 = ~v_89 | ~v_173 | v_1688;
assign x_26628 = ~v_84 | ~v_174 | v_1687;
assign x_26629 = ~v_74 | v_173 | v_1686;
assign x_26630 = ~v_69 | v_174 | v_1685;
assign x_26631 = ~v_88 | ~v_175 | v_1684;
assign x_26632 = ~v_80 | ~v_176 | v_1683;
assign x_26633 = ~v_73 | v_175 | v_1682;
assign x_26634 = ~v_65 | v_176 | v_1681;
assign x_26635 = v_1680 | ~v_1568;
assign x_26636 = v_1680 | ~v_1569;
assign x_26637 = v_1680 | ~v_1570;
assign x_26638 = v_1680 | ~v_1571;
assign x_26639 = v_1680 | ~v_1644;
assign x_26640 = v_1680 | ~v_1645;
assign x_26641 = v_1680 | ~v_1646;
assign x_26642 = v_1680 | ~v_1647;
assign x_26643 = v_1680 | ~v_1672;
assign x_26644 = v_1680 | ~v_1673;
assign x_26645 = v_1680 | ~v_1674;
assign x_26646 = v_1680 | ~v_1675;
assign x_26647 = v_1680 | ~v_1576;
assign x_26648 = v_1680 | ~v_1579;
assign x_26649 = v_1680 | ~v_1676;
assign x_26650 = v_1680 | ~v_1677;
assign x_26651 = v_1680 | ~v_1678;
assign x_26652 = v_1680 | ~v_1679;
assign x_26653 = v_1680 | ~v_1648;
assign x_26654 = v_1680 | ~v_1649;
assign x_26655 = v_1680 | ~v_1650;
assign x_26656 = v_1680 | ~v_1651;
assign x_26657 = v_1680 | ~v_1586;
assign x_26658 = v_1680 | ~v_1589;
assign x_26659 = v_1680 | ~v_1199;
assign x_26660 = v_1680 | ~v_1200;
assign x_26661 = v_1680 | ~v_1163;
assign x_26662 = v_1680 | ~v_1164;
assign x_26663 = v_1680 | ~v_897;
assign x_26664 = v_1680 | ~v_898;
assign x_26665 = v_1680 | ~v_1201;
assign x_26666 = v_1680 | ~v_1202;
assign x_26667 = v_1680 | ~v_182;
assign x_26668 = v_1680 | ~v_164;
assign x_26669 = v_1680 | ~v_163;
assign x_26670 = v_1680 | ~v_161;
assign x_26671 = v_1680 | ~v_137;
assign x_26672 = v_1680 | ~v_136;
assign x_26673 = v_1680 | ~v_135;
assign x_26674 = v_1680 | ~v_134;
assign x_26675 = v_1680 | ~v_17;
assign x_26676 = v_1680 | ~v_16;
assign x_26677 = v_1680 | ~v_15;
assign x_26678 = v_1680 | ~v_9;
assign x_26679 = ~v_47 | ~v_173 | v_1679;
assign x_26680 = ~v_42 | ~v_174 | v_1678;
assign x_26681 = ~v_32 | v_173 | v_1677;
assign x_26682 = ~v_27 | v_174 | v_1676;
assign x_26683 = ~v_46 | ~v_175 | v_1675;
assign x_26684 = ~v_38 | ~v_176 | v_1674;
assign x_26685 = ~v_31 | v_175 | v_1673;
assign x_26686 = ~v_23 | v_176 | v_1672;
assign x_26687 = ~v_1670 | ~v_1661 | ~v_1652 | v_1671;
assign x_26688 = v_1670 | ~v_1618;
assign x_26689 = v_1670 | ~v_1619;
assign x_26690 = v_1670 | ~v_1620;
assign x_26691 = v_1670 | ~v_1621;
assign x_26692 = v_1670 | ~v_1662;
assign x_26693 = v_1670 | ~v_1663;
assign x_26694 = v_1670 | ~v_1664;
assign x_26695 = v_1670 | ~v_1665;
assign x_26696 = v_1670 | ~v_1622;
assign x_26697 = v_1670 | ~v_1623;
assign x_26698 = v_1670 | ~v_1624;
assign x_26699 = v_1670 | ~v_1625;
assign x_26700 = v_1670 | ~v_1626;
assign x_26701 = v_1670 | ~v_1629;
assign x_26702 = v_1670 | ~v_1632;
assign x_26703 = v_1670 | ~v_1633;
assign x_26704 = v_1670 | ~v_1634;
assign x_26705 = v_1670 | ~v_1635;
assign x_26706 = v_1670 | ~v_1666;
assign x_26707 = v_1670 | ~v_1667;
assign x_26708 = v_1670 | ~v_1668;
assign x_26709 = v_1670 | ~v_1669;
assign x_26710 = v_1670 | ~v_1636;
assign x_26711 = v_1670 | ~v_1639;
assign x_26712 = v_1670 | ~v_1225;
assign x_26713 = v_1670 | ~v_1226;
assign x_26714 = v_1670 | ~v_1227;
assign x_26715 = v_1670 | ~v_1228;
assign x_26716 = v_1670 | ~v_1193;
assign x_26717 = v_1670 | ~v_1194;
assign x_26718 = v_1670 | ~v_975;
assign x_26719 = v_1670 | ~v_976;
assign x_26720 = v_1670 | ~v_184;
assign x_26721 = v_1670 | ~v_171;
assign x_26722 = v_1670 | ~v_169;
assign x_26723 = v_1670 | ~v_150;
assign x_26724 = v_1670 | ~v_148;
assign x_26725 = v_1670 | ~v_103;
assign x_26726 = v_1670 | ~v_102;
assign x_26727 = v_1670 | ~v_101;
assign x_26728 = v_1670 | ~v_100;
assign x_26729 = v_1670 | ~v_97;
assign x_26730 = v_1670 | ~v_95;
assign x_26731 = v_1670 | ~v_94;
assign x_26732 = ~v_128 | ~v_154 | v_1669;
assign x_26733 = ~v_125 | ~v_154 | v_1668;
assign x_26734 = ~v_113 | v_154 | v_1667;
assign x_26735 = ~v_110 | v_154 | v_1666;
assign x_26736 = ~v_127 | ~v_177 | v_1665;
assign x_26737 = ~v_121 | ~v_178 | v_1664;
assign x_26738 = ~v_112 | v_177 | v_1663;
assign x_26739 = ~v_106 | v_178 | v_1662;
assign x_26740 = v_1661 | ~v_1593;
assign x_26741 = v_1661 | ~v_1594;
assign x_26742 = v_1661 | ~v_1595;
assign x_26743 = v_1661 | ~v_1596;
assign x_26744 = v_1661 | ~v_1653;
assign x_26745 = v_1661 | ~v_1654;
assign x_26746 = v_1661 | ~v_1655;
assign x_26747 = v_1661 | ~v_1656;
assign x_26748 = v_1661 | ~v_1597;
assign x_26749 = v_1661 | ~v_1598;
assign x_26750 = v_1661 | ~v_1599;
assign x_26751 = v_1661 | ~v_1600;
assign x_26752 = v_1661 | ~v_1601;
assign x_26753 = v_1661 | ~v_1604;
assign x_26754 = v_1661 | ~v_1607;
assign x_26755 = v_1661 | ~v_1608;
assign x_26756 = v_1661 | ~v_1609;
assign x_26757 = v_1661 | ~v_1610;
assign x_26758 = v_1661 | ~v_1657;
assign x_26759 = v_1661 | ~v_1658;
assign x_26760 = v_1661 | ~v_1659;
assign x_26761 = v_1661 | ~v_1660;
assign x_26762 = v_1661 | ~v_1611;
assign x_26763 = v_1661 | ~v_1614;
assign x_26764 = v_1661 | ~v_1220;
assign x_26765 = v_1661 | ~v_1221;
assign x_26766 = v_1661 | ~v_1222;
assign x_26767 = v_1661 | ~v_1223;
assign x_26768 = v_1661 | ~v_1178;
assign x_26769 = v_1661 | ~v_1179;
assign x_26770 = v_1661 | ~v_960;
assign x_26771 = v_1661 | ~v_961;
assign x_26772 = v_1661 | ~v_183;
assign x_26773 = v_1661 | ~v_167;
assign x_26774 = v_1661 | ~v_165;
assign x_26775 = v_1661 | ~v_145;
assign x_26776 = v_1661 | ~v_143;
assign x_26777 = v_1661 | ~v_61;
assign x_26778 = v_1661 | ~v_60;
assign x_26779 = v_1661 | ~v_59;
assign x_26780 = v_1661 | ~v_58;
assign x_26781 = v_1661 | ~v_55;
assign x_26782 = v_1661 | ~v_53;
assign x_26783 = v_1661 | ~v_52;
assign x_26784 = ~v_86 | ~v_154 | v_1660;
assign x_26785 = ~v_83 | ~v_154 | v_1659;
assign x_26786 = ~v_71 | v_154 | v_1658;
assign x_26787 = ~v_68 | v_154 | v_1657;
assign x_26788 = ~v_85 | ~v_177 | v_1656;
assign x_26789 = ~v_79 | ~v_178 | v_1655;
assign x_26790 = ~v_70 | v_177 | v_1654;
assign x_26791 = ~v_64 | v_178 | v_1653;
assign x_26792 = v_1652 | ~v_1568;
assign x_26793 = v_1652 | ~v_1569;
assign x_26794 = v_1652 | ~v_1570;
assign x_26795 = v_1652 | ~v_1571;
assign x_26796 = v_1652 | ~v_1644;
assign x_26797 = v_1652 | ~v_1645;
assign x_26798 = v_1652 | ~v_1646;
assign x_26799 = v_1652 | ~v_1647;
assign x_26800 = v_1652 | ~v_1572;
assign x_26801 = v_1652 | ~v_1573;
assign x_26802 = v_1652 | ~v_1574;
assign x_26803 = v_1652 | ~v_1575;
assign x_26804 = v_1652 | ~v_1576;
assign x_26805 = v_1652 | ~v_1579;
assign x_26806 = v_1652 | ~v_1582;
assign x_26807 = v_1652 | ~v_1583;
assign x_26808 = v_1652 | ~v_1584;
assign x_26809 = v_1652 | ~v_1585;
assign x_26810 = v_1652 | ~v_1648;
assign x_26811 = v_1652 | ~v_1649;
assign x_26812 = v_1652 | ~v_1650;
assign x_26813 = v_1652 | ~v_1651;
assign x_26814 = v_1652 | ~v_1586;
assign x_26815 = v_1652 | ~v_1589;
assign x_26816 = v_1652 | ~v_1215;
assign x_26817 = v_1652 | ~v_1216;
assign x_26818 = v_1652 | ~v_1217;
assign x_26819 = v_1652 | ~v_1218;
assign x_26820 = v_1652 | ~v_1163;
assign x_26821 = v_1652 | ~v_1164;
assign x_26822 = v_1652 | ~v_945;
assign x_26823 = v_1652 | ~v_946;
assign x_26824 = v_1652 | ~v_182;
assign x_26825 = v_1652 | ~v_163;
assign x_26826 = v_1652 | ~v_161;
assign x_26827 = v_1652 | ~v_137;
assign x_26828 = v_1652 | ~v_135;
assign x_26829 = v_1652 | ~v_18;
assign x_26830 = v_1652 | ~v_17;
assign x_26831 = v_1652 | ~v_16;
assign x_26832 = v_1652 | ~v_15;
assign x_26833 = v_1652 | ~v_12;
assign x_26834 = v_1652 | ~v_10;
assign x_26835 = v_1652 | ~v_9;
assign x_26836 = ~v_44 | ~v_154 | v_1651;
assign x_26837 = ~v_41 | ~v_154 | v_1650;
assign x_26838 = ~v_29 | v_154 | v_1649;
assign x_26839 = ~v_26 | v_154 | v_1648;
assign x_26840 = ~v_43 | ~v_177 | v_1647;
assign x_26841 = ~v_37 | ~v_178 | v_1646;
assign x_26842 = ~v_28 | v_177 | v_1645;
assign x_26843 = ~v_22 | v_178 | v_1644;
assign x_26844 = ~v_1642 | ~v_1617 | ~v_1592 | v_1643;
assign x_26845 = v_1642 | ~v_1618;
assign x_26846 = v_1642 | ~v_1619;
assign x_26847 = v_1642 | ~v_1620;
assign x_26848 = v_1642 | ~v_1621;
assign x_26849 = v_1642 | ~v_1622;
assign x_26850 = v_1642 | ~v_1623;
assign x_26851 = v_1642 | ~v_1624;
assign x_26852 = v_1642 | ~v_1625;
assign x_26853 = v_1642 | ~v_1626;
assign x_26854 = v_1642 | ~v_1627;
assign x_26855 = v_1642 | ~v_1628;
assign x_26856 = v_1642 | ~v_1629;
assign x_26857 = v_1642 | ~v_1630;
assign x_26858 = v_1642 | ~v_1631;
assign x_26859 = v_1642 | ~v_1632;
assign x_26860 = v_1642 | ~v_1633;
assign x_26861 = v_1642 | ~v_1634;
assign x_26862 = v_1642 | ~v_1635;
assign x_26863 = v_1642 | ~v_1636;
assign x_26864 = v_1642 | ~v_1637;
assign x_26865 = v_1642 | ~v_1638;
assign x_26866 = v_1642 | ~v_1639;
assign x_26867 = v_1642 | ~v_1640;
assign x_26868 = v_1642 | ~v_1641;
assign x_26869 = v_1642 | ~v_1147;
assign x_26870 = v_1642 | ~v_1148;
assign x_26871 = v_1642 | ~v_975;
assign x_26872 = v_1642 | ~v_976;
assign x_26873 = v_1642 | ~v_839;
assign x_26874 = v_1642 | ~v_840;
assign x_26875 = v_1642 | ~v_1149;
assign x_26876 = v_1642 | ~v_1150;
assign x_26877 = v_1642 | ~v_184;
assign x_26878 = v_1642 | ~v_170;
assign x_26879 = v_1642 | ~v_169;
assign x_26880 = v_1642 | ~v_150;
assign x_26881 = v_1642 | ~v_148;
assign x_26882 = v_1642 | ~v_147;
assign x_26883 = v_1642 | ~v_103;
assign x_26884 = v_1642 | ~v_102;
assign x_26885 = v_1642 | ~v_101;
assign x_26886 = v_1642 | ~v_100;
assign x_26887 = v_1642 | ~v_98;
assign x_26888 = v_1642 | ~v_97;
assign x_26889 = ~v_128 | ~v_152 | v_1641;
assign x_26890 = ~v_125 | ~v_153 | v_1640;
assign x_26891 = ~v_124 | ~v_154 | v_1639;
assign x_26892 = ~v_113 | v_152 | v_1638;
assign x_26893 = ~v_110 | v_153 | v_1637;
assign x_26894 = ~v_109 | v_154 | v_1636;
assign x_26895 = ~v_131 | ~v_154 | v_1635;
assign x_26896 = ~v_126 | ~v_154 | v_1634;
assign x_26897 = ~v_116 | v_154 | v_1633;
assign x_26898 = ~v_111 | v_154 | v_1632;
assign x_26899 = ~v_127 | ~v_156 | v_1631;
assign x_26900 = ~v_121 | ~v_157 | v_1630;
assign x_26901 = ~v_119 | ~v_158 | v_1629;
assign x_26902 = ~v_112 | v_156 | v_1628;
assign x_26903 = ~v_106 | v_157 | v_1627;
assign x_26904 = ~v_104 | v_158 | v_1626;
assign x_26905 = ~v_130 | ~v_177 | v_1625;
assign x_26906 = ~v_122 | ~v_178 | v_1624;
assign x_26907 = ~v_115 | v_177 | v_1623;
assign x_26908 = ~v_107 | v_178 | v_1622;
assign x_26909 = ~v_123 | ~v_177 | v_1621;
assign x_26910 = ~v_120 | ~v_178 | v_1620;
assign x_26911 = ~v_108 | v_177 | v_1619;
assign x_26912 = ~v_105 | v_178 | v_1618;
assign x_26913 = v_1617 | ~v_1593;
assign x_26914 = v_1617 | ~v_1594;
assign x_26915 = v_1617 | ~v_1595;
assign x_26916 = v_1617 | ~v_1596;
assign x_26917 = v_1617 | ~v_1597;
assign x_26918 = v_1617 | ~v_1598;
assign x_26919 = v_1617 | ~v_1599;
assign x_26920 = v_1617 | ~v_1600;
assign x_26921 = v_1617 | ~v_1601;
assign x_26922 = v_1617 | ~v_1602;
assign x_26923 = v_1617 | ~v_1603;
assign x_26924 = v_1617 | ~v_1604;
assign x_26925 = v_1617 | ~v_1605;
assign x_26926 = v_1617 | ~v_1606;
assign x_26927 = v_1617 | ~v_1607;
assign x_26928 = v_1617 | ~v_1608;
assign x_26929 = v_1617 | ~v_1609;
assign x_26930 = v_1617 | ~v_1610;
assign x_26931 = v_1617 | ~v_1611;
assign x_26932 = v_1617 | ~v_1612;
assign x_26933 = v_1617 | ~v_1613;
assign x_26934 = v_1617 | ~v_1614;
assign x_26935 = v_1617 | ~v_1615;
assign x_26936 = v_1617 | ~v_1616;
assign x_26937 = v_1617 | ~v_1142;
assign x_26938 = v_1617 | ~v_1143;
assign x_26939 = v_1617 | ~v_960;
assign x_26940 = v_1617 | ~v_961;
assign x_26941 = v_1617 | ~v_806;
assign x_26942 = v_1617 | ~v_807;
assign x_26943 = v_1617 | ~v_1144;
assign x_26944 = v_1617 | ~v_1145;
assign x_26945 = v_1617 | ~v_183;
assign x_26946 = v_1617 | ~v_166;
assign x_26947 = v_1617 | ~v_165;
assign x_26948 = v_1617 | ~v_145;
assign x_26949 = v_1617 | ~v_143;
assign x_26950 = v_1617 | ~v_142;
assign x_26951 = v_1617 | ~v_61;
assign x_26952 = v_1617 | ~v_60;
assign x_26953 = v_1617 | ~v_59;
assign x_26954 = v_1617 | ~v_58;
assign x_26955 = v_1617 | ~v_56;
assign x_26956 = v_1617 | ~v_55;
assign x_26957 = ~v_86 | ~v_152 | v_1616;
assign x_26958 = ~v_83 | ~v_153 | v_1615;
assign x_26959 = ~v_82 | ~v_154 | v_1614;
assign x_26960 = ~v_71 | v_152 | v_1613;
assign x_26961 = ~v_68 | v_153 | v_1612;
assign x_26962 = ~v_67 | v_154 | v_1611;
assign x_26963 = ~v_89 | ~v_154 | v_1610;
assign x_26964 = ~v_84 | ~v_154 | v_1609;
assign x_26965 = ~v_74 | v_154 | v_1608;
assign x_26966 = ~v_69 | v_154 | v_1607;
assign x_26967 = ~v_85 | ~v_156 | v_1606;
assign x_26968 = ~v_79 | ~v_157 | v_1605;
assign x_26969 = ~v_77 | ~v_158 | v_1604;
assign x_26970 = ~v_70 | v_156 | v_1603;
assign x_26971 = ~v_64 | v_157 | v_1602;
assign x_26972 = ~v_62 | v_158 | v_1601;
assign x_26973 = ~v_88 | ~v_177 | v_1600;
assign x_26974 = ~v_80 | ~v_178 | v_1599;
assign x_26975 = ~v_73 | v_177 | v_1598;
assign x_26976 = ~v_65 | v_178 | v_1597;
assign x_26977 = ~v_81 | ~v_177 | v_1596;
assign x_26978 = ~v_78 | ~v_178 | v_1595;
assign x_26979 = ~v_66 | v_177 | v_1594;
assign x_26980 = ~v_63 | v_178 | v_1593;
assign x_26981 = v_1592 | ~v_1568;
assign x_26982 = v_1592 | ~v_1569;
assign x_26983 = v_1592 | ~v_1570;
assign x_26984 = v_1592 | ~v_1571;
assign x_26985 = v_1592 | ~v_1572;
assign x_26986 = v_1592 | ~v_1573;
assign x_26987 = v_1592 | ~v_1574;
assign x_26988 = v_1592 | ~v_1575;
assign x_26989 = v_1592 | ~v_1576;
assign x_26990 = v_1592 | ~v_1577;
assign x_26991 = v_1592 | ~v_1578;
assign x_26992 = v_1592 | ~v_1579;
assign x_26993 = v_1592 | ~v_1580;
assign x_26994 = v_1592 | ~v_1581;
assign x_26995 = v_1592 | ~v_1582;
assign x_26996 = v_1592 | ~v_1583;
assign x_26997 = v_1592 | ~v_1584;
assign x_26998 = v_1592 | ~v_1585;
assign x_26999 = v_1592 | ~v_1586;
assign x_27000 = v_1592 | ~v_1587;
assign x_27001 = v_1592 | ~v_1588;
assign x_27002 = v_1592 | ~v_1589;
assign x_27003 = v_1592 | ~v_1590;
assign x_27004 = v_1592 | ~v_1591;
assign x_27005 = v_1592 | ~v_1137;
assign x_27006 = v_1592 | ~v_1138;
assign x_27007 = v_1592 | ~v_945;
assign x_27008 = v_1592 | ~v_946;
assign x_27009 = v_1592 | ~v_773;
assign x_27010 = v_1592 | ~v_774;
assign x_27011 = v_1592 | ~v_1139;
assign x_27012 = v_1592 | ~v_1140;
assign x_27013 = v_1592 | ~v_182;
assign x_27014 = v_1592 | ~v_162;
assign x_27015 = v_1592 | ~v_161;
assign x_27016 = v_1592 | ~v_137;
assign x_27017 = v_1592 | ~v_135;
assign x_27018 = v_1592 | ~v_134;
assign x_27019 = v_1592 | ~v_18;
assign x_27020 = v_1592 | ~v_17;
assign x_27021 = v_1592 | ~v_16;
assign x_27022 = v_1592 | ~v_15;
assign x_27023 = v_1592 | ~v_13;
assign x_27024 = v_1592 | ~v_12;
assign x_27025 = ~v_44 | ~v_152 | v_1591;
assign x_27026 = ~v_41 | ~v_153 | v_1590;
assign x_27027 = ~v_40 | ~v_154 | v_1589;
assign x_27028 = ~v_29 | v_152 | v_1588;
assign x_27029 = ~v_26 | v_153 | v_1587;
assign x_27030 = ~v_25 | v_154 | v_1586;
assign x_27031 = ~v_47 | ~v_154 | v_1585;
assign x_27032 = ~v_42 | ~v_154 | v_1584;
assign x_27033 = ~v_32 | v_154 | v_1583;
assign x_27034 = ~v_27 | v_154 | v_1582;
assign x_27035 = ~v_43 | ~v_156 | v_1581;
assign x_27036 = ~v_37 | ~v_157 | v_1580;
assign x_27037 = ~v_35 | ~v_158 | v_1579;
assign x_27038 = ~v_28 | v_156 | v_1578;
assign x_27039 = ~v_22 | v_157 | v_1577;
assign x_27040 = ~v_20 | v_158 | v_1576;
assign x_27041 = ~v_46 | ~v_177 | v_1575;
assign x_27042 = ~v_38 | ~v_178 | v_1574;
assign x_27043 = ~v_31 | v_177 | v_1573;
assign x_27044 = ~v_23 | v_178 | v_1572;
assign x_27045 = ~v_39 | ~v_177 | v_1571;
assign x_27046 = ~v_36 | ~v_178 | v_1570;
assign x_27047 = ~v_24 | v_177 | v_1569;
assign x_27048 = ~v_21 | v_178 | v_1568;
assign x_27049 = v_1567 | ~v_1566;
assign x_27050 = v_1567 | ~v_727;
assign x_27051 = v_152 | v_153 | ~v_1565 | ~v_1564 | v_1566;
assign x_27052 = v_1565 | ~v_728;
assign x_27053 = v_1565 | ~v_731;
assign x_27054 = v_1564 | ~v_727;
assign x_27055 = v_1564 | ~v_730;
assign x_27056 = v_1563 | ~v_1562;
assign x_27057 = v_1563 | ~v_735;
assign x_27058 = v_174 | v_173 | ~v_1561 | ~v_1560 | v_1562;
assign x_27059 = v_1561 | ~v_737;
assign x_27060 = v_1561 | ~v_728;
assign x_27061 = v_1560 | ~v_735;
assign x_27062 = v_1560 | ~v_730;
assign x_27063 = ~v_725 | ~v_724 | ~v_723 | ~v_722 | ~v_1558 | ~v_1554 | ~v_1550 | ~v_1546 | ~v_1542 | ~v_1514 | ~v_1510 | ~v_1506 | ~v_1502 | ~v_1498 | ~v_1470 | ~v_1466 | ~v_1438 | ~v_1410 | ~v_1382 | ~v_1354 | ~v_1278 | v_1559;
assign x_27064 = v_1558 | ~v_1555;
assign x_27065 = v_1558 | ~v_1556;
assign x_27066 = v_1558 | ~v_1557;
assign x_27067 = v_98 | v_103 | v_101 | v_100 | v_95 | v_99 | v_102 | ~v_719 | ~v_718 | v_170 | v_169 | v_149 | v_148 | v_184 | ~v_483 | ~v_717 | ~v_299 | ~v_482 | ~v_716 | ~v_298 | ~v_1464 | ~v_1352 | ~v_1463 | ~v_1351 | ~v_1350 | ~v_1462 | ~v_1349 | ~v_1461 | ~v_1348 | ~v_1347 | ~v_1460 | ~v_1342 | ~v_1459 | ~v_1341 | ~v_1340 | ~v_1458 | ~v_1339 | ~v_1457 | ~v_1338 | ~v_1337 | ~v_1332 | ~v_1331 | ~v_1330 | ~v_1329 | v_1557;
assign x_27068 = v_53 | v_56 | v_61 | v_60 | v_59 | v_58 | v_57 | ~v_714 | ~v_713 | v_144 | v_143 | v_166 | v_165 | v_183 | ~v_266 | ~v_468 | ~v_712 | ~v_467 | ~v_711 | ~v_265 | ~v_1455 | ~v_1327 | ~v_1454 | ~v_1326 | ~v_1325 | ~v_1453 | ~v_1324 | ~v_1452 | ~v_1323 | ~v_1322 | ~v_1451 | ~v_1317 | ~v_1450 | ~v_1316 | ~v_1315 | ~v_1449 | ~v_1314 | ~v_1448 | ~v_1313 | ~v_1312 | ~v_1307 | ~v_1306 | ~v_1305 | ~v_1304 | v_1556;
assign x_27069 = v_13 | v_18 | v_17 | v_16 | v_15 | v_14 | v_10 | ~v_453 | ~v_709 | ~v_452 | ~v_708 | v_136 | v_135 | ~v_707 | ~v_706 | v_162 | v_161 | v_182 | ~v_233 | ~v_232 | ~v_1446 | ~v_1302 | ~v_1445 | ~v_1301 | ~v_1300 | ~v_1444 | ~v_1299 | ~v_1443 | ~v_1298 | ~v_1297 | ~v_1442 | ~v_1292 | ~v_1441 | ~v_1291 | ~v_1290 | ~v_1440 | ~v_1289 | ~v_1439 | ~v_1288 | ~v_1287 | ~v_1282 | ~v_1281 | ~v_1280 | ~v_1279 | v_1555;
assign x_27070 = v_1554 | ~v_1551;
assign x_27071 = v_1554 | ~v_1552;
assign x_27072 = v_1554 | ~v_1553;
assign x_27073 = v_103 | v_101 | v_99 | v_93 | v_102 | v_171 | v_170 | v_149 | v_148 | v_147 | v_184 | v_181 | ~v_483 | ~v_482 | ~v_481 | ~v_480 | ~v_345 | ~v_479 | ~v_478 | ~v_344 | ~v_1464 | ~v_1463 | ~v_1350 | ~v_1462 | ~v_1461 | ~v_1347 | ~v_1540 | ~v_1539 | ~v_1538 | ~v_1537 | ~v_1460 | ~v_1459 | ~v_1340 | ~v_1458 | ~v_1457 | ~v_1337 | ~v_1536 | ~v_1535 | ~v_1534 | ~v_1533 | ~v_1332 | ~v_1331 | ~v_1330 | ~v_1329 | v_1553;
assign x_27074 = v_61 | v_51 | v_60 | v_59 | v_57 | v_144 | v_180 | v_143 | v_142 | v_167 | v_166 | v_183 | ~v_468 | ~v_467 | ~v_466 | ~v_465 | ~v_330 | ~v_464 | ~v_463 | ~v_329 | ~v_1455 | ~v_1454 | ~v_1325 | ~v_1453 | ~v_1452 | ~v_1322 | ~v_1531 | ~v_1530 | ~v_1529 | ~v_1528 | ~v_1451 | ~v_1450 | ~v_1315 | ~v_1449 | ~v_1448 | ~v_1312 | ~v_1527 | ~v_1526 | ~v_1525 | ~v_1524 | ~v_1307 | ~v_1306 | ~v_1305 | ~v_1304 | v_1552;
assign x_27075 = v_18 | v_17 | v_16 | v_8 | v_14 | ~v_453 | ~v_452 | v_136 | v_135 | v_134 | v_179 | v_163 | v_162 | v_182 | ~v_451 | ~v_450 | ~v_315 | ~v_449 | ~v_448 | ~v_314 | ~v_1446 | ~v_1445 | ~v_1300 | ~v_1444 | ~v_1443 | ~v_1297 | ~v_1522 | ~v_1521 | ~v_1520 | ~v_1519 | ~v_1442 | ~v_1441 | ~v_1290 | ~v_1440 | ~v_1439 | ~v_1287 | ~v_1518 | ~v_1517 | ~v_1516 | ~v_1515 | ~v_1282 | ~v_1281 | ~v_1280 | ~v_1279 | v_1551;
assign x_27076 = v_1550 | ~v_1547;
assign x_27077 = v_1550 | ~v_1548;
assign x_27078 = v_1550 | ~v_1549;
assign x_27079 = v_103 | v_96 | v_95 | v_93 | v_102 | v_171 | v_170 | v_160 | v_150 | v_149 | v_184 | v_181 | ~v_297 | ~v_296 | ~v_345 | ~v_344 | ~v_343 | ~v_342 | ~v_341 | ~v_340 | ~v_1350 | ~v_1347 | ~v_1436 | ~v_1435 | ~v_1434 | ~v_1433 | ~v_1540 | ~v_1539 | ~v_1538 | ~v_1537 | ~v_1340 | ~v_1337 | ~v_1536 | ~v_1535 | ~v_1534 | ~v_1533 | ~v_1432 | ~v_1431 | ~v_1430 | ~v_1429 | ~v_1332 | ~v_1331 | ~v_1330 | ~v_1329 | v_1549;
assign x_27080 = v_54 | v_53 | v_61 | v_51 | v_60 | v_144 | v_180 | v_159 | v_145 | v_167 | v_166 | v_183 | ~v_264 | ~v_263 | ~v_330 | ~v_329 | ~v_328 | ~v_327 | ~v_326 | ~v_325 | ~v_1325 | ~v_1322 | ~v_1427 | ~v_1426 | ~v_1425 | ~v_1424 | ~v_1531 | ~v_1530 | ~v_1529 | ~v_1528 | ~v_1315 | ~v_1312 | ~v_1527 | ~v_1526 | ~v_1525 | ~v_1524 | ~v_1423 | ~v_1422 | ~v_1421 | ~v_1420 | ~v_1307 | ~v_1306 | ~v_1305 | ~v_1304 | v_1548;
assign x_27081 = v_18 | v_17 | v_8 | v_11 | v_10 | v_136 | v_137 | v_179 | v_163 | v_162 | v_155 | v_182 | ~v_231 | ~v_230 | ~v_315 | ~v_314 | ~v_313 | ~v_312 | ~v_311 | ~v_310 | ~v_1300 | ~v_1297 | ~v_1418 | ~v_1417 | ~v_1416 | ~v_1415 | ~v_1522 | ~v_1521 | ~v_1520 | ~v_1519 | ~v_1290 | ~v_1287 | ~v_1518 | ~v_1517 | ~v_1516 | ~v_1515 | ~v_1414 | ~v_1413 | ~v_1412 | ~v_1411 | ~v_1282 | ~v_1281 | ~v_1280 | ~v_1279 | v_1547;
assign x_27082 = v_1546 | ~v_1543;
assign x_27083 = v_1546 | ~v_1544;
assign x_27084 = v_1546 | ~v_1545;
assign x_27085 = v_103 | v_101 | v_93 | v_102 | v_171 | v_170 | v_150 | v_149 | v_148 | v_147 | v_184 | v_181 | ~v_391 | ~v_390 | ~v_387 | ~v_386 | ~v_345 | ~v_344 | ~v_385 | ~v_384 | ~v_1350 | ~v_1347 | ~v_1408 | ~v_1407 | ~v_1406 | ~v_1405 | ~v_1540 | ~v_1539 | ~v_1538 | ~v_1537 | ~v_1340 | ~v_1337 | ~v_1536 | ~v_1535 | ~v_1534 | ~v_1533 | ~v_1404 | ~v_1403 | ~v_1402 | ~v_1401 | ~v_1332 | ~v_1331 | ~v_1330 | ~v_1329 | v_1545;
assign x_27086 = v_61 | v_51 | v_60 | v_59 | v_144 | v_180 | v_145 | v_143 | v_142 | v_167 | v_166 | v_183 | ~v_376 | ~v_375 | ~v_372 | ~v_371 | ~v_330 | ~v_329 | ~v_370 | ~v_369 | ~v_1325 | ~v_1322 | ~v_1399 | ~v_1398 | ~v_1397 | ~v_1396 | ~v_1531 | ~v_1530 | ~v_1529 | ~v_1528 | ~v_1315 | ~v_1312 | ~v_1527 | ~v_1526 | ~v_1525 | ~v_1524 | ~v_1395 | ~v_1394 | ~v_1393 | ~v_1392 | ~v_1307 | ~v_1306 | ~v_1305 | ~v_1304 | v_1544;
assign x_27087 = v_18 | v_17 | v_16 | v_8 | v_136 | v_135 | v_134 | v_137 | v_179 | v_163 | v_162 | v_182 | ~v_361 | ~v_360 | ~v_357 | ~v_356 | ~v_315 | ~v_314 | ~v_355 | ~v_354 | ~v_1300 | ~v_1297 | ~v_1390 | ~v_1389 | ~v_1388 | ~v_1387 | ~v_1522 | ~v_1521 | ~v_1520 | ~v_1519 | ~v_1290 | ~v_1287 | ~v_1518 | ~v_1517 | ~v_1516 | ~v_1515 | ~v_1386 | ~v_1385 | ~v_1384 | ~v_1383 | ~v_1282 | ~v_1281 | ~v_1280 | ~v_1279 | v_1543;
assign x_27088 = v_1542 | ~v_1523;
assign x_27089 = v_1542 | ~v_1532;
assign x_27090 = v_1542 | ~v_1541;
assign x_27091 = v_101 | v_97 | v_93 | v_102 | v_172 | v_171 | v_170 | v_150 | v_148 | v_147 | v_184 | v_181 | ~v_437 | ~v_436 | ~v_435 | ~v_434 | ~v_345 | ~v_344 | ~v_433 | ~v_432 | ~v_1350 | ~v_1347 | ~v_1346 | ~v_1345 | ~v_1344 | ~v_1343 | ~v_1540 | ~v_1539 | ~v_1538 | ~v_1537 | ~v_1340 | ~v_1337 | ~v_1536 | ~v_1535 | ~v_1534 | ~v_1533 | ~v_1336 | ~v_1335 | ~v_1334 | ~v_1333 | ~v_1332 | ~v_1331 | ~v_1330 | ~v_1329 | v_1541;
assign x_27092 = v_1540 | v_178;
assign x_27093 = v_1540 | v_128;
assign x_27094 = v_1539 | v_177;
assign x_27095 = v_1539 | v_125;
assign x_27096 = v_1538 | ~v_178;
assign x_27097 = v_1538 | v_113;
assign x_27098 = v_1537 | ~v_177;
assign x_27099 = v_1537 | v_110;
assign x_27100 = v_1536 | v_158;
assign x_27101 = v_1536 | v_127;
assign x_27102 = v_1535 | v_158;
assign x_27103 = v_1535 | v_121;
assign x_27104 = v_1534 | ~v_158;
assign x_27105 = v_1534 | v_112;
assign x_27106 = v_1533 | ~v_158;
assign x_27107 = v_1533 | v_106;
assign x_27108 = v_55 | v_51 | v_60 | v_59 | v_180 | v_145 | v_143 | v_142 | v_168 | v_167 | v_166 | v_183 | ~v_422 | ~v_421 | ~v_420 | ~v_419 | ~v_330 | ~v_329 | ~v_418 | ~v_417 | ~v_1325 | ~v_1322 | ~v_1321 | ~v_1320 | ~v_1319 | ~v_1318 | ~v_1531 | ~v_1530 | ~v_1529 | ~v_1528 | ~v_1315 | ~v_1312 | ~v_1527 | ~v_1526 | ~v_1525 | ~v_1524 | ~v_1311 | ~v_1310 | ~v_1309 | ~v_1308 | ~v_1307 | ~v_1306 | ~v_1305 | ~v_1304 | v_1532;
assign x_27109 = v_1531 | v_178;
assign x_27110 = v_1531 | v_86;
assign x_27111 = v_1530 | v_177;
assign x_27112 = v_1530 | v_83;
assign x_27113 = v_1529 | ~v_178;
assign x_27114 = v_1529 | v_71;
assign x_27115 = v_1528 | ~v_177;
assign x_27116 = v_1528 | v_68;
assign x_27117 = v_1527 | v_158;
assign x_27118 = v_1527 | v_85;
assign x_27119 = v_1526 | v_158;
assign x_27120 = v_1526 | v_79;
assign x_27121 = v_1525 | ~v_158;
assign x_27122 = v_1525 | v_70;
assign x_27123 = v_1524 | ~v_158;
assign x_27124 = v_1524 | v_64;
assign x_27125 = v_17 | v_16 | v_8 | v_12 | v_135 | v_134 | v_137 | v_179 | v_164 | v_163 | v_162 | v_182 | ~v_407 | ~v_406 | ~v_405 | ~v_404 | ~v_315 | ~v_314 | ~v_403 | ~v_402 | ~v_1300 | ~v_1297 | ~v_1296 | ~v_1295 | ~v_1294 | ~v_1293 | ~v_1522 | ~v_1521 | ~v_1520 | ~v_1519 | ~v_1290 | ~v_1287 | ~v_1518 | ~v_1517 | ~v_1516 | ~v_1515 | ~v_1286 | ~v_1285 | ~v_1284 | ~v_1283 | ~v_1282 | ~v_1281 | ~v_1280 | ~v_1279 | v_1523;
assign x_27126 = v_1522 | v_178;
assign x_27127 = v_1522 | v_44;
assign x_27128 = v_1521 | v_177;
assign x_27129 = v_1521 | v_41;
assign x_27130 = v_1520 | ~v_178;
assign x_27131 = v_1520 | v_29;
assign x_27132 = v_1519 | ~v_177;
assign x_27133 = v_1519 | v_26;
assign x_27134 = v_1518 | v_158;
assign x_27135 = v_1518 | v_43;
assign x_27136 = v_1517 | v_158;
assign x_27137 = v_1517 | v_37;
assign x_27138 = v_1516 | ~v_158;
assign x_27139 = v_1516 | v_28;
assign x_27140 = v_1515 | ~v_158;
assign x_27141 = v_1515 | v_22;
assign x_27142 = v_1514 | ~v_1511;
assign x_27143 = v_1514 | ~v_1512;
assign x_27144 = v_1514 | ~v_1513;
assign x_27145 = v_98 | v_103 | v_96 | v_100 | v_102 | v_170 | v_169 | v_160 | v_150 | v_149 | v_147 | v_184 | ~v_299 | ~v_298 | ~v_297 | ~v_296 | ~v_295 | ~v_294 | ~v_293 | ~v_292 | ~v_1352 | ~v_1351 | ~v_1350 | ~v_1349 | ~v_1348 | ~v_1347 | ~v_1436 | ~v_1435 | ~v_1434 | ~v_1433 | ~v_1342 | ~v_1341 | ~v_1340 | ~v_1339 | ~v_1338 | ~v_1337 | ~v_1432 | ~v_1431 | ~v_1430 | ~v_1429 | ~v_1332 | ~v_1331 | ~v_1330 | ~v_1329 | v_1513;
assign x_27146 = v_54 | v_56 | v_61 | v_60 | v_58 | v_144 | v_159 | v_145 | v_142 | v_166 | v_165 | v_183 | ~v_266 | ~v_265 | ~v_264 | ~v_263 | ~v_262 | ~v_261 | ~v_260 | ~v_259 | ~v_1327 | ~v_1326 | ~v_1325 | ~v_1324 | ~v_1323 | ~v_1322 | ~v_1427 | ~v_1426 | ~v_1425 | ~v_1424 | ~v_1317 | ~v_1316 | ~v_1315 | ~v_1314 | ~v_1313 | ~v_1312 | ~v_1423 | ~v_1422 | ~v_1421 | ~v_1420 | ~v_1307 | ~v_1306 | ~v_1305 | ~v_1304 | v_1512;
assign x_27147 = v_13 | v_18 | v_17 | v_15 | v_11 | v_136 | v_134 | v_137 | v_162 | v_161 | v_155 | v_182 | ~v_233 | ~v_232 | ~v_231 | ~v_230 | ~v_229 | ~v_228 | ~v_227 | ~v_226 | ~v_1302 | ~v_1301 | ~v_1300 | ~v_1299 | ~v_1298 | ~v_1297 | ~v_1418 | ~v_1417 | ~v_1416 | ~v_1415 | ~v_1292 | ~v_1291 | ~v_1290 | ~v_1289 | ~v_1288 | ~v_1287 | ~v_1414 | ~v_1413 | ~v_1412 | ~v_1411 | ~v_1282 | ~v_1281 | ~v_1280 | ~v_1279 | v_1511;
assign x_27148 = v_1510 | ~v_1507;
assign x_27149 = v_1510 | ~v_1508;
assign x_27150 = v_1510 | ~v_1509;
assign x_27151 = v_101 | v_100 | v_99 | v_102 | v_172 | v_171 | v_170 | v_169 | v_149 | v_148 | v_147 | v_184 | ~v_483 | ~v_482 | ~v_593 | ~v_592 | ~v_545 | ~v_591 | ~v_590 | ~v_544 | ~v_1464 | ~v_1463 | ~v_1350 | ~v_1462 | ~v_1461 | ~v_1347 | ~v_1496 | ~v_1495 | ~v_1494 | ~v_1493 | ~v_1460 | ~v_1459 | ~v_1340 | ~v_1458 | ~v_1457 | ~v_1337 | ~v_1492 | ~v_1491 | ~v_1490 | ~v_1489 | ~v_1332 | ~v_1331 | ~v_1330 | ~v_1329 | v_1509;
assign x_27152 = v_60 | v_59 | v_58 | v_57 | v_144 | v_143 | v_142 | v_168 | v_167 | v_166 | v_165 | v_183 | ~v_468 | ~v_467 | ~v_588 | ~v_587 | ~v_530 | ~v_586 | ~v_585 | ~v_529 | ~v_1455 | ~v_1454 | ~v_1325 | ~v_1453 | ~v_1452 | ~v_1322 | ~v_1487 | ~v_1486 | ~v_1485 | ~v_1484 | ~v_1451 | ~v_1450 | ~v_1315 | ~v_1449 | ~v_1448 | ~v_1312 | ~v_1483 | ~v_1482 | ~v_1481 | ~v_1480 | ~v_1307 | ~v_1306 | ~v_1305 | ~v_1304 | v_1508;
assign x_27153 = v_17 | v_16 | v_15 | v_14 | ~v_453 | ~v_452 | v_136 | v_135 | v_134 | v_164 | v_163 | v_162 | v_161 | v_182 | ~v_583 | ~v_582 | ~v_515 | ~v_581 | ~v_580 | ~v_514 | ~v_1446 | ~v_1445 | ~v_1300 | ~v_1444 | ~v_1443 | ~v_1297 | ~v_1478 | ~v_1477 | ~v_1476 | ~v_1475 | ~v_1442 | ~v_1441 | ~v_1290 | ~v_1440 | ~v_1439 | ~v_1287 | ~v_1474 | ~v_1473 | ~v_1472 | ~v_1471 | ~v_1282 | ~v_1281 | ~v_1280 | ~v_1279 | v_1507;
assign x_27154 = v_1506 | ~v_1503;
assign x_27155 = v_1506 | ~v_1504;
assign x_27156 = v_1506 | ~v_1505;
assign x_27157 = v_103 | v_96 | v_100 | v_102 | v_171 | v_170 | v_169 | v_160 | v_150 | v_149 | v_147 | v_184 | ~v_545 | ~v_544 | ~v_543 | ~v_542 | ~v_541 | ~v_540 | ~v_297 | ~v_296 | ~v_1350 | ~v_1347 | ~v_1436 | ~v_1435 | ~v_1434 | ~v_1433 | ~v_1496 | ~v_1495 | ~v_1494 | ~v_1493 | ~v_1340 | ~v_1337 | ~v_1432 | ~v_1431 | ~v_1430 | ~v_1429 | ~v_1492 | ~v_1491 | ~v_1490 | ~v_1489 | ~v_1332 | ~v_1331 | ~v_1330 | ~v_1329 | v_1505;
assign x_27158 = v_54 | v_61 | v_60 | v_58 | v_144 | v_159 | v_145 | v_142 | v_167 | v_166 | v_165 | v_183 | ~v_530 | ~v_529 | ~v_528 | ~v_527 | ~v_526 | ~v_525 | ~v_264 | ~v_263 | ~v_1325 | ~v_1322 | ~v_1427 | ~v_1426 | ~v_1425 | ~v_1424 | ~v_1487 | ~v_1486 | ~v_1485 | ~v_1484 | ~v_1315 | ~v_1312 | ~v_1423 | ~v_1422 | ~v_1421 | ~v_1420 | ~v_1483 | ~v_1482 | ~v_1481 | ~v_1480 | ~v_1307 | ~v_1306 | ~v_1305 | ~v_1304 | v_1504;
assign x_27159 = v_18 | v_17 | v_15 | v_11 | v_136 | v_134 | v_137 | v_163 | v_162 | v_161 | v_155 | v_182 | ~v_515 | ~v_514 | ~v_513 | ~v_512 | ~v_511 | ~v_510 | ~v_231 | ~v_230 | ~v_1300 | ~v_1297 | ~v_1418 | ~v_1417 | ~v_1416 | ~v_1415 | ~v_1478 | ~v_1477 | ~v_1476 | ~v_1475 | ~v_1290 | ~v_1287 | ~v_1414 | ~v_1413 | ~v_1412 | ~v_1411 | ~v_1474 | ~v_1473 | ~v_1472 | ~v_1471 | ~v_1282 | ~v_1281 | ~v_1280 | ~v_1279 | v_1503;
assign x_27160 = v_1502 | ~v_1499;
assign x_27161 = v_1502 | ~v_1500;
assign x_27162 = v_1502 | ~v_1501;
assign x_27163 = v_103 | v_101 | v_100 | v_95 | v_102 | v_171 | v_170 | v_169 | v_150 | v_149 | v_148 | v_184 | ~v_545 | ~v_544 | ~v_561 | ~v_560 | ~v_559 | ~v_558 | ~v_387 | ~v_386 | ~v_1350 | ~v_1347 | ~v_1408 | ~v_1407 | ~v_1406 | ~v_1405 | ~v_1496 | ~v_1495 | ~v_1494 | ~v_1493 | ~v_1340 | ~v_1337 | ~v_1404 | ~v_1403 | ~v_1402 | ~v_1401 | ~v_1492 | ~v_1491 | ~v_1490 | ~v_1489 | ~v_1332 | ~v_1331 | ~v_1330 | ~v_1329 | v_1501;
assign x_27164 = v_53 | v_61 | v_60 | v_59 | v_58 | v_144 | v_145 | v_143 | v_167 | v_166 | v_165 | v_183 | ~v_530 | ~v_529 | ~v_556 | ~v_555 | ~v_554 | ~v_553 | ~v_372 | ~v_371 | ~v_1325 | ~v_1322 | ~v_1399 | ~v_1398 | ~v_1397 | ~v_1396 | ~v_1487 | ~v_1486 | ~v_1485 | ~v_1484 | ~v_1315 | ~v_1312 | ~v_1395 | ~v_1394 | ~v_1393 | ~v_1392 | ~v_1483 | ~v_1482 | ~v_1481 | ~v_1480 | ~v_1307 | ~v_1306 | ~v_1305 | ~v_1304 | v_1500;
assign x_27165 = v_18 | v_17 | v_16 | v_15 | v_10 | v_136 | v_135 | v_137 | v_163 | v_162 | v_161 | v_182 | ~v_515 | ~v_514 | ~v_551 | ~v_550 | ~v_549 | ~v_548 | ~v_357 | ~v_356 | ~v_1300 | ~v_1297 | ~v_1390 | ~v_1389 | ~v_1388 | ~v_1387 | ~v_1478 | ~v_1477 | ~v_1476 | ~v_1475 | ~v_1290 | ~v_1287 | ~v_1386 | ~v_1385 | ~v_1384 | ~v_1383 | ~v_1474 | ~v_1473 | ~v_1472 | ~v_1471 | ~v_1282 | ~v_1281 | ~v_1280 | ~v_1279 | v_1499;
assign x_27166 = v_1498 | ~v_1479;
assign x_27167 = v_1498 | ~v_1488;
assign x_27168 = v_1498 | ~v_1497;
assign x_27169 = v_103 | v_101 | v_97 | v_100 | v_151 | v_171 | v_170 | v_169 | v_150 | v_148 | v_147 | v_184 | ~v_577 | ~v_576 | ~v_545 | ~v_544 | ~v_575 | ~v_574 | ~v_435 | ~v_434 | ~v_1350 | ~v_1347 | ~v_1346 | ~v_1345 | ~v_1344 | ~v_1343 | ~v_1496 | ~v_1495 | ~v_1494 | ~v_1493 | ~v_1340 | ~v_1337 | ~v_1336 | ~v_1335 | ~v_1334 | ~v_1333 | ~v_1492 | ~v_1491 | ~v_1490 | ~v_1489 | ~v_1332 | ~v_1331 | ~v_1330 | ~v_1329 | v_1497;
assign x_27170 = v_1496 | v_173;
assign x_27171 = v_1496 | v_128;
assign x_27172 = v_1495 | v_174;
assign x_27173 = v_1495 | v_125;
assign x_27174 = v_1494 | ~v_173;
assign x_27175 = v_1494 | v_113;
assign x_27176 = v_1493 | ~v_174;
assign x_27177 = v_1493 | v_110;
assign x_27178 = v_1492 | v_175;
assign x_27179 = v_1492 | v_127;
assign x_27180 = v_1491 | v_176;
assign x_27181 = v_1491 | v_121;
assign x_27182 = v_1490 | ~v_175;
assign x_27183 = v_1490 | v_112;
assign x_27184 = v_1489 | ~v_176;
assign x_27185 = v_1489 | v_106;
assign x_27186 = v_55 | v_61 | v_59 | v_58 | v_145 | v_143 | v_142 | v_167 | v_166 | v_165 | v_146 | v_183 | ~v_572 | ~v_571 | ~v_530 | ~v_529 | ~v_570 | ~v_569 | ~v_420 | ~v_419 | ~v_1325 | ~v_1322 | ~v_1321 | ~v_1320 | ~v_1319 | ~v_1318 | ~v_1487 | ~v_1486 | ~v_1485 | ~v_1484 | ~v_1315 | ~v_1312 | ~v_1311 | ~v_1310 | ~v_1309 | ~v_1308 | ~v_1483 | ~v_1482 | ~v_1481 | ~v_1480 | ~v_1307 | ~v_1306 | ~v_1305 | ~v_1304 | v_1488;
assign x_27187 = v_1487 | v_173;
assign x_27188 = v_1487 | v_86;
assign x_27189 = v_1486 | v_174;
assign x_27190 = v_1486 | v_83;
assign x_27191 = v_1485 | ~v_173;
assign x_27192 = v_1485 | v_71;
assign x_27193 = v_1484 | ~v_174;
assign x_27194 = v_1484 | v_68;
assign x_27195 = v_1483 | v_175;
assign x_27196 = v_1483 | v_85;
assign x_27197 = v_1482 | v_176;
assign x_27198 = v_1482 | v_79;
assign x_27199 = v_1481 | ~v_175;
assign x_27200 = v_1481 | v_70;
assign x_27201 = v_1480 | ~v_176;
assign x_27202 = v_1480 | v_64;
assign x_27203 = v_18 | v_16 | v_15 | v_12 | v_135 | v_134 | v_137 | v_138 | v_163 | v_162 | v_161 | v_182 | ~v_567 | ~v_566 | ~v_515 | ~v_514 | ~v_565 | ~v_564 | ~v_405 | ~v_404 | ~v_1300 | ~v_1297 | ~v_1296 | ~v_1295 | ~v_1294 | ~v_1293 | ~v_1478 | ~v_1477 | ~v_1476 | ~v_1475 | ~v_1290 | ~v_1287 | ~v_1286 | ~v_1285 | ~v_1284 | ~v_1283 | ~v_1474 | ~v_1473 | ~v_1472 | ~v_1471 | ~v_1282 | ~v_1281 | ~v_1280 | ~v_1279 | v_1479;
assign x_27204 = v_1478 | v_173;
assign x_27205 = v_1478 | v_44;
assign x_27206 = v_1477 | v_174;
assign x_27207 = v_1477 | v_41;
assign x_27208 = v_1476 | ~v_173;
assign x_27209 = v_1476 | v_29;
assign x_27210 = v_1475 | ~v_174;
assign x_27211 = v_1475 | v_26;
assign x_27212 = v_1474 | v_175;
assign x_27213 = v_1474 | v_43;
assign x_27214 = v_1473 | v_176;
assign x_27215 = v_1473 | v_37;
assign x_27216 = v_1472 | ~v_175;
assign x_27217 = v_1472 | v_28;
assign x_27218 = v_1471 | ~v_176;
assign x_27219 = v_1471 | v_22;
assign x_27220 = v_1470 | ~v_1467;
assign x_27221 = v_1470 | ~v_1468;
assign x_27222 = v_1470 | ~v_1469;
assign x_27223 = v_98 | v_103 | v_101 | v_100 | v_151 | v_170 | v_169 | v_150 | v_149 | v_148 | v_147 | v_184 | ~v_299 | ~v_298 | ~v_387 | ~v_386 | ~v_499 | ~v_498 | ~v_497 | ~v_496 | ~v_1352 | ~v_1351 | ~v_1350 | ~v_1349 | ~v_1348 | ~v_1347 | ~v_1408 | ~v_1407 | ~v_1406 | ~v_1405 | ~v_1342 | ~v_1341 | ~v_1340 | ~v_1339 | ~v_1338 | ~v_1337 | ~v_1404 | ~v_1403 | ~v_1402 | ~v_1401 | ~v_1332 | ~v_1331 | ~v_1330 | ~v_1329 | v_1469;
assign x_27224 = v_56 | v_61 | v_59 | v_58 | v_144 | v_145 | v_143 | v_142 | v_166 | v_165 | v_146 | v_183 | ~v_266 | ~v_265 | ~v_372 | ~v_371 | ~v_494 | ~v_493 | ~v_492 | ~v_491 | ~v_1327 | ~v_1326 | ~v_1325 | ~v_1324 | ~v_1323 | ~v_1322 | ~v_1399 | ~v_1398 | ~v_1397 | ~v_1396 | ~v_1317 | ~v_1316 | ~v_1315 | ~v_1314 | ~v_1313 | ~v_1312 | ~v_1395 | ~v_1394 | ~v_1393 | ~v_1392 | ~v_1307 | ~v_1306 | ~v_1305 | ~v_1304 | v_1468;
assign x_27225 = v_13 | v_18 | v_16 | v_15 | v_136 | v_135 | v_134 | v_137 | v_138 | v_162 | v_161 | v_182 | ~v_233 | ~v_232 | ~v_357 | ~v_356 | ~v_489 | ~v_488 | ~v_487 | ~v_486 | ~v_1302 | ~v_1301 | ~v_1300 | ~v_1299 | ~v_1298 | ~v_1297 | ~v_1390 | ~v_1389 | ~v_1388 | ~v_1387 | ~v_1292 | ~v_1291 | ~v_1290 | ~v_1289 | ~v_1288 | ~v_1287 | ~v_1386 | ~v_1385 | ~v_1384 | ~v_1383 | ~v_1282 | ~v_1281 | ~v_1280 | ~v_1279 | v_1467;
assign x_27226 = v_1466 | ~v_1447;
assign x_27227 = v_1466 | ~v_1456;
assign x_27228 = v_1466 | ~v_1465;
assign x_27229 = v_103 | v_101 | v_100 | v_94 | v_99 | v_102 | v_171 | v_169 | v_149 | v_148 | v_147 | v_184 | ~v_703 | ~v_702 | ~v_483 | ~v_482 | ~v_701 | ~v_653 | ~v_700 | ~v_652 | ~v_1464 | ~v_1463 | ~v_1350 | ~v_1462 | ~v_1461 | ~v_1347 | ~v_1380 | ~v_1379 | ~v_1378 | ~v_1377 | ~v_1460 | ~v_1459 | ~v_1340 | ~v_1458 | ~v_1457 | ~v_1337 | ~v_1376 | ~v_1375 | ~v_1374 | ~v_1373 | ~v_1332 | ~v_1331 | ~v_1330 | ~v_1329 | v_1465;
assign x_27230 = v_1464 | v_152;
assign x_27231 = v_1464 | v_131;
assign x_27232 = v_1463 | v_153;
assign x_27233 = v_1463 | v_126;
assign x_27234 = v_1462 | ~v_152;
assign x_27235 = v_1462 | v_116;
assign x_27236 = v_1461 | ~v_153;
assign x_27237 = v_1461 | v_111;
assign x_27238 = v_1460 | v_156;
assign x_27239 = v_1460 | v_130;
assign x_27240 = v_1459 | v_157;
assign x_27241 = v_1459 | v_122;
assign x_27242 = v_1458 | ~v_156;
assign x_27243 = v_1458 | v_115;
assign x_27244 = v_1457 | ~v_157;
assign x_27245 = v_1457 | v_107;
assign x_27246 = v_61 | v_52 | v_60 | v_59 | v_58 | v_57 | v_144 | v_143 | v_142 | v_167 | v_165 | v_183 | ~v_698 | ~v_697 | ~v_468 | ~v_467 | ~v_696 | ~v_638 | ~v_695 | ~v_637 | ~v_1455 | ~v_1454 | ~v_1325 | ~v_1453 | ~v_1452 | ~v_1322 | ~v_1371 | ~v_1370 | ~v_1369 | ~v_1368 | ~v_1451 | ~v_1450 | ~v_1315 | ~v_1449 | ~v_1448 | ~v_1312 | ~v_1367 | ~v_1366 | ~v_1365 | ~v_1364 | ~v_1307 | ~v_1306 | ~v_1305 | ~v_1304 | v_1456;
assign x_27247 = v_1455 | v_152;
assign x_27248 = v_1455 | v_89;
assign x_27249 = v_1454 | v_153;
assign x_27250 = v_1454 | v_84;
assign x_27251 = v_1453 | ~v_152;
assign x_27252 = v_1453 | v_74;
assign x_27253 = v_1452 | ~v_153;
assign x_27254 = v_1452 | v_69;
assign x_27255 = v_1451 | v_156;
assign x_27256 = v_1451 | v_88;
assign x_27257 = v_1450 | v_157;
assign x_27258 = v_1450 | v_80;
assign x_27259 = v_1449 | ~v_156;
assign x_27260 = v_1449 | v_73;
assign x_27261 = v_1448 | ~v_157;
assign x_27262 = v_1448 | v_65;
assign x_27263 = v_9 | v_18 | v_17 | v_16 | v_15 | v_14 | ~v_453 | ~v_452 | v_136 | v_135 | v_134 | v_163 | v_161 | v_182 | ~v_693 | ~v_692 | ~v_691 | ~v_623 | ~v_690 | ~v_622 | ~v_1446 | ~v_1445 | ~v_1300 | ~v_1444 | ~v_1443 | ~v_1297 | ~v_1362 | ~v_1361 | ~v_1360 | ~v_1359 | ~v_1442 | ~v_1441 | ~v_1290 | ~v_1440 | ~v_1439 | ~v_1287 | ~v_1358 | ~v_1357 | ~v_1356 | ~v_1355 | ~v_1282 | ~v_1281 | ~v_1280 | ~v_1279 | v_1447;
assign x_27264 = v_1446 | v_152;
assign x_27265 = v_1446 | v_47;
assign x_27266 = v_1445 | v_153;
assign x_27267 = v_1445 | v_42;
assign x_27268 = v_1444 | ~v_152;
assign x_27269 = v_1444 | v_32;
assign x_27270 = v_1443 | ~v_153;
assign x_27271 = v_1443 | v_27;
assign x_27272 = v_1442 | v_156;
assign x_27273 = v_1442 | v_46;
assign x_27274 = v_1441 | v_157;
assign x_27275 = v_1441 | v_38;
assign x_27276 = v_1440 | ~v_156;
assign x_27277 = v_1440 | v_31;
assign x_27278 = v_1439 | ~v_157;
assign x_27279 = v_1439 | v_23;
assign x_27280 = v_1438 | ~v_1419;
assign x_27281 = v_1438 | ~v_1428;
assign x_27282 = v_1438 | ~v_1437;
assign x_27283 = v_103 | v_96 | v_100 | v_94 | v_151 | v_171 | v_169 | v_160 | v_150 | v_149 | v_147 | v_184 | ~v_655 | ~v_654 | ~v_297 | ~v_296 | ~v_653 | ~v_652 | ~v_651 | ~v_650 | ~v_1350 | ~v_1347 | ~v_1380 | ~v_1379 | ~v_1378 | ~v_1377 | ~v_1436 | ~v_1435 | ~v_1434 | ~v_1433 | ~v_1340 | ~v_1337 | ~v_1432 | ~v_1431 | ~v_1430 | ~v_1429 | ~v_1376 | ~v_1375 | ~v_1374 | ~v_1373 | ~v_1332 | ~v_1331 | ~v_1330 | ~v_1329 | v_1437;
assign x_27284 = v_1436 | v_178;
assign x_27285 = v_1436 | v_131;
assign x_27286 = v_1435 | v_177;
assign x_27287 = v_1435 | v_126;
assign x_27288 = v_1434 | ~v_178;
assign x_27289 = v_1434 | v_116;
assign x_27290 = v_1433 | ~v_177;
assign x_27291 = v_1433 | v_111;
assign x_27292 = v_1432 | v_158;
assign x_27293 = v_1432 | v_130;
assign x_27294 = v_1431 | v_158;
assign x_27295 = v_1431 | v_122;
assign x_27296 = v_1430 | ~v_158;
assign x_27297 = v_1430 | v_115;
assign x_27298 = v_1429 | ~v_158;
assign x_27299 = v_1429 | v_107;
assign x_27300 = v_54 | v_61 | v_52 | v_58 | v_144 | v_159 | v_145 | v_142 | v_167 | v_165 | v_146 | v_183 | ~v_640 | ~v_639 | ~v_264 | ~v_263 | ~v_638 | ~v_637 | ~v_636 | ~v_635 | ~v_1325 | ~v_1322 | ~v_1371 | ~v_1370 | ~v_1369 | ~v_1368 | ~v_1427 | ~v_1426 | ~v_1425 | ~v_1424 | ~v_1315 | ~v_1312 | ~v_1423 | ~v_1422 | ~v_1421 | ~v_1420 | ~v_1367 | ~v_1366 | ~v_1365 | ~v_1364 | ~v_1307 | ~v_1306 | ~v_1305 | ~v_1304 | v_1428;
assign x_27301 = v_1427 | v_178;
assign x_27302 = v_1427 | v_89;
assign x_27303 = v_1426 | v_177;
assign x_27304 = v_1426 | v_84;
assign x_27305 = v_1425 | ~v_178;
assign x_27306 = v_1425 | v_74;
assign x_27307 = v_1424 | ~v_177;
assign x_27308 = v_1424 | v_69;
assign x_27309 = v_1423 | v_158;
assign x_27310 = v_1423 | v_88;
assign x_27311 = v_1422 | v_158;
assign x_27312 = v_1422 | v_80;
assign x_27313 = v_1421 | ~v_158;
assign x_27314 = v_1421 | v_73;
assign x_27315 = v_1420 | ~v_158;
assign x_27316 = v_1420 | v_65;
assign x_27317 = v_9 | v_18 | v_15 | v_11 | v_136 | v_134 | v_137 | v_138 | v_163 | v_161 | v_155 | v_182 | ~v_625 | ~v_624 | ~v_231 | ~v_230 | ~v_623 | ~v_622 | ~v_621 | ~v_620 | ~v_1300 | ~v_1297 | ~v_1362 | ~v_1361 | ~v_1360 | ~v_1359 | ~v_1418 | ~v_1417 | ~v_1416 | ~v_1415 | ~v_1290 | ~v_1287 | ~v_1414 | ~v_1413 | ~v_1412 | ~v_1411 | ~v_1358 | ~v_1357 | ~v_1356 | ~v_1355 | ~v_1282 | ~v_1281 | ~v_1280 | ~v_1279 | v_1419;
assign x_27318 = v_1418 | v_178;
assign x_27319 = v_1418 | v_47;
assign x_27320 = v_1417 | v_177;
assign x_27321 = v_1417 | v_42;
assign x_27322 = v_1416 | ~v_178;
assign x_27323 = v_1416 | v_32;
assign x_27324 = v_1415 | ~v_177;
assign x_27325 = v_1415 | v_27;
assign x_27326 = v_1414 | v_158;
assign x_27327 = v_1414 | v_46;
assign x_27328 = v_1413 | v_158;
assign x_27329 = v_1413 | v_38;
assign x_27330 = v_1412 | ~v_158;
assign x_27331 = v_1412 | v_31;
assign x_27332 = v_1411 | ~v_158;
assign x_27333 = v_1411 | v_23;
assign x_27334 = v_1410 | ~v_1391;
assign x_27335 = v_1410 | ~v_1400;
assign x_27336 = v_1410 | ~v_1409;
assign x_27337 = v_101 | v_100 | v_94 | v_102 | v_172 | v_171 | v_169 | v_150 | v_149 | v_148 | v_147 | v_184 | ~v_671 | ~v_670 | ~v_387 | ~v_386 | ~v_653 | ~v_652 | ~v_669 | ~v_668 | ~v_1350 | ~v_1347 | ~v_1380 | ~v_1379 | ~v_1378 | ~v_1377 | ~v_1408 | ~v_1407 | ~v_1406 | ~v_1405 | ~v_1340 | ~v_1337 | ~v_1404 | ~v_1403 | ~v_1402 | ~v_1401 | ~v_1376 | ~v_1375 | ~v_1374 | ~v_1373 | ~v_1332 | ~v_1331 | ~v_1330 | ~v_1329 | v_1409;
assign x_27338 = v_1408 | v_173;
assign x_27339 = v_1408 | v_131;
assign x_27340 = v_1407 | v_174;
assign x_27341 = v_1407 | v_126;
assign x_27342 = v_1406 | ~v_173;
assign x_27343 = v_1406 | v_116;
assign x_27344 = v_1405 | ~v_174;
assign x_27345 = v_1405 | v_111;
assign x_27346 = v_1404 | v_175;
assign x_27347 = v_1404 | v_130;
assign x_27348 = v_1403 | v_176;
assign x_27349 = v_1403 | v_122;
assign x_27350 = v_1402 | ~v_175;
assign x_27351 = v_1402 | v_115;
assign x_27352 = v_1401 | ~v_176;
assign x_27353 = v_1401 | v_107;
assign x_27354 = v_52 | v_60 | v_59 | v_58 | v_144 | v_145 | v_143 | v_142 | v_168 | v_167 | v_165 | v_183 | ~v_666 | ~v_665 | ~v_372 | ~v_371 | ~v_638 | ~v_637 | ~v_664 | ~v_663 | ~v_1325 | ~v_1322 | ~v_1371 | ~v_1370 | ~v_1369 | ~v_1368 | ~v_1399 | ~v_1398 | ~v_1397 | ~v_1396 | ~v_1315 | ~v_1312 | ~v_1395 | ~v_1394 | ~v_1393 | ~v_1392 | ~v_1367 | ~v_1366 | ~v_1365 | ~v_1364 | ~v_1307 | ~v_1306 | ~v_1305 | ~v_1304 | v_1400;
assign x_27355 = v_1399 | v_173;
assign x_27356 = v_1399 | v_89;
assign x_27357 = v_1398 | v_174;
assign x_27358 = v_1398 | v_84;
assign x_27359 = v_1397 | ~v_173;
assign x_27360 = v_1397 | v_74;
assign x_27361 = v_1396 | ~v_174;
assign x_27362 = v_1396 | v_69;
assign x_27363 = v_1395 | v_175;
assign x_27364 = v_1395 | v_88;
assign x_27365 = v_1394 | v_176;
assign x_27366 = v_1394 | v_80;
assign x_27367 = v_1393 | ~v_175;
assign x_27368 = v_1393 | v_73;
assign x_27369 = v_1392 | ~v_176;
assign x_27370 = v_1392 | v_65;
assign x_27371 = v_9 | v_17 | v_16 | v_15 | v_136 | v_135 | v_134 | v_137 | v_164 | v_163 | v_161 | v_182 | ~v_661 | ~v_660 | ~v_357 | ~v_356 | ~v_623 | ~v_622 | ~v_659 | ~v_658 | ~v_1300 | ~v_1297 | ~v_1362 | ~v_1361 | ~v_1360 | ~v_1359 | ~v_1390 | ~v_1389 | ~v_1388 | ~v_1387 | ~v_1290 | ~v_1287 | ~v_1386 | ~v_1385 | ~v_1384 | ~v_1383 | ~v_1358 | ~v_1357 | ~v_1356 | ~v_1355 | ~v_1282 | ~v_1281 | ~v_1280 | ~v_1279 | v_1391;
assign x_27372 = v_1390 | v_173;
assign x_27373 = v_1390 | v_47;
assign x_27374 = v_1389 | v_174;
assign x_27375 = v_1389 | v_42;
assign x_27376 = v_1388 | ~v_173;
assign x_27377 = v_1388 | v_32;
assign x_27378 = v_1387 | ~v_174;
assign x_27379 = v_1387 | v_27;
assign x_27380 = v_1386 | v_175;
assign x_27381 = v_1386 | v_46;
assign x_27382 = v_1385 | v_176;
assign x_27383 = v_1385 | v_38;
assign x_27384 = v_1384 | ~v_175;
assign x_27385 = v_1384 | v_31;
assign x_27386 = v_1383 | ~v_176;
assign x_27387 = v_1383 | v_23;
assign x_27388 = v_1382 | ~v_1363;
assign x_27389 = v_1382 | ~v_1372;
assign x_27390 = v_1382 | ~v_1381;
assign x_27391 = v_103 | v_101 | v_97 | v_100 | v_95 | v_94 | v_102 | v_171 | v_169 | v_150 | v_148 | v_184 | ~v_435 | ~v_434 | ~v_653 | ~v_652 | ~v_687 | ~v_686 | ~v_685 | ~v_684 | ~v_1350 | ~v_1347 | ~v_1380 | ~v_1379 | ~v_1378 | ~v_1377 | ~v_1346 | ~v_1345 | ~v_1344 | ~v_1343 | ~v_1340 | ~v_1337 | ~v_1336 | ~v_1335 | ~v_1334 | ~v_1333 | ~v_1376 | ~v_1375 | ~v_1374 | ~v_1373 | ~v_1332 | ~v_1331 | ~v_1330 | ~v_1329 | v_1381;
assign x_27392 = v_1380 | v_154;
assign x_27393 = v_1380 | v_128;
assign x_27394 = v_1379 | v_154;
assign x_27395 = v_1379 | v_125;
assign x_27396 = v_1378 | ~v_154;
assign x_27397 = v_1378 | v_113;
assign x_27398 = v_1377 | ~v_154;
assign x_27399 = v_1377 | v_110;
assign x_27400 = v_1376 | v_177;
assign x_27401 = v_1376 | v_127;
assign x_27402 = v_1375 | v_178;
assign x_27403 = v_1375 | v_121;
assign x_27404 = v_1374 | ~v_177;
assign x_27405 = v_1374 | v_112;
assign x_27406 = v_1373 | ~v_178;
assign x_27407 = v_1373 | v_106;
assign x_27408 = v_53 | v_55 | v_61 | v_52 | v_60 | v_59 | v_58 | v_145 | v_143 | v_167 | v_165 | v_183 | ~v_420 | ~v_419 | ~v_638 | ~v_637 | ~v_682 | ~v_681 | ~v_680 | ~v_679 | ~v_1325 | ~v_1322 | ~v_1371 | ~v_1370 | ~v_1369 | ~v_1368 | ~v_1321 | ~v_1320 | ~v_1319 | ~v_1318 | ~v_1315 | ~v_1312 | ~v_1311 | ~v_1310 | ~v_1309 | ~v_1308 | ~v_1367 | ~v_1366 | ~v_1365 | ~v_1364 | ~v_1307 | ~v_1306 | ~v_1305 | ~v_1304 | v_1372;
assign x_27409 = v_1371 | v_154;
assign x_27410 = v_1371 | v_86;
assign x_27411 = v_1370 | v_154;
assign x_27412 = v_1370 | v_83;
assign x_27413 = v_1369 | ~v_154;
assign x_27414 = v_1369 | v_71;
assign x_27415 = v_1368 | ~v_154;
assign x_27416 = v_1368 | v_68;
assign x_27417 = v_1367 | v_177;
assign x_27418 = v_1367 | v_85;
assign x_27419 = v_1366 | v_178;
assign x_27420 = v_1366 | v_79;
assign x_27421 = v_1365 | ~v_177;
assign x_27422 = v_1365 | v_70;
assign x_27423 = v_1364 | ~v_178;
assign x_27424 = v_1364 | v_64;
assign x_27425 = v_9 | v_18 | v_17 | v_16 | v_15 | v_12 | v_10 | v_135 | v_137 | v_163 | v_161 | v_182 | ~v_405 | ~v_404 | ~v_623 | ~v_622 | ~v_677 | ~v_676 | ~v_675 | ~v_674 | ~v_1300 | ~v_1297 | ~v_1362 | ~v_1361 | ~v_1360 | ~v_1359 | ~v_1296 | ~v_1295 | ~v_1294 | ~v_1293 | ~v_1290 | ~v_1287 | ~v_1286 | ~v_1285 | ~v_1284 | ~v_1283 | ~v_1358 | ~v_1357 | ~v_1356 | ~v_1355 | ~v_1282 | ~v_1281 | ~v_1280 | ~v_1279 | v_1363;
assign x_27426 = v_1362 | v_154;
assign x_27427 = v_1362 | v_44;
assign x_27428 = v_1361 | v_154;
assign x_27429 = v_1361 | v_41;
assign x_27430 = v_1360 | ~v_154;
assign x_27431 = v_1360 | v_29;
assign x_27432 = v_1359 | ~v_154;
assign x_27433 = v_1359 | v_26;
assign x_27434 = v_1358 | v_177;
assign x_27435 = v_1358 | v_43;
assign x_27436 = v_1357 | v_178;
assign x_27437 = v_1357 | v_37;
assign x_27438 = v_1356 | ~v_177;
assign x_27439 = v_1356 | v_28;
assign x_27440 = v_1355 | ~v_178;
assign x_27441 = v_1355 | v_22;
assign x_27442 = v_1354 | ~v_1303;
assign x_27443 = v_1354 | ~v_1328;
assign x_27444 = v_1354 | ~v_1353;
assign x_27445 = v_98 | v_103 | v_101 | v_97 | v_100 | v_102 | v_170 | v_169 | v_150 | v_148 | v_147 | v_184 | ~v_609 | ~v_608 | ~v_299 | ~v_298 | ~v_435 | ~v_434 | ~v_607 | ~v_606 | ~v_1352 | ~v_1351 | ~v_1350 | ~v_1349 | ~v_1348 | ~v_1347 | ~v_1346 | ~v_1345 | ~v_1344 | ~v_1343 | ~v_1342 | ~v_1341 | ~v_1340 | ~v_1339 | ~v_1338 | ~v_1337 | ~v_1336 | ~v_1335 | ~v_1334 | ~v_1333 | ~v_1332 | ~v_1331 | ~v_1330 | ~v_1329 | v_1353;
assign x_27446 = v_1352 | v_152;
assign x_27447 = v_1352 | v_128;
assign x_27448 = v_1351 | v_153;
assign x_27449 = v_1351 | v_125;
assign x_27450 = v_1350 | v_154;
assign x_27451 = v_1350 | v_124;
assign x_27452 = v_1349 | ~v_152;
assign x_27453 = v_1349 | v_113;
assign x_27454 = v_1348 | ~v_153;
assign x_27455 = v_1348 | v_110;
assign x_27456 = v_1347 | ~v_154;
assign x_27457 = v_1347 | v_109;
assign x_27458 = v_1346 | v_154;
assign x_27459 = v_1346 | v_131;
assign x_27460 = v_1345 | v_154;
assign x_27461 = v_1345 | v_126;
assign x_27462 = v_1344 | ~v_154;
assign x_27463 = v_1344 | v_116;
assign x_27464 = v_1343 | ~v_154;
assign x_27465 = v_1343 | v_111;
assign x_27466 = v_1342 | v_156;
assign x_27467 = v_1342 | v_127;
assign x_27468 = v_1341 | v_157;
assign x_27469 = v_1341 | v_121;
assign x_27470 = v_1340 | v_158;
assign x_27471 = v_1340 | v_119;
assign x_27472 = v_1339 | ~v_156;
assign x_27473 = v_1339 | v_112;
assign x_27474 = v_1338 | ~v_157;
assign x_27475 = v_1338 | v_106;
assign x_27476 = v_1337 | ~v_158;
assign x_27477 = v_1337 | v_104;
assign x_27478 = v_1336 | v_177;
assign x_27479 = v_1336 | v_130;
assign x_27480 = v_1335 | v_178;
assign x_27481 = v_1335 | v_122;
assign x_27482 = v_1334 | ~v_177;
assign x_27483 = v_1334 | v_115;
assign x_27484 = v_1333 | ~v_178;
assign x_27485 = v_1333 | v_107;
assign x_27486 = v_1332 | v_177;
assign x_27487 = v_1332 | v_123;
assign x_27488 = v_1331 | v_178;
assign x_27489 = v_1331 | v_120;
assign x_27490 = v_1330 | ~v_177;
assign x_27491 = v_1330 | v_108;
assign x_27492 = v_1329 | ~v_178;
assign x_27493 = v_1329 | v_105;
assign x_27494 = v_56 | v_55 | v_61 | v_60 | v_59 | v_58 | v_145 | v_143 | v_142 | v_166 | v_165 | v_183 | ~v_604 | ~v_603 | ~v_266 | ~v_265 | ~v_420 | ~v_419 | ~v_602 | ~v_601 | ~v_1327 | ~v_1326 | ~v_1325 | ~v_1324 | ~v_1323 | ~v_1322 | ~v_1321 | ~v_1320 | ~v_1319 | ~v_1318 | ~v_1317 | ~v_1316 | ~v_1315 | ~v_1314 | ~v_1313 | ~v_1312 | ~v_1311 | ~v_1310 | ~v_1309 | ~v_1308 | ~v_1307 | ~v_1306 | ~v_1305 | ~v_1304 | v_1328;
assign x_27495 = v_1327 | v_152;
assign x_27496 = v_1327 | v_86;
assign x_27497 = v_1326 | v_153;
assign x_27498 = v_1326 | v_83;
assign x_27499 = v_1325 | v_154;
assign x_27500 = v_1325 | v_82;
assign x_27501 = v_1324 | ~v_152;
assign x_27502 = v_1324 | v_71;
assign x_27503 = v_1323 | ~v_153;
assign x_27504 = v_1323 | v_68;
assign x_27505 = v_1322 | ~v_154;
assign x_27506 = v_1322 | v_67;
assign x_27507 = v_1321 | v_154;
assign x_27508 = v_1321 | v_89;
assign x_27509 = v_1320 | v_154;
assign x_27510 = v_1320 | v_84;
assign x_27511 = v_1319 | ~v_154;
assign x_27512 = v_1319 | v_74;
assign x_27513 = v_1318 | ~v_154;
assign x_27514 = v_1318 | v_69;
assign x_27515 = v_1317 | v_156;
assign x_27516 = v_1317 | v_85;
assign x_27517 = v_1316 | v_157;
assign x_27518 = v_1316 | v_79;
assign x_27519 = v_1315 | v_158;
assign x_27520 = v_1315 | v_77;
assign x_27521 = v_1314 | ~v_156;
assign x_27522 = v_1314 | v_70;
assign x_27523 = v_1313 | ~v_157;
assign x_27524 = v_1313 | v_64;
assign x_27525 = v_1312 | ~v_158;
assign x_27526 = v_1312 | v_62;
assign x_27527 = v_1311 | v_177;
assign x_27528 = v_1311 | v_88;
assign x_27529 = v_1310 | v_178;
assign x_27530 = v_1310 | v_80;
assign x_27531 = v_1309 | ~v_177;
assign x_27532 = v_1309 | v_73;
assign x_27533 = v_1308 | ~v_178;
assign x_27534 = v_1308 | v_65;
assign x_27535 = v_1307 | v_177;
assign x_27536 = v_1307 | v_81;
assign x_27537 = v_1306 | v_178;
assign x_27538 = v_1306 | v_78;
assign x_27539 = v_1305 | ~v_177;
assign x_27540 = v_1305 | v_66;
assign x_27541 = v_1304 | ~v_178;
assign x_27542 = v_1304 | v_63;
assign x_27543 = v_13 | v_18 | v_17 | v_16 | v_15 | v_12 | v_135 | v_134 | v_137 | v_162 | v_161 | v_182 | ~v_599 | ~v_598 | ~v_233 | ~v_232 | ~v_405 | ~v_404 | ~v_597 | ~v_596 | ~v_1302 | ~v_1301 | ~v_1300 | ~v_1299 | ~v_1298 | ~v_1297 | ~v_1296 | ~v_1295 | ~v_1294 | ~v_1293 | ~v_1292 | ~v_1291 | ~v_1290 | ~v_1289 | ~v_1288 | ~v_1287 | ~v_1286 | ~v_1285 | ~v_1284 | ~v_1283 | ~v_1282 | ~v_1281 | ~v_1280 | ~v_1279 | v_1303;
assign x_27544 = v_1302 | v_152;
assign x_27545 = v_1302 | v_44;
assign x_27546 = v_1301 | v_153;
assign x_27547 = v_1301 | v_41;
assign x_27548 = v_1300 | v_154;
assign x_27549 = v_1300 | v_40;
assign x_27550 = v_1299 | ~v_152;
assign x_27551 = v_1299 | v_29;
assign x_27552 = v_1298 | ~v_153;
assign x_27553 = v_1298 | v_26;
assign x_27554 = v_1297 | ~v_154;
assign x_27555 = v_1297 | v_25;
assign x_27556 = v_1296 | v_154;
assign x_27557 = v_1296 | v_47;
assign x_27558 = v_1295 | v_154;
assign x_27559 = v_1295 | v_42;
assign x_27560 = v_1294 | ~v_154;
assign x_27561 = v_1294 | v_32;
assign x_27562 = v_1293 | ~v_154;
assign x_27563 = v_1293 | v_27;
assign x_27564 = v_1292 | v_156;
assign x_27565 = v_1292 | v_43;
assign x_27566 = v_1291 | v_157;
assign x_27567 = v_1291 | v_37;
assign x_27568 = v_1290 | v_158;
assign x_27569 = v_1290 | v_35;
assign x_27570 = v_1289 | ~v_156;
assign x_27571 = v_1289 | v_28;
assign x_27572 = v_1288 | ~v_157;
assign x_27573 = v_1288 | v_22;
assign x_27574 = v_1287 | ~v_158;
assign x_27575 = v_1287 | v_20;
assign x_27576 = v_1286 | v_177;
assign x_27577 = v_1286 | v_46;
assign x_27578 = v_1285 | v_178;
assign x_27579 = v_1285 | v_38;
assign x_27580 = v_1284 | ~v_177;
assign x_27581 = v_1284 | v_31;
assign x_27582 = v_1283 | ~v_178;
assign x_27583 = v_1283 | v_23;
assign x_27584 = v_1282 | v_177;
assign x_27585 = v_1282 | v_39;
assign x_27586 = v_1281 | v_178;
assign x_27587 = v_1281 | v_36;
assign x_27588 = v_1280 | ~v_177;
assign x_27589 = v_1280 | v_24;
assign x_27590 = v_1279 | ~v_178;
assign x_27591 = v_1279 | v_21;
assign x_27592 = v_1278 | ~v_1273;
assign x_27593 = v_1278 | ~v_1277;
assign x_27594 = v_1278 | ~v_199;
assign x_27595 = v_1278 | ~v_200;
assign x_27596 = v_1278 | ~v_178;
assign x_27597 = v_1278 | ~v_177;
assign x_27598 = ~v_185 | ~v_1276 | v_1277;
assign x_27599 = v_1276 | ~v_1274;
assign x_27600 = v_1276 | ~v_1275;
assign x_27601 = v_1276 | ~v_153;
assign x_27602 = v_1276 | ~v_152;
assign x_27603 = ~v_189 | ~v_186 | v_1275;
assign x_27604 = ~v_188 | ~v_185 | v_1274;
assign x_27605 = ~v_195 | ~v_1272 | v_1273;
assign x_27606 = v_1272 | ~v_1270;
assign x_27607 = v_1272 | ~v_1271;
assign x_27608 = v_1272 | ~v_174;
assign x_27609 = v_1272 | ~v_173;
assign x_27610 = ~v_186 | ~v_193 | v_1271;
assign x_27611 = ~v_188 | ~v_195 | v_1270;
assign x_27612 = v_1269 | ~v_726;
assign x_27613 = v_1269 | ~v_1268;
assign x_27614 = v_177 | v_178 | ~v_1267 | ~v_742 | ~v_741 | ~v_740 | ~v_734 | v_1268;
assign x_27615 = v_1267 | ~v_842;
assign x_27616 = v_1267 | ~v_888;
assign x_27617 = v_1267 | ~v_934;
assign x_27618 = v_1267 | ~v_980;
assign x_27619 = v_1267 | ~v_1026;
assign x_27620 = v_1267 | ~v_1042;
assign x_27621 = v_1267 | ~v_1088;
assign x_27622 = v_1267 | ~v_1104;
assign x_27623 = v_1267 | ~v_1120;
assign x_27624 = v_1267 | ~v_1136;
assign x_27625 = v_1267 | ~v_1152;
assign x_27626 = v_1267 | ~v_1198;
assign x_27627 = v_1267 | ~v_1214;
assign x_27628 = v_1267 | ~v_1230;
assign x_27629 = v_1267 | ~v_1246;
assign x_27630 = v_1267 | ~v_1262;
assign x_27631 = v_1267 | ~v_1263;
assign x_27632 = v_1267 | ~v_1264;
assign x_27633 = v_1267 | ~v_1265;
assign x_27634 = v_1267 | ~v_1266;
assign x_27635 = ~v_5 | v_4 | v_1266;
assign x_27636 = ~v_4 | v_6 | v_1265;
assign x_27637 = ~v_3 | v_2 | v_1264;
assign x_27638 = ~v_2 | v_1 | v_1263;
assign x_27639 = ~v_1261 | ~v_1256 | ~v_1251 | v_1262;
assign x_27640 = v_1261 | ~v_809;
assign x_27641 = v_1261 | ~v_810;
assign x_27642 = v_1261 | ~v_811;
assign x_27643 = v_1261 | ~v_812;
assign x_27644 = v_1261 | ~v_817;
assign x_27645 = v_1261 | ~v_818;
assign x_27646 = v_1261 | ~v_1011;
assign x_27647 = v_1261 | ~v_819;
assign x_27648 = v_1261 | ~v_1012;
assign x_27649 = v_1261 | ~v_820;
assign x_27650 = v_1261 | ~v_821;
assign x_27651 = v_1261 | ~v_1013;
assign x_27652 = v_1261 | ~v_822;
assign x_27653 = v_1261 | ~v_1014;
assign x_27654 = v_1261 | ~v_827;
assign x_27655 = v_1261 | ~v_828;
assign x_27656 = v_1261 | ~v_1015;
assign x_27657 = v_1261 | ~v_829;
assign x_27658 = v_1261 | ~v_1016;
assign x_27659 = v_1261 | ~v_830;
assign x_27660 = v_1261 | ~v_831;
assign x_27661 = v_1261 | ~v_1017;
assign x_27662 = v_1261 | ~v_832;
assign x_27663 = v_1261 | ~v_1018;
assign x_27664 = v_1261 | ~v_839;
assign x_27665 = v_1261 | ~v_1257;
assign x_27666 = v_1261 | ~v_1023;
assign x_27667 = v_1261 | ~v_840;
assign x_27668 = v_1261 | ~v_1258;
assign x_27669 = v_1261 | ~v_1024;
assign x_27670 = v_1261 | ~v_184;
assign x_27671 = v_1261 | ~v_170;
assign x_27672 = v_1261 | ~v_169;
assign x_27673 = v_1261 | ~v_149;
assign x_27674 = v_1261 | ~v_148;
assign x_27675 = v_1261 | ~v_1259;
assign x_27676 = v_1261 | ~v_1260;
assign x_27677 = v_1261 | ~v_103;
assign x_27678 = v_1261 | ~v_102;
assign x_27679 = v_1261 | ~v_101;
assign x_27680 = v_1261 | ~v_100;
assign x_27681 = v_1261 | ~v_99;
assign x_27682 = v_1261 | ~v_98;
assign x_27683 = v_1261 | ~v_95;
assign x_27684 = ~v_6 | ~v_19 | v_1260;
assign x_27685 = ~v_3 | v_19 | v_1259;
assign x_27686 = ~v_19 | ~v_132 | v_1258;
assign x_27687 = v_19 | ~v_117 | v_1257;
assign x_27688 = v_1256 | ~v_776;
assign x_27689 = v_1256 | ~v_777;
assign x_27690 = v_1256 | ~v_778;
assign x_27691 = v_1256 | ~v_779;
assign x_27692 = v_1256 | ~v_784;
assign x_27693 = v_1256 | ~v_785;
assign x_27694 = v_1256 | ~v_996;
assign x_27695 = v_1256 | ~v_786;
assign x_27696 = v_1256 | ~v_997;
assign x_27697 = v_1256 | ~v_787;
assign x_27698 = v_1256 | ~v_788;
assign x_27699 = v_1256 | ~v_998;
assign x_27700 = v_1256 | ~v_789;
assign x_27701 = v_1256 | ~v_999;
assign x_27702 = v_1256 | ~v_794;
assign x_27703 = v_1256 | ~v_795;
assign x_27704 = v_1256 | ~v_1000;
assign x_27705 = v_1256 | ~v_796;
assign x_27706 = v_1256 | ~v_1001;
assign x_27707 = v_1256 | ~v_797;
assign x_27708 = v_1256 | ~v_798;
assign x_27709 = v_1256 | ~v_1002;
assign x_27710 = v_1256 | ~v_799;
assign x_27711 = v_1256 | ~v_1003;
assign x_27712 = v_1256 | ~v_806;
assign x_27713 = v_1256 | ~v_1252;
assign x_27714 = v_1256 | ~v_1008;
assign x_27715 = v_1256 | ~v_1253;
assign x_27716 = v_1256 | ~v_1009;
assign x_27717 = v_1256 | ~v_807;
assign x_27718 = v_1256 | ~v_183;
assign x_27719 = v_1256 | ~v_166;
assign x_27720 = v_1256 | ~v_165;
assign x_27721 = v_1256 | ~v_144;
assign x_27722 = v_1256 | ~v_143;
assign x_27723 = v_1256 | ~v_1254;
assign x_27724 = v_1256 | ~v_1255;
assign x_27725 = v_1256 | ~v_61;
assign x_27726 = v_1256 | ~v_60;
assign x_27727 = v_1256 | ~v_59;
assign x_27728 = v_1256 | ~v_58;
assign x_27729 = v_1256 | ~v_57;
assign x_27730 = v_1256 | ~v_56;
assign x_27731 = v_1256 | ~v_53;
assign x_27732 = ~v_4 | ~v_19 | v_1255;
assign x_27733 = ~v_2 | v_19 | v_1254;
assign x_27734 = ~v_19 | ~v_90 | v_1253;
assign x_27735 = v_19 | ~v_75 | v_1252;
assign x_27736 = v_1251 | ~v_743;
assign x_27737 = v_1251 | ~v_744;
assign x_27738 = v_1251 | ~v_745;
assign x_27739 = v_1251 | ~v_746;
assign x_27740 = v_1251 | ~v_751;
assign x_27741 = v_1251 | ~v_752;
assign x_27742 = v_1251 | ~v_981;
assign x_27743 = v_1251 | ~v_753;
assign x_27744 = v_1251 | ~v_982;
assign x_27745 = v_1251 | ~v_754;
assign x_27746 = v_1251 | ~v_755;
assign x_27747 = v_1251 | ~v_983;
assign x_27748 = v_1251 | ~v_756;
assign x_27749 = v_1251 | ~v_984;
assign x_27750 = v_1251 | ~v_761;
assign x_27751 = v_1251 | ~v_762;
assign x_27752 = v_1251 | ~v_985;
assign x_27753 = v_1251 | ~v_763;
assign x_27754 = v_1251 | ~v_986;
assign x_27755 = v_1251 | ~v_764;
assign x_27756 = v_1251 | ~v_765;
assign x_27757 = v_1251 | ~v_987;
assign x_27758 = v_1251 | ~v_766;
assign x_27759 = v_1251 | ~v_988;
assign x_27760 = v_1251 | ~v_773;
assign x_27761 = v_1251 | ~v_774;
assign x_27762 = v_1251 | ~v_182;
assign x_27763 = v_1251 | ~v_162;
assign x_27764 = v_1251 | ~v_161;
assign x_27765 = v_1251 | ~v_1247;
assign x_27766 = v_1251 | ~v_1248;
assign x_27767 = v_1251 | ~v_136;
assign x_27768 = v_1251 | ~v_135;
assign x_27769 = v_1251 | ~v_1249;
assign x_27770 = v_1251 | ~v_993;
assign x_27771 = v_1251 | ~v_1250;
assign x_27772 = v_1251 | ~v_994;
assign x_27773 = v_1251 | ~v_18;
assign x_27774 = v_1251 | ~v_17;
assign x_27775 = v_1251 | ~v_16;
assign x_27776 = v_1251 | ~v_15;
assign x_27777 = v_1251 | ~v_14;
assign x_27778 = v_1251 | ~v_13;
assign x_27779 = v_1251 | ~v_10;
assign x_27780 = ~v_19 | ~v_48 | v_1250;
assign x_27781 = ~v_33 | v_19 | v_1249;
assign x_27782 = ~v_5 | ~v_19 | v_1248;
assign x_27783 = ~v_1 | v_19 | v_1247;
assign x_27784 = ~v_1245 | ~v_1240 | ~v_1235 | v_1246;
assign x_27785 = v_1245 | ~v_809;
assign x_27786 = v_1245 | ~v_810;
assign x_27787 = v_1245 | ~v_811;
assign x_27788 = v_1245 | ~v_812;
assign x_27789 = v_1245 | ~v_1183;
assign x_27790 = v_1245 | ~v_1184;
assign x_27791 = v_1245 | ~v_1185;
assign x_27792 = v_1245 | ~v_1186;
assign x_27793 = v_1245 | ~v_817;
assign x_27794 = v_1245 | ~v_1011;
assign x_27795 = v_1245 | ~v_1012;
assign x_27796 = v_1245 | ~v_820;
assign x_27797 = v_1245 | ~v_1013;
assign x_27798 = v_1245 | ~v_1014;
assign x_27799 = v_1245 | ~v_1187;
assign x_27800 = v_1245 | ~v_1188;
assign x_27801 = v_1245 | ~v_1189;
assign x_27802 = v_1245 | ~v_1190;
assign x_27803 = v_1245 | ~v_827;
assign x_27804 = v_1245 | ~v_1015;
assign x_27805 = v_1245 | ~v_1016;
assign x_27806 = v_1245 | ~v_830;
assign x_27807 = v_1245 | ~v_1017;
assign x_27808 = v_1245 | ~v_1018;
assign x_27809 = v_1245 | ~v_1193;
assign x_27810 = v_1245 | ~v_1241;
assign x_27811 = v_1245 | ~v_1194;
assign x_27812 = v_1245 | ~v_1242;
assign x_27813 = v_1245 | ~v_1023;
assign x_27814 = v_1245 | ~v_1024;
assign x_27815 = v_1245 | ~v_1243;
assign x_27816 = v_1245 | ~v_1244;
assign x_27817 = v_1245 | ~v_184;
assign x_27818 = v_1245 | ~v_171;
assign x_27819 = v_1245 | ~v_170;
assign x_27820 = v_1245 | ~v_149;
assign x_27821 = v_1245 | ~v_148;
assign x_27822 = v_1245 | ~v_147;
assign x_27823 = v_1245 | ~v_103;
assign x_27824 = v_1245 | ~v_102;
assign x_27825 = v_1245 | ~v_101;
assign x_27826 = v_1245 | ~v_100;
assign x_27827 = v_1245 | ~v_99;
assign x_27828 = v_1245 | ~v_93;
assign x_27829 = ~v_132 | ~v_152 | v_1244;
assign x_27830 = ~v_117 | v_152 | v_1243;
assign x_27831 = ~v_6 | ~v_153 | v_1242;
assign x_27832 = ~v_3 | v_153 | v_1241;
assign x_27833 = v_1240 | ~v_776;
assign x_27834 = v_1240 | ~v_777;
assign x_27835 = v_1240 | ~v_778;
assign x_27836 = v_1240 | ~v_779;
assign x_27837 = v_1240 | ~v_1168;
assign x_27838 = v_1240 | ~v_1169;
assign x_27839 = v_1240 | ~v_1170;
assign x_27840 = v_1240 | ~v_1171;
assign x_27841 = v_1240 | ~v_784;
assign x_27842 = v_1240 | ~v_996;
assign x_27843 = v_1240 | ~v_997;
assign x_27844 = v_1240 | ~v_787;
assign x_27845 = v_1240 | ~v_998;
assign x_27846 = v_1240 | ~v_999;
assign x_27847 = v_1240 | ~v_1172;
assign x_27848 = v_1240 | ~v_1173;
assign x_27849 = v_1240 | ~v_1174;
assign x_27850 = v_1240 | ~v_1175;
assign x_27851 = v_1240 | ~v_794;
assign x_27852 = v_1240 | ~v_1000;
assign x_27853 = v_1240 | ~v_1001;
assign x_27854 = v_1240 | ~v_797;
assign x_27855 = v_1240 | ~v_1002;
assign x_27856 = v_1240 | ~v_1003;
assign x_27857 = v_1240 | ~v_1178;
assign x_27858 = v_1240 | ~v_1236;
assign x_27859 = v_1240 | ~v_1179;
assign x_27860 = v_1240 | ~v_1237;
assign x_27861 = v_1240 | ~v_1008;
assign x_27862 = v_1240 | ~v_1009;
assign x_27863 = v_1240 | ~v_1238;
assign x_27864 = v_1240 | ~v_1239;
assign x_27865 = v_1240 | ~v_183;
assign x_27866 = v_1240 | ~v_167;
assign x_27867 = v_1240 | ~v_166;
assign x_27868 = v_1240 | ~v_144;
assign x_27869 = v_1240 | ~v_143;
assign x_27870 = v_1240 | ~v_142;
assign x_27871 = v_1240 | ~v_61;
assign x_27872 = v_1240 | ~v_60;
assign x_27873 = v_1240 | ~v_59;
assign x_27874 = v_1240 | ~v_58;
assign x_27875 = v_1240 | ~v_57;
assign x_27876 = v_1240 | ~v_51;
assign x_27877 = ~v_90 | ~v_152 | v_1239;
assign x_27878 = ~v_75 | v_152 | v_1238;
assign x_27879 = ~v_4 | ~v_153 | v_1237;
assign x_27880 = ~v_2 | v_153 | v_1236;
assign x_27881 = v_1235 | ~v_743;
assign x_27882 = v_1235 | ~v_744;
assign x_27883 = v_1235 | ~v_745;
assign x_27884 = v_1235 | ~v_746;
assign x_27885 = v_1235 | ~v_1153;
assign x_27886 = v_1235 | ~v_1154;
assign x_27887 = v_1235 | ~v_1155;
assign x_27888 = v_1235 | ~v_1156;
assign x_27889 = v_1235 | ~v_751;
assign x_27890 = v_1235 | ~v_981;
assign x_27891 = v_1235 | ~v_982;
assign x_27892 = v_1235 | ~v_754;
assign x_27893 = v_1235 | ~v_983;
assign x_27894 = v_1235 | ~v_984;
assign x_27895 = v_1235 | ~v_1157;
assign x_27896 = v_1235 | ~v_1158;
assign x_27897 = v_1235 | ~v_1159;
assign x_27898 = v_1235 | ~v_1160;
assign x_27899 = v_1235 | ~v_761;
assign x_27900 = v_1235 | ~v_985;
assign x_27901 = v_1235 | ~v_986;
assign x_27902 = v_1235 | ~v_764;
assign x_27903 = v_1235 | ~v_987;
assign x_27904 = v_1235 | ~v_988;
assign x_27905 = v_1235 | ~v_1163;
assign x_27906 = v_1235 | ~v_1231;
assign x_27907 = v_1235 | ~v_1164;
assign x_27908 = v_1235 | ~v_1232;
assign x_27909 = v_1235 | ~v_1233;
assign x_27910 = v_1235 | ~v_1234;
assign x_27911 = v_1235 | ~v_182;
assign x_27912 = v_1235 | ~v_163;
assign x_27913 = v_1235 | ~v_162;
assign x_27914 = v_1235 | ~v_136;
assign x_27915 = v_1235 | ~v_135;
assign x_27916 = v_1235 | ~v_134;
assign x_27917 = v_1235 | ~v_993;
assign x_27918 = v_1235 | ~v_994;
assign x_27919 = v_1235 | ~v_18;
assign x_27920 = v_1235 | ~v_17;
assign x_27921 = v_1235 | ~v_16;
assign x_27922 = v_1235 | ~v_15;
assign x_27923 = v_1235 | ~v_14;
assign x_27924 = v_1235 | ~v_8;
assign x_27925 = ~v_48 | ~v_152 | v_1234;
assign x_27926 = ~v_33 | v_152 | v_1233;
assign x_27927 = ~v_5 | ~v_153 | v_1232;
assign x_27928 = ~v_1 | v_153 | v_1231;
assign x_27929 = ~v_1229 | ~v_1224 | ~v_1219 | v_1230;
assign x_27930 = v_1229 | ~v_809;
assign x_27931 = v_1229 | ~v_810;
assign x_27932 = v_1229 | ~v_811;
assign x_27933 = v_1229 | ~v_812;
assign x_27934 = v_1229 | ~v_1183;
assign x_27935 = v_1229 | ~v_1184;
assign x_27936 = v_1229 | ~v_1185;
assign x_27937 = v_1229 | ~v_1186;
assign x_27938 = v_1229 | ~v_965;
assign x_27939 = v_1229 | ~v_966;
assign x_27940 = v_1229 | ~v_967;
assign x_27941 = v_1229 | ~v_968;
assign x_27942 = v_1229 | ~v_817;
assign x_27943 = v_1229 | ~v_820;
assign x_27944 = v_1229 | ~v_969;
assign x_27945 = v_1229 | ~v_970;
assign x_27946 = v_1229 | ~v_971;
assign x_27947 = v_1229 | ~v_972;
assign x_27948 = v_1229 | ~v_1187;
assign x_27949 = v_1229 | ~v_1188;
assign x_27950 = v_1229 | ~v_1189;
assign x_27951 = v_1229 | ~v_1190;
assign x_27952 = v_1229 | ~v_827;
assign x_27953 = v_1229 | ~v_830;
assign x_27954 = v_1229 | ~v_1225;
assign x_27955 = v_1229 | ~v_1226;
assign x_27956 = v_1229 | ~v_1227;
assign x_27957 = v_1229 | ~v_1228;
assign x_27958 = v_1229 | ~v_1193;
assign x_27959 = v_1229 | ~v_1194;
assign x_27960 = v_1229 | ~v_975;
assign x_27961 = v_1229 | ~v_976;
assign x_27962 = v_1229 | ~v_184;
assign x_27963 = v_1229 | ~v_171;
assign x_27964 = v_1229 | ~v_170;
assign x_27965 = v_1229 | ~v_150;
assign x_27966 = v_1229 | ~v_149;
assign x_27967 = v_1229 | ~v_103;
assign x_27968 = v_1229 | ~v_102;
assign x_27969 = v_1229 | ~v_101;
assign x_27970 = v_1229 | ~v_100;
assign x_27971 = v_1229 | ~v_96;
assign x_27972 = v_1229 | ~v_95;
assign x_27973 = v_1229 | ~v_93;
assign x_27974 = ~v_132 | ~v_154 | v_1228;
assign x_27975 = ~v_6 | ~v_154 | v_1227;
assign x_27976 = ~v_117 | v_154 | v_1226;
assign x_27977 = ~v_3 | v_154 | v_1225;
assign x_27978 = v_1224 | ~v_776;
assign x_27979 = v_1224 | ~v_777;
assign x_27980 = v_1224 | ~v_778;
assign x_27981 = v_1224 | ~v_779;
assign x_27982 = v_1224 | ~v_1168;
assign x_27983 = v_1224 | ~v_1169;
assign x_27984 = v_1224 | ~v_1170;
assign x_27985 = v_1224 | ~v_1171;
assign x_27986 = v_1224 | ~v_950;
assign x_27987 = v_1224 | ~v_951;
assign x_27988 = v_1224 | ~v_952;
assign x_27989 = v_1224 | ~v_953;
assign x_27990 = v_1224 | ~v_784;
assign x_27991 = v_1224 | ~v_787;
assign x_27992 = v_1224 | ~v_954;
assign x_27993 = v_1224 | ~v_955;
assign x_27994 = v_1224 | ~v_956;
assign x_27995 = v_1224 | ~v_957;
assign x_27996 = v_1224 | ~v_1172;
assign x_27997 = v_1224 | ~v_1173;
assign x_27998 = v_1224 | ~v_1174;
assign x_27999 = v_1224 | ~v_1175;
assign x_28000 = v_1224 | ~v_794;
assign x_28001 = v_1224 | ~v_797;
assign x_28002 = v_1224 | ~v_1220;
assign x_28003 = v_1224 | ~v_1221;
assign x_28004 = v_1224 | ~v_1222;
assign x_28005 = v_1224 | ~v_1223;
assign x_28006 = v_1224 | ~v_1178;
assign x_28007 = v_1224 | ~v_1179;
assign x_28008 = v_1224 | ~v_960;
assign x_28009 = v_1224 | ~v_961;
assign x_28010 = v_1224 | ~v_183;
assign x_28011 = v_1224 | ~v_167;
assign x_28012 = v_1224 | ~v_166;
assign x_28013 = v_1224 | ~v_145;
assign x_28014 = v_1224 | ~v_144;
assign x_28015 = v_1224 | ~v_61;
assign x_28016 = v_1224 | ~v_60;
assign x_28017 = v_1224 | ~v_59;
assign x_28018 = v_1224 | ~v_58;
assign x_28019 = v_1224 | ~v_54;
assign x_28020 = v_1224 | ~v_53;
assign x_28021 = v_1224 | ~v_51;
assign x_28022 = ~v_90 | ~v_154 | v_1223;
assign x_28023 = ~v_4 | ~v_154 | v_1222;
assign x_28024 = ~v_75 | v_154 | v_1221;
assign x_28025 = ~v_2 | v_154 | v_1220;
assign x_28026 = v_1219 | ~v_743;
assign x_28027 = v_1219 | ~v_744;
assign x_28028 = v_1219 | ~v_745;
assign x_28029 = v_1219 | ~v_746;
assign x_28030 = v_1219 | ~v_1153;
assign x_28031 = v_1219 | ~v_1154;
assign x_28032 = v_1219 | ~v_1155;
assign x_28033 = v_1219 | ~v_1156;
assign x_28034 = v_1219 | ~v_935;
assign x_28035 = v_1219 | ~v_936;
assign x_28036 = v_1219 | ~v_937;
assign x_28037 = v_1219 | ~v_938;
assign x_28038 = v_1219 | ~v_751;
assign x_28039 = v_1219 | ~v_754;
assign x_28040 = v_1219 | ~v_939;
assign x_28041 = v_1219 | ~v_940;
assign x_28042 = v_1219 | ~v_941;
assign x_28043 = v_1219 | ~v_942;
assign x_28044 = v_1219 | ~v_1157;
assign x_28045 = v_1219 | ~v_1158;
assign x_28046 = v_1219 | ~v_1159;
assign x_28047 = v_1219 | ~v_1160;
assign x_28048 = v_1219 | ~v_761;
assign x_28049 = v_1219 | ~v_764;
assign x_28050 = v_1219 | ~v_1215;
assign x_28051 = v_1219 | ~v_1216;
assign x_28052 = v_1219 | ~v_1217;
assign x_28053 = v_1219 | ~v_1218;
assign x_28054 = v_1219 | ~v_1163;
assign x_28055 = v_1219 | ~v_1164;
assign x_28056 = v_1219 | ~v_945;
assign x_28057 = v_1219 | ~v_946;
assign x_28058 = v_1219 | ~v_182;
assign x_28059 = v_1219 | ~v_163;
assign x_28060 = v_1219 | ~v_162;
assign x_28061 = v_1219 | ~v_137;
assign x_28062 = v_1219 | ~v_136;
assign x_28063 = v_1219 | ~v_18;
assign x_28064 = v_1219 | ~v_17;
assign x_28065 = v_1219 | ~v_16;
assign x_28066 = v_1219 | ~v_15;
assign x_28067 = v_1219 | ~v_11;
assign x_28068 = v_1219 | ~v_10;
assign x_28069 = v_1219 | ~v_8;
assign x_28070 = ~v_48 | ~v_154 | v_1218;
assign x_28071 = ~v_5 | ~v_154 | v_1217;
assign x_28072 = ~v_33 | v_154 | v_1216;
assign x_28073 = ~v_1 | v_154 | v_1215;
assign x_28074 = ~v_1213 | ~v_1208 | ~v_1203 | v_1214;
assign x_28075 = v_1213 | ~v_809;
assign x_28076 = v_1213 | ~v_810;
assign x_28077 = v_1213 | ~v_811;
assign x_28078 = v_1213 | ~v_812;
assign x_28079 = v_1213 | ~v_1183;
assign x_28080 = v_1213 | ~v_1184;
assign x_28081 = v_1213 | ~v_1185;
assign x_28082 = v_1213 | ~v_1186;
assign x_28083 = v_1213 | ~v_919;
assign x_28084 = v_1213 | ~v_920;
assign x_28085 = v_1213 | ~v_817;
assign x_28086 = v_1213 | ~v_820;
assign x_28087 = v_1213 | ~v_921;
assign x_28088 = v_1213 | ~v_922;
assign x_28089 = v_1213 | ~v_923;
assign x_28090 = v_1213 | ~v_924;
assign x_28091 = v_1213 | ~v_1187;
assign x_28092 = v_1213 | ~v_1188;
assign x_28093 = v_1213 | ~v_1189;
assign x_28094 = v_1213 | ~v_1190;
assign x_28095 = v_1213 | ~v_827;
assign x_28096 = v_1213 | ~v_830;
assign x_28097 = v_1213 | ~v_1209;
assign x_28098 = v_1213 | ~v_1210;
assign x_28099 = v_1213 | ~v_1193;
assign x_28100 = v_1213 | ~v_1194;
assign x_28101 = v_1213 | ~v_927;
assign x_28102 = v_1213 | ~v_928;
assign x_28103 = v_1213 | ~v_931;
assign x_28104 = v_1213 | ~v_932;
assign x_28105 = v_1213 | ~v_1211;
assign x_28106 = v_1213 | ~v_1212;
assign x_28107 = v_1213 | ~v_184;
assign x_28108 = v_1213 | ~v_172;
assign x_28109 = v_1213 | ~v_171;
assign x_28110 = v_1213 | ~v_170;
assign x_28111 = v_1213 | ~v_150;
assign x_28112 = v_1213 | ~v_149;
assign x_28113 = v_1213 | ~v_148;
assign x_28114 = v_1213 | ~v_147;
assign x_28115 = v_1213 | ~v_102;
assign x_28116 = v_1213 | ~v_101;
assign x_28117 = v_1213 | ~v_100;
assign x_28118 = v_1213 | ~v_93;
assign x_28119 = ~v_132 | ~v_173 | v_1212;
assign x_28120 = ~v_117 | v_173 | v_1211;
assign x_28121 = ~v_6 | ~v_174 | v_1210;
assign x_28122 = ~v_3 | v_174 | v_1209;
assign x_28123 = v_1208 | ~v_776;
assign x_28124 = v_1208 | ~v_777;
assign x_28125 = v_1208 | ~v_778;
assign x_28126 = v_1208 | ~v_779;
assign x_28127 = v_1208 | ~v_1168;
assign x_28128 = v_1208 | ~v_1169;
assign x_28129 = v_1208 | ~v_1170;
assign x_28130 = v_1208 | ~v_1171;
assign x_28131 = v_1208 | ~v_904;
assign x_28132 = v_1208 | ~v_905;
assign x_28133 = v_1208 | ~v_784;
assign x_28134 = v_1208 | ~v_787;
assign x_28135 = v_1208 | ~v_906;
assign x_28136 = v_1208 | ~v_907;
assign x_28137 = v_1208 | ~v_908;
assign x_28138 = v_1208 | ~v_909;
assign x_28139 = v_1208 | ~v_1172;
assign x_28140 = v_1208 | ~v_1173;
assign x_28141 = v_1208 | ~v_1174;
assign x_28142 = v_1208 | ~v_1175;
assign x_28143 = v_1208 | ~v_794;
assign x_28144 = v_1208 | ~v_797;
assign x_28145 = v_1208 | ~v_1204;
assign x_28146 = v_1208 | ~v_1205;
assign x_28147 = v_1208 | ~v_1178;
assign x_28148 = v_1208 | ~v_1179;
assign x_28149 = v_1208 | ~v_912;
assign x_28150 = v_1208 | ~v_913;
assign x_28151 = v_1208 | ~v_916;
assign x_28152 = v_1208 | ~v_917;
assign x_28153 = v_1208 | ~v_1206;
assign x_28154 = v_1208 | ~v_1207;
assign x_28155 = v_1208 | ~v_183;
assign x_28156 = v_1208 | ~v_168;
assign x_28157 = v_1208 | ~v_167;
assign x_28158 = v_1208 | ~v_166;
assign x_28159 = v_1208 | ~v_145;
assign x_28160 = v_1208 | ~v_144;
assign x_28161 = v_1208 | ~v_143;
assign x_28162 = v_1208 | ~v_142;
assign x_28163 = v_1208 | ~v_60;
assign x_28164 = v_1208 | ~v_59;
assign x_28165 = v_1208 | ~v_58;
assign x_28166 = v_1208 | ~v_51;
assign x_28167 = ~v_90 | ~v_173 | v_1207;
assign x_28168 = ~v_75 | v_173 | v_1206;
assign x_28169 = ~v_4 | ~v_174 | v_1205;
assign x_28170 = ~v_2 | v_174 | v_1204;
assign x_28171 = v_1203 | ~v_743;
assign x_28172 = v_1203 | ~v_744;
assign x_28173 = v_1203 | ~v_745;
assign x_28174 = v_1203 | ~v_746;
assign x_28175 = v_1203 | ~v_1153;
assign x_28176 = v_1203 | ~v_1154;
assign x_28177 = v_1203 | ~v_1155;
assign x_28178 = v_1203 | ~v_1156;
assign x_28179 = v_1203 | ~v_889;
assign x_28180 = v_1203 | ~v_890;
assign x_28181 = v_1203 | ~v_751;
assign x_28182 = v_1203 | ~v_754;
assign x_28183 = v_1203 | ~v_891;
assign x_28184 = v_1203 | ~v_892;
assign x_28185 = v_1203 | ~v_893;
assign x_28186 = v_1203 | ~v_894;
assign x_28187 = v_1203 | ~v_1157;
assign x_28188 = v_1203 | ~v_1158;
assign x_28189 = v_1203 | ~v_1159;
assign x_28190 = v_1203 | ~v_1160;
assign x_28191 = v_1203 | ~v_761;
assign x_28192 = v_1203 | ~v_764;
assign x_28193 = v_1203 | ~v_1199;
assign x_28194 = v_1203 | ~v_1200;
assign x_28195 = v_1203 | ~v_1163;
assign x_28196 = v_1203 | ~v_1164;
assign x_28197 = v_1203 | ~v_897;
assign x_28198 = v_1203 | ~v_898;
assign x_28199 = v_1203 | ~v_901;
assign x_28200 = v_1203 | ~v_902;
assign x_28201 = v_1203 | ~v_1201;
assign x_28202 = v_1203 | ~v_1202;
assign x_28203 = v_1203 | ~v_182;
assign x_28204 = v_1203 | ~v_164;
assign x_28205 = v_1203 | ~v_163;
assign x_28206 = v_1203 | ~v_162;
assign x_28207 = v_1203 | ~v_137;
assign x_28208 = v_1203 | ~v_136;
assign x_28209 = v_1203 | ~v_135;
assign x_28210 = v_1203 | ~v_134;
assign x_28211 = v_1203 | ~v_17;
assign x_28212 = v_1203 | ~v_16;
assign x_28213 = v_1203 | ~v_15;
assign x_28214 = v_1203 | ~v_8;
assign x_28215 = ~v_48 | ~v_173 | v_1202;
assign x_28216 = ~v_33 | v_173 | v_1201;
assign x_28217 = ~v_5 | ~v_174 | v_1200;
assign x_28218 = ~v_1 | v_174 | v_1199;
assign x_28219 = ~v_1197 | ~v_1182 | ~v_1167 | v_1198;
assign x_28220 = v_1197 | ~v_809;
assign x_28221 = v_1197 | ~v_810;
assign x_28222 = v_1197 | ~v_811;
assign x_28223 = v_1197 | ~v_812;
assign x_28224 = v_1197 | ~v_1183;
assign x_28225 = v_1197 | ~v_1184;
assign x_28226 = v_1197 | ~v_1185;
assign x_28227 = v_1197 | ~v_1186;
assign x_28228 = v_1197 | ~v_813;
assign x_28229 = v_1197 | ~v_814;
assign x_28230 = v_1197 | ~v_815;
assign x_28231 = v_1197 | ~v_816;
assign x_28232 = v_1197 | ~v_817;
assign x_28233 = v_1197 | ~v_820;
assign x_28234 = v_1197 | ~v_823;
assign x_28235 = v_1197 | ~v_824;
assign x_28236 = v_1197 | ~v_825;
assign x_28237 = v_1197 | ~v_826;
assign x_28238 = v_1197 | ~v_1187;
assign x_28239 = v_1197 | ~v_1188;
assign x_28240 = v_1197 | ~v_1189;
assign x_28241 = v_1197 | ~v_1190;
assign x_28242 = v_1197 | ~v_827;
assign x_28243 = v_1197 | ~v_830;
assign x_28244 = v_1197 | ~v_1191;
assign x_28245 = v_1197 | ~v_1192;
assign x_28246 = v_1197 | ~v_1193;
assign x_28247 = v_1197 | ~v_1194;
assign x_28248 = v_1197 | ~v_837;
assign x_28249 = v_1197 | ~v_838;
assign x_28250 = v_1197 | ~v_1195;
assign x_28251 = v_1197 | ~v_1196;
assign x_28252 = v_1197 | ~v_184;
assign x_28253 = v_1197 | ~v_171;
assign x_28254 = v_1197 | ~v_170;
assign x_28255 = v_1197 | ~v_160;
assign x_28256 = v_1197 | ~v_151;
assign x_28257 = v_1197 | ~v_150;
assign x_28258 = v_1197 | ~v_148;
assign x_28259 = v_1197 | ~v_147;
assign x_28260 = v_1197 | ~v_103;
assign x_28261 = v_1197 | ~v_100;
assign x_28262 = v_1197 | ~v_97;
assign x_28263 = v_1197 | ~v_93;
assign x_28264 = ~v_132 | ~v_178 | v_1196;
assign x_28265 = ~v_117 | v_178 | v_1195;
assign x_28266 = ~v_129 | ~v_154 | v_1194;
assign x_28267 = ~v_114 | v_154 | v_1193;
assign x_28268 = ~v_6 | ~v_177 | v_1192;
assign x_28269 = ~v_3 | v_177 | v_1191;
assign x_28270 = ~v_127 | ~v_154 | v_1190;
assign x_28271 = ~v_121 | ~v_154 | v_1189;
assign x_28272 = ~v_112 | v_154 | v_1188;
assign x_28273 = ~v_106 | v_154 | v_1187;
assign x_28274 = ~v_128 | ~v_177 | v_1186;
assign x_28275 = ~v_125 | ~v_178 | v_1185;
assign x_28276 = ~v_113 | v_177 | v_1184;
assign x_28277 = ~v_110 | v_178 | v_1183;
assign x_28278 = v_1182 | ~v_776;
assign x_28279 = v_1182 | ~v_777;
assign x_28280 = v_1182 | ~v_778;
assign x_28281 = v_1182 | ~v_779;
assign x_28282 = v_1182 | ~v_1168;
assign x_28283 = v_1182 | ~v_1169;
assign x_28284 = v_1182 | ~v_1170;
assign x_28285 = v_1182 | ~v_1171;
assign x_28286 = v_1182 | ~v_780;
assign x_28287 = v_1182 | ~v_781;
assign x_28288 = v_1182 | ~v_782;
assign x_28289 = v_1182 | ~v_783;
assign x_28290 = v_1182 | ~v_784;
assign x_28291 = v_1182 | ~v_787;
assign x_28292 = v_1182 | ~v_790;
assign x_28293 = v_1182 | ~v_791;
assign x_28294 = v_1182 | ~v_792;
assign x_28295 = v_1182 | ~v_793;
assign x_28296 = v_1182 | ~v_1172;
assign x_28297 = v_1182 | ~v_1173;
assign x_28298 = v_1182 | ~v_1174;
assign x_28299 = v_1182 | ~v_1175;
assign x_28300 = v_1182 | ~v_794;
assign x_28301 = v_1182 | ~v_797;
assign x_28302 = v_1182 | ~v_1176;
assign x_28303 = v_1182 | ~v_1177;
assign x_28304 = v_1182 | ~v_1178;
assign x_28305 = v_1182 | ~v_1179;
assign x_28306 = v_1182 | ~v_804;
assign x_28307 = v_1182 | ~v_805;
assign x_28308 = v_1182 | ~v_1180;
assign x_28309 = v_1182 | ~v_1181;
assign x_28310 = v_1182 | ~v_183;
assign x_28311 = v_1182 | ~v_167;
assign x_28312 = v_1182 | ~v_166;
assign x_28313 = v_1182 | ~v_159;
assign x_28314 = v_1182 | ~v_146;
assign x_28315 = v_1182 | ~v_145;
assign x_28316 = v_1182 | ~v_143;
assign x_28317 = v_1182 | ~v_142;
assign x_28318 = v_1182 | ~v_61;
assign x_28319 = v_1182 | ~v_58;
assign x_28320 = v_1182 | ~v_55;
assign x_28321 = v_1182 | ~v_51;
assign x_28322 = ~v_90 | ~v_178 | v_1181;
assign x_28323 = ~v_75 | v_178 | v_1180;
assign x_28324 = ~v_87 | ~v_154 | v_1179;
assign x_28325 = ~v_72 | v_154 | v_1178;
assign x_28326 = ~v_4 | ~v_177 | v_1177;
assign x_28327 = ~v_2 | v_177 | v_1176;
assign x_28328 = ~v_85 | ~v_154 | v_1175;
assign x_28329 = ~v_79 | ~v_154 | v_1174;
assign x_28330 = ~v_70 | v_154 | v_1173;
assign x_28331 = ~v_64 | v_154 | v_1172;
assign x_28332 = ~v_86 | ~v_177 | v_1171;
assign x_28333 = ~v_83 | ~v_178 | v_1170;
assign x_28334 = ~v_71 | v_177 | v_1169;
assign x_28335 = ~v_68 | v_178 | v_1168;
assign x_28336 = v_1167 | ~v_743;
assign x_28337 = v_1167 | ~v_744;
assign x_28338 = v_1167 | ~v_745;
assign x_28339 = v_1167 | ~v_746;
assign x_28340 = v_1167 | ~v_1153;
assign x_28341 = v_1167 | ~v_1154;
assign x_28342 = v_1167 | ~v_1155;
assign x_28343 = v_1167 | ~v_1156;
assign x_28344 = v_1167 | ~v_747;
assign x_28345 = v_1167 | ~v_748;
assign x_28346 = v_1167 | ~v_749;
assign x_28347 = v_1167 | ~v_750;
assign x_28348 = v_1167 | ~v_751;
assign x_28349 = v_1167 | ~v_754;
assign x_28350 = v_1167 | ~v_757;
assign x_28351 = v_1167 | ~v_758;
assign x_28352 = v_1167 | ~v_759;
assign x_28353 = v_1167 | ~v_760;
assign x_28354 = v_1167 | ~v_1157;
assign x_28355 = v_1167 | ~v_1158;
assign x_28356 = v_1167 | ~v_1159;
assign x_28357 = v_1167 | ~v_1160;
assign x_28358 = v_1167 | ~v_761;
assign x_28359 = v_1167 | ~v_764;
assign x_28360 = v_1167 | ~v_1161;
assign x_28361 = v_1167 | ~v_1162;
assign x_28362 = v_1167 | ~v_1163;
assign x_28363 = v_1167 | ~v_1164;
assign x_28364 = v_1167 | ~v_771;
assign x_28365 = v_1167 | ~v_772;
assign x_28366 = v_1167 | ~v_1165;
assign x_28367 = v_1167 | ~v_1166;
assign x_28368 = v_1167 | ~v_182;
assign x_28369 = v_1167 | ~v_163;
assign x_28370 = v_1167 | ~v_162;
assign x_28371 = v_1167 | ~v_155;
assign x_28372 = v_1167 | ~v_138;
assign x_28373 = v_1167 | ~v_137;
assign x_28374 = v_1167 | ~v_135;
assign x_28375 = v_1167 | ~v_134;
assign x_28376 = v_1167 | ~v_18;
assign x_28377 = v_1167 | ~v_15;
assign x_28378 = v_1167 | ~v_12;
assign x_28379 = v_1167 | ~v_8;
assign x_28380 = ~v_48 | ~v_178 | v_1166;
assign x_28381 = ~v_33 | v_178 | v_1165;
assign x_28382 = ~v_45 | ~v_154 | v_1164;
assign x_28383 = ~v_30 | v_154 | v_1163;
assign x_28384 = ~v_5 | ~v_177 | v_1162;
assign x_28385 = ~v_1 | v_177 | v_1161;
assign x_28386 = ~v_43 | ~v_154 | v_1160;
assign x_28387 = ~v_37 | ~v_154 | v_1159;
assign x_28388 = ~v_28 | v_154 | v_1158;
assign x_28389 = ~v_22 | v_154 | v_1157;
assign x_28390 = ~v_44 | ~v_177 | v_1156;
assign x_28391 = ~v_41 | ~v_178 | v_1155;
assign x_28392 = ~v_29 | v_177 | v_1154;
assign x_28393 = ~v_26 | v_178 | v_1153;
assign x_28394 = ~v_1151 | ~v_1146 | ~v_1141 | v_1152;
assign x_28395 = v_1151 | ~v_809;
assign x_28396 = v_1151 | ~v_810;
assign x_28397 = v_1151 | ~v_811;
assign x_28398 = v_1151 | ~v_812;
assign x_28399 = v_1151 | ~v_965;
assign x_28400 = v_1151 | ~v_966;
assign x_28401 = v_1151 | ~v_967;
assign x_28402 = v_1151 | ~v_968;
assign x_28403 = v_1151 | ~v_817;
assign x_28404 = v_1151 | ~v_818;
assign x_28405 = v_1151 | ~v_819;
assign x_28406 = v_1151 | ~v_820;
assign x_28407 = v_1151 | ~v_821;
assign x_28408 = v_1151 | ~v_822;
assign x_28409 = v_1151 | ~v_969;
assign x_28410 = v_1151 | ~v_970;
assign x_28411 = v_1151 | ~v_971;
assign x_28412 = v_1151 | ~v_972;
assign x_28413 = v_1151 | ~v_827;
assign x_28414 = v_1151 | ~v_828;
assign x_28415 = v_1151 | ~v_829;
assign x_28416 = v_1151 | ~v_830;
assign x_28417 = v_1151 | ~v_831;
assign x_28418 = v_1151 | ~v_832;
assign x_28419 = v_1151 | ~v_1147;
assign x_28420 = v_1151 | ~v_1148;
assign x_28421 = v_1151 | ~v_975;
assign x_28422 = v_1151 | ~v_976;
assign x_28423 = v_1151 | ~v_839;
assign x_28424 = v_1151 | ~v_840;
assign x_28425 = v_1151 | ~v_1149;
assign x_28426 = v_1151 | ~v_1150;
assign x_28427 = v_1151 | ~v_184;
assign x_28428 = v_1151 | ~v_170;
assign x_28429 = v_1151 | ~v_169;
assign x_28430 = v_1151 | ~v_150;
assign x_28431 = v_1151 | ~v_149;
assign x_28432 = v_1151 | ~v_147;
assign x_28433 = v_1151 | ~v_103;
assign x_28434 = v_1151 | ~v_102;
assign x_28435 = v_1151 | ~v_101;
assign x_28436 = v_1151 | ~v_100;
assign x_28437 = v_1151 | ~v_98;
assign x_28438 = v_1151 | ~v_96;
assign x_28439 = ~v_117 | v_153 | v_1150;
assign x_28440 = ~v_132 | ~v_153 | v_1149;
assign x_28441 = ~v_6 | ~v_152 | v_1148;
assign x_28442 = ~v_3 | v_152 | v_1147;
assign x_28443 = v_1146 | ~v_776;
assign x_28444 = v_1146 | ~v_777;
assign x_28445 = v_1146 | ~v_778;
assign x_28446 = v_1146 | ~v_779;
assign x_28447 = v_1146 | ~v_950;
assign x_28448 = v_1146 | ~v_951;
assign x_28449 = v_1146 | ~v_952;
assign x_28450 = v_1146 | ~v_953;
assign x_28451 = v_1146 | ~v_784;
assign x_28452 = v_1146 | ~v_785;
assign x_28453 = v_1146 | ~v_786;
assign x_28454 = v_1146 | ~v_787;
assign x_28455 = v_1146 | ~v_788;
assign x_28456 = v_1146 | ~v_789;
assign x_28457 = v_1146 | ~v_954;
assign x_28458 = v_1146 | ~v_955;
assign x_28459 = v_1146 | ~v_956;
assign x_28460 = v_1146 | ~v_957;
assign x_28461 = v_1146 | ~v_794;
assign x_28462 = v_1146 | ~v_795;
assign x_28463 = v_1146 | ~v_796;
assign x_28464 = v_1146 | ~v_797;
assign x_28465 = v_1146 | ~v_798;
assign x_28466 = v_1146 | ~v_799;
assign x_28467 = v_1146 | ~v_1142;
assign x_28468 = v_1146 | ~v_1143;
assign x_28469 = v_1146 | ~v_960;
assign x_28470 = v_1146 | ~v_961;
assign x_28471 = v_1146 | ~v_806;
assign x_28472 = v_1146 | ~v_807;
assign x_28473 = v_1146 | ~v_1144;
assign x_28474 = v_1146 | ~v_1145;
assign x_28475 = v_1146 | ~v_183;
assign x_28476 = v_1146 | ~v_166;
assign x_28477 = v_1146 | ~v_165;
assign x_28478 = v_1146 | ~v_145;
assign x_28479 = v_1146 | ~v_144;
assign x_28480 = v_1146 | ~v_142;
assign x_28481 = v_1146 | ~v_61;
assign x_28482 = v_1146 | ~v_60;
assign x_28483 = v_1146 | ~v_59;
assign x_28484 = v_1146 | ~v_58;
assign x_28485 = v_1146 | ~v_56;
assign x_28486 = v_1146 | ~v_54;
assign x_28487 = ~v_75 | v_153 | v_1145;
assign x_28488 = ~v_90 | ~v_153 | v_1144;
assign x_28489 = ~v_4 | ~v_152 | v_1143;
assign x_28490 = ~v_2 | v_152 | v_1142;
assign x_28491 = v_1141 | ~v_743;
assign x_28492 = v_1141 | ~v_744;
assign x_28493 = v_1141 | ~v_745;
assign x_28494 = v_1141 | ~v_746;
assign x_28495 = v_1141 | ~v_935;
assign x_28496 = v_1141 | ~v_936;
assign x_28497 = v_1141 | ~v_937;
assign x_28498 = v_1141 | ~v_938;
assign x_28499 = v_1141 | ~v_751;
assign x_28500 = v_1141 | ~v_752;
assign x_28501 = v_1141 | ~v_753;
assign x_28502 = v_1141 | ~v_754;
assign x_28503 = v_1141 | ~v_755;
assign x_28504 = v_1141 | ~v_756;
assign x_28505 = v_1141 | ~v_939;
assign x_28506 = v_1141 | ~v_940;
assign x_28507 = v_1141 | ~v_941;
assign x_28508 = v_1141 | ~v_942;
assign x_28509 = v_1141 | ~v_761;
assign x_28510 = v_1141 | ~v_762;
assign x_28511 = v_1141 | ~v_763;
assign x_28512 = v_1141 | ~v_764;
assign x_28513 = v_1141 | ~v_765;
assign x_28514 = v_1141 | ~v_766;
assign x_28515 = v_1141 | ~v_1137;
assign x_28516 = v_1141 | ~v_1138;
assign x_28517 = v_1141 | ~v_945;
assign x_28518 = v_1141 | ~v_946;
assign x_28519 = v_1141 | ~v_773;
assign x_28520 = v_1141 | ~v_774;
assign x_28521 = v_1141 | ~v_1139;
assign x_28522 = v_1141 | ~v_1140;
assign x_28523 = v_1141 | ~v_182;
assign x_28524 = v_1141 | ~v_162;
assign x_28525 = v_1141 | ~v_161;
assign x_28526 = v_1141 | ~v_137;
assign x_28527 = v_1141 | ~v_136;
assign x_28528 = v_1141 | ~v_134;
assign x_28529 = v_1141 | ~v_18;
assign x_28530 = v_1141 | ~v_17;
assign x_28531 = v_1141 | ~v_16;
assign x_28532 = v_1141 | ~v_15;
assign x_28533 = v_1141 | ~v_13;
assign x_28534 = v_1141 | ~v_11;
assign x_28535 = ~v_33 | v_153 | v_1140;
assign x_28536 = ~v_48 | ~v_153 | v_1139;
assign x_28537 = ~v_5 | ~v_152 | v_1138;
assign x_28538 = ~v_1 | v_152 | v_1137;
assign x_28539 = ~v_1135 | ~v_1130 | ~v_1125 | v_1136;
assign x_28540 = v_1135 | ~v_809;
assign x_28541 = v_1135 | ~v_810;
assign x_28542 = v_1135 | ~v_811;
assign x_28543 = v_1135 | ~v_812;
assign x_28544 = v_1135 | ~v_1073;
assign x_28545 = v_1135 | ~v_1074;
assign x_28546 = v_1135 | ~v_1075;
assign x_28547 = v_1135 | ~v_1076;
assign x_28548 = v_1135 | ~v_817;
assign x_28549 = v_1135 | ~v_1011;
assign x_28550 = v_1135 | ~v_1012;
assign x_28551 = v_1135 | ~v_820;
assign x_28552 = v_1135 | ~v_1013;
assign x_28553 = v_1135 | ~v_1014;
assign x_28554 = v_1135 | ~v_1077;
assign x_28555 = v_1135 | ~v_1078;
assign x_28556 = v_1135 | ~v_1079;
assign x_28557 = v_1135 | ~v_1080;
assign x_28558 = v_1135 | ~v_827;
assign x_28559 = v_1135 | ~v_1015;
assign x_28560 = v_1135 | ~v_1016;
assign x_28561 = v_1135 | ~v_830;
assign x_28562 = v_1135 | ~v_1017;
assign x_28563 = v_1135 | ~v_1018;
assign x_28564 = v_1135 | ~v_1085;
assign x_28565 = v_1135 | ~v_1131;
assign x_28566 = v_1135 | ~v_1132;
assign x_28567 = v_1135 | ~v_1086;
assign x_28568 = v_1135 | ~v_1133;
assign x_28569 = v_1135 | ~v_1134;
assign x_28570 = v_1135 | ~v_1023;
assign x_28571 = v_1135 | ~v_1024;
assign x_28572 = v_1135 | ~v_184;
assign x_28573 = v_1135 | ~v_172;
assign x_28574 = v_1135 | ~v_171;
assign x_28575 = v_1135 | ~v_170;
assign x_28576 = v_1135 | ~v_169;
assign x_28577 = v_1135 | ~v_149;
assign x_28578 = v_1135 | ~v_148;
assign x_28579 = v_1135 | ~v_147;
assign x_28580 = v_1135 | ~v_102;
assign x_28581 = v_1135 | ~v_101;
assign x_28582 = v_1135 | ~v_100;
assign x_28583 = v_1135 | ~v_99;
assign x_28584 = ~v_132 | ~v_139 | v_1134;
assign x_28585 = ~v_6 | ~v_140 | v_1133;
assign x_28586 = ~v_117 | v_139 | v_1132;
assign x_28587 = ~v_3 | v_140 | v_1131;
assign x_28588 = v_1130 | ~v_776;
assign x_28589 = v_1130 | ~v_777;
assign x_28590 = v_1130 | ~v_778;
assign x_28591 = v_1130 | ~v_779;
assign x_28592 = v_1130 | ~v_1058;
assign x_28593 = v_1130 | ~v_1059;
assign x_28594 = v_1130 | ~v_1060;
assign x_28595 = v_1130 | ~v_1061;
assign x_28596 = v_1130 | ~v_784;
assign x_28597 = v_1130 | ~v_996;
assign x_28598 = v_1130 | ~v_997;
assign x_28599 = v_1130 | ~v_787;
assign x_28600 = v_1130 | ~v_998;
assign x_28601 = v_1130 | ~v_999;
assign x_28602 = v_1130 | ~v_1062;
assign x_28603 = v_1130 | ~v_1063;
assign x_28604 = v_1130 | ~v_1064;
assign x_28605 = v_1130 | ~v_1065;
assign x_28606 = v_1130 | ~v_794;
assign x_28607 = v_1130 | ~v_1000;
assign x_28608 = v_1130 | ~v_1001;
assign x_28609 = v_1130 | ~v_797;
assign x_28610 = v_1130 | ~v_1002;
assign x_28611 = v_1130 | ~v_1003;
assign x_28612 = v_1130 | ~v_1070;
assign x_28613 = v_1130 | ~v_1126;
assign x_28614 = v_1130 | ~v_1127;
assign x_28615 = v_1130 | ~v_1071;
assign x_28616 = v_1130 | ~v_1128;
assign x_28617 = v_1130 | ~v_1129;
assign x_28618 = v_1130 | ~v_1008;
assign x_28619 = v_1130 | ~v_1009;
assign x_28620 = v_1130 | ~v_183;
assign x_28621 = v_1130 | ~v_168;
assign x_28622 = v_1130 | ~v_167;
assign x_28623 = v_1130 | ~v_166;
assign x_28624 = v_1130 | ~v_165;
assign x_28625 = v_1130 | ~v_144;
assign x_28626 = v_1130 | ~v_143;
assign x_28627 = v_1130 | ~v_142;
assign x_28628 = v_1130 | ~v_60;
assign x_28629 = v_1130 | ~v_59;
assign x_28630 = v_1130 | ~v_58;
assign x_28631 = v_1130 | ~v_57;
assign x_28632 = ~v_90 | ~v_139 | v_1129;
assign x_28633 = ~v_4 | ~v_140 | v_1128;
assign x_28634 = ~v_75 | v_139 | v_1127;
assign x_28635 = ~v_2 | v_140 | v_1126;
assign x_28636 = v_1125 | ~v_743;
assign x_28637 = v_1125 | ~v_744;
assign x_28638 = v_1125 | ~v_745;
assign x_28639 = v_1125 | ~v_746;
assign x_28640 = v_1125 | ~v_1043;
assign x_28641 = v_1125 | ~v_1044;
assign x_28642 = v_1125 | ~v_1045;
assign x_28643 = v_1125 | ~v_1046;
assign x_28644 = v_1125 | ~v_751;
assign x_28645 = v_1125 | ~v_981;
assign x_28646 = v_1125 | ~v_982;
assign x_28647 = v_1125 | ~v_754;
assign x_28648 = v_1125 | ~v_983;
assign x_28649 = v_1125 | ~v_984;
assign x_28650 = v_1125 | ~v_1047;
assign x_28651 = v_1125 | ~v_1048;
assign x_28652 = v_1125 | ~v_1049;
assign x_28653 = v_1125 | ~v_1050;
assign x_28654 = v_1125 | ~v_761;
assign x_28655 = v_1125 | ~v_985;
assign x_28656 = v_1125 | ~v_986;
assign x_28657 = v_1125 | ~v_764;
assign x_28658 = v_1125 | ~v_987;
assign x_28659 = v_1125 | ~v_988;
assign x_28660 = v_1125 | ~v_1055;
assign x_28661 = v_1125 | ~v_1121;
assign x_28662 = v_1125 | ~v_1122;
assign x_28663 = v_1125 | ~v_1056;
assign x_28664 = v_1125 | ~v_1123;
assign x_28665 = v_1125 | ~v_1124;
assign x_28666 = v_1125 | ~v_182;
assign x_28667 = v_1125 | ~v_164;
assign x_28668 = v_1125 | ~v_163;
assign x_28669 = v_1125 | ~v_162;
assign x_28670 = v_1125 | ~v_161;
assign x_28671 = v_1125 | ~v_136;
assign x_28672 = v_1125 | ~v_135;
assign x_28673 = v_1125 | ~v_134;
assign x_28674 = v_1125 | ~v_993;
assign x_28675 = v_1125 | ~v_994;
assign x_28676 = v_1125 | ~v_17;
assign x_28677 = v_1125 | ~v_16;
assign x_28678 = v_1125 | ~v_15;
assign x_28679 = v_1125 | ~v_14;
assign x_28680 = ~v_48 | ~v_139 | v_1124;
assign x_28681 = ~v_5 | ~v_140 | v_1123;
assign x_28682 = ~v_33 | v_139 | v_1122;
assign x_28683 = ~v_1 | v_140 | v_1121;
assign x_28684 = ~v_1119 | ~v_1114 | ~v_1109 | v_1120;
assign x_28685 = v_1119 | ~v_809;
assign x_28686 = v_1119 | ~v_810;
assign x_28687 = v_1119 | ~v_811;
assign x_28688 = v_1119 | ~v_812;
assign x_28689 = v_1119 | ~v_1073;
assign x_28690 = v_1119 | ~v_1074;
assign x_28691 = v_1119 | ~v_1075;
assign x_28692 = v_1119 | ~v_1076;
assign x_28693 = v_1119 | ~v_965;
assign x_28694 = v_1119 | ~v_966;
assign x_28695 = v_1119 | ~v_967;
assign x_28696 = v_1119 | ~v_968;
assign x_28697 = v_1119 | ~v_817;
assign x_28698 = v_1119 | ~v_820;
assign x_28699 = v_1119 | ~v_1077;
assign x_28700 = v_1119 | ~v_1078;
assign x_28701 = v_1119 | ~v_1079;
assign x_28702 = v_1119 | ~v_1080;
assign x_28703 = v_1119 | ~v_969;
assign x_28704 = v_1119 | ~v_970;
assign x_28705 = v_1119 | ~v_971;
assign x_28706 = v_1119 | ~v_972;
assign x_28707 = v_1119 | ~v_827;
assign x_28708 = v_1119 | ~v_830;
assign x_28709 = v_1119 | ~v_975;
assign x_28710 = v_1119 | ~v_976;
assign x_28711 = v_1119 | ~v_1115;
assign x_28712 = v_1119 | ~v_1116;
assign x_28713 = v_1119 | ~v_1085;
assign x_28714 = v_1119 | ~v_1086;
assign x_28715 = v_1119 | ~v_1117;
assign x_28716 = v_1119 | ~v_1118;
assign x_28717 = v_1119 | ~v_184;
assign x_28718 = v_1119 | ~v_171;
assign x_28719 = v_1119 | ~v_170;
assign x_28720 = v_1119 | ~v_169;
assign x_28721 = v_1119 | ~v_151;
assign x_28722 = v_1119 | ~v_150;
assign x_28723 = v_1119 | ~v_149;
assign x_28724 = v_1119 | ~v_147;
assign x_28725 = v_1119 | ~v_103;
assign x_28726 = v_1119 | ~v_101;
assign x_28727 = v_1119 | ~v_100;
assign x_28728 = v_1119 | ~v_96;
assign x_28729 = ~v_132 | ~v_174 | v_1118;
assign x_28730 = ~v_117 | v_174 | v_1117;
assign x_28731 = ~v_6 | ~v_173 | v_1116;
assign x_28732 = ~v_3 | v_173 | v_1115;
assign x_28733 = v_1114 | ~v_776;
assign x_28734 = v_1114 | ~v_777;
assign x_28735 = v_1114 | ~v_778;
assign x_28736 = v_1114 | ~v_779;
assign x_28737 = v_1114 | ~v_1058;
assign x_28738 = v_1114 | ~v_1059;
assign x_28739 = v_1114 | ~v_1060;
assign x_28740 = v_1114 | ~v_1061;
assign x_28741 = v_1114 | ~v_950;
assign x_28742 = v_1114 | ~v_951;
assign x_28743 = v_1114 | ~v_952;
assign x_28744 = v_1114 | ~v_953;
assign x_28745 = v_1114 | ~v_784;
assign x_28746 = v_1114 | ~v_787;
assign x_28747 = v_1114 | ~v_1062;
assign x_28748 = v_1114 | ~v_1063;
assign x_28749 = v_1114 | ~v_1064;
assign x_28750 = v_1114 | ~v_1065;
assign x_28751 = v_1114 | ~v_954;
assign x_28752 = v_1114 | ~v_955;
assign x_28753 = v_1114 | ~v_956;
assign x_28754 = v_1114 | ~v_957;
assign x_28755 = v_1114 | ~v_794;
assign x_28756 = v_1114 | ~v_797;
assign x_28757 = v_1114 | ~v_960;
assign x_28758 = v_1114 | ~v_961;
assign x_28759 = v_1114 | ~v_1110;
assign x_28760 = v_1114 | ~v_1111;
assign x_28761 = v_1114 | ~v_1070;
assign x_28762 = v_1114 | ~v_1071;
assign x_28763 = v_1114 | ~v_1112;
assign x_28764 = v_1114 | ~v_1113;
assign x_28765 = v_1114 | ~v_183;
assign x_28766 = v_1114 | ~v_167;
assign x_28767 = v_1114 | ~v_166;
assign x_28768 = v_1114 | ~v_165;
assign x_28769 = v_1114 | ~v_146;
assign x_28770 = v_1114 | ~v_145;
assign x_28771 = v_1114 | ~v_144;
assign x_28772 = v_1114 | ~v_142;
assign x_28773 = v_1114 | ~v_61;
assign x_28774 = v_1114 | ~v_59;
assign x_28775 = v_1114 | ~v_58;
assign x_28776 = v_1114 | ~v_54;
assign x_28777 = ~v_90 | ~v_174 | v_1113;
assign x_28778 = ~v_75 | v_174 | v_1112;
assign x_28779 = ~v_4 | ~v_173 | v_1111;
assign x_28780 = ~v_2 | v_173 | v_1110;
assign x_28781 = v_1109 | ~v_743;
assign x_28782 = v_1109 | ~v_744;
assign x_28783 = v_1109 | ~v_745;
assign x_28784 = v_1109 | ~v_746;
assign x_28785 = v_1109 | ~v_1043;
assign x_28786 = v_1109 | ~v_1044;
assign x_28787 = v_1109 | ~v_1045;
assign x_28788 = v_1109 | ~v_1046;
assign x_28789 = v_1109 | ~v_935;
assign x_28790 = v_1109 | ~v_936;
assign x_28791 = v_1109 | ~v_937;
assign x_28792 = v_1109 | ~v_938;
assign x_28793 = v_1109 | ~v_751;
assign x_28794 = v_1109 | ~v_754;
assign x_28795 = v_1109 | ~v_1047;
assign x_28796 = v_1109 | ~v_1048;
assign x_28797 = v_1109 | ~v_1049;
assign x_28798 = v_1109 | ~v_1050;
assign x_28799 = v_1109 | ~v_939;
assign x_28800 = v_1109 | ~v_940;
assign x_28801 = v_1109 | ~v_941;
assign x_28802 = v_1109 | ~v_942;
assign x_28803 = v_1109 | ~v_761;
assign x_28804 = v_1109 | ~v_764;
assign x_28805 = v_1109 | ~v_945;
assign x_28806 = v_1109 | ~v_946;
assign x_28807 = v_1109 | ~v_1105;
assign x_28808 = v_1109 | ~v_1106;
assign x_28809 = v_1109 | ~v_1055;
assign x_28810 = v_1109 | ~v_1056;
assign x_28811 = v_1109 | ~v_1107;
assign x_28812 = v_1109 | ~v_1108;
assign x_28813 = v_1109 | ~v_182;
assign x_28814 = v_1109 | ~v_163;
assign x_28815 = v_1109 | ~v_162;
assign x_28816 = v_1109 | ~v_161;
assign x_28817 = v_1109 | ~v_138;
assign x_28818 = v_1109 | ~v_137;
assign x_28819 = v_1109 | ~v_136;
assign x_28820 = v_1109 | ~v_134;
assign x_28821 = v_1109 | ~v_18;
assign x_28822 = v_1109 | ~v_16;
assign x_28823 = v_1109 | ~v_15;
assign x_28824 = v_1109 | ~v_11;
assign x_28825 = ~v_48 | ~v_174 | v_1108;
assign x_28826 = ~v_33 | v_174 | v_1107;
assign x_28827 = ~v_5 | ~v_173 | v_1106;
assign x_28828 = ~v_1 | v_173 | v_1105;
assign x_28829 = ~v_1103 | ~v_1098 | ~v_1093 | v_1104;
assign x_28830 = v_1103 | ~v_809;
assign x_28831 = v_1103 | ~v_810;
assign x_28832 = v_1103 | ~v_811;
assign x_28833 = v_1103 | ~v_812;
assign x_28834 = v_1103 | ~v_1073;
assign x_28835 = v_1103 | ~v_1074;
assign x_28836 = v_1103 | ~v_1075;
assign x_28837 = v_1103 | ~v_1076;
assign x_28838 = v_1103 | ~v_919;
assign x_28839 = v_1103 | ~v_920;
assign x_28840 = v_1103 | ~v_817;
assign x_28841 = v_1103 | ~v_820;
assign x_28842 = v_1103 | ~v_1077;
assign x_28843 = v_1103 | ~v_1078;
assign x_28844 = v_1103 | ~v_1079;
assign x_28845 = v_1103 | ~v_1080;
assign x_28846 = v_1103 | ~v_921;
assign x_28847 = v_1103 | ~v_922;
assign x_28848 = v_1103 | ~v_923;
assign x_28849 = v_1103 | ~v_924;
assign x_28850 = v_1103 | ~v_827;
assign x_28851 = v_1103 | ~v_830;
assign x_28852 = v_1103 | ~v_927;
assign x_28853 = v_1103 | ~v_928;
assign x_28854 = v_1103 | ~v_1099;
assign x_28855 = v_1103 | ~v_1100;
assign x_28856 = v_1103 | ~v_1101;
assign x_28857 = v_1103 | ~v_1102;
assign x_28858 = v_1103 | ~v_1085;
assign x_28859 = v_1103 | ~v_1086;
assign x_28860 = v_1103 | ~v_931;
assign x_28861 = v_1103 | ~v_932;
assign x_28862 = v_1103 | ~v_184;
assign x_28863 = v_1103 | ~v_171;
assign x_28864 = v_1103 | ~v_170;
assign x_28865 = v_1103 | ~v_169;
assign x_28866 = v_1103 | ~v_150;
assign x_28867 = v_1103 | ~v_149;
assign x_28868 = v_1103 | ~v_148;
assign x_28869 = v_1103 | ~v_103;
assign x_28870 = v_1103 | ~v_102;
assign x_28871 = v_1103 | ~v_101;
assign x_28872 = v_1103 | ~v_100;
assign x_28873 = v_1103 | ~v_95;
assign x_28874 = ~v_132 | ~v_141 | v_1102;
assign x_28875 = ~v_6 | ~v_141 | v_1101;
assign x_28876 = ~v_117 | v_141 | v_1100;
assign x_28877 = ~v_3 | v_141 | v_1099;
assign x_28878 = v_1098 | ~v_776;
assign x_28879 = v_1098 | ~v_777;
assign x_28880 = v_1098 | ~v_778;
assign x_28881 = v_1098 | ~v_779;
assign x_28882 = v_1098 | ~v_1058;
assign x_28883 = v_1098 | ~v_1059;
assign x_28884 = v_1098 | ~v_1060;
assign x_28885 = v_1098 | ~v_1061;
assign x_28886 = v_1098 | ~v_904;
assign x_28887 = v_1098 | ~v_905;
assign x_28888 = v_1098 | ~v_784;
assign x_28889 = v_1098 | ~v_787;
assign x_28890 = v_1098 | ~v_1062;
assign x_28891 = v_1098 | ~v_1063;
assign x_28892 = v_1098 | ~v_1064;
assign x_28893 = v_1098 | ~v_1065;
assign x_28894 = v_1098 | ~v_906;
assign x_28895 = v_1098 | ~v_907;
assign x_28896 = v_1098 | ~v_908;
assign x_28897 = v_1098 | ~v_909;
assign x_28898 = v_1098 | ~v_794;
assign x_28899 = v_1098 | ~v_797;
assign x_28900 = v_1098 | ~v_912;
assign x_28901 = v_1098 | ~v_913;
assign x_28902 = v_1098 | ~v_1094;
assign x_28903 = v_1098 | ~v_1095;
assign x_28904 = v_1098 | ~v_1096;
assign x_28905 = v_1098 | ~v_1097;
assign x_28906 = v_1098 | ~v_1070;
assign x_28907 = v_1098 | ~v_1071;
assign x_28908 = v_1098 | ~v_916;
assign x_28909 = v_1098 | ~v_917;
assign x_28910 = v_1098 | ~v_183;
assign x_28911 = v_1098 | ~v_167;
assign x_28912 = v_1098 | ~v_166;
assign x_28913 = v_1098 | ~v_165;
assign x_28914 = v_1098 | ~v_145;
assign x_28915 = v_1098 | ~v_144;
assign x_28916 = v_1098 | ~v_143;
assign x_28917 = v_1098 | ~v_61;
assign x_28918 = v_1098 | ~v_60;
assign x_28919 = v_1098 | ~v_59;
assign x_28920 = v_1098 | ~v_58;
assign x_28921 = v_1098 | ~v_53;
assign x_28922 = ~v_90 | ~v_141 | v_1097;
assign x_28923 = ~v_4 | ~v_141 | v_1096;
assign x_28924 = ~v_75 | v_141 | v_1095;
assign x_28925 = ~v_2 | v_141 | v_1094;
assign x_28926 = v_1093 | ~v_743;
assign x_28927 = v_1093 | ~v_744;
assign x_28928 = v_1093 | ~v_745;
assign x_28929 = v_1093 | ~v_746;
assign x_28930 = v_1093 | ~v_1043;
assign x_28931 = v_1093 | ~v_1044;
assign x_28932 = v_1093 | ~v_1045;
assign x_28933 = v_1093 | ~v_1046;
assign x_28934 = v_1093 | ~v_889;
assign x_28935 = v_1093 | ~v_890;
assign x_28936 = v_1093 | ~v_751;
assign x_28937 = v_1093 | ~v_754;
assign x_28938 = v_1093 | ~v_1047;
assign x_28939 = v_1093 | ~v_1048;
assign x_28940 = v_1093 | ~v_1049;
assign x_28941 = v_1093 | ~v_1050;
assign x_28942 = v_1093 | ~v_891;
assign x_28943 = v_1093 | ~v_892;
assign x_28944 = v_1093 | ~v_893;
assign x_28945 = v_1093 | ~v_894;
assign x_28946 = v_1093 | ~v_761;
assign x_28947 = v_1093 | ~v_764;
assign x_28948 = v_1093 | ~v_897;
assign x_28949 = v_1093 | ~v_898;
assign x_28950 = v_1093 | ~v_1089;
assign x_28951 = v_1093 | ~v_1090;
assign x_28952 = v_1093 | ~v_1091;
assign x_28953 = v_1093 | ~v_1092;
assign x_28954 = v_1093 | ~v_1055;
assign x_28955 = v_1093 | ~v_1056;
assign x_28956 = v_1093 | ~v_901;
assign x_28957 = v_1093 | ~v_902;
assign x_28958 = v_1093 | ~v_182;
assign x_28959 = v_1093 | ~v_163;
assign x_28960 = v_1093 | ~v_162;
assign x_28961 = v_1093 | ~v_161;
assign x_28962 = v_1093 | ~v_137;
assign x_28963 = v_1093 | ~v_136;
assign x_28964 = v_1093 | ~v_135;
assign x_28965 = v_1093 | ~v_18;
assign x_28966 = v_1093 | ~v_17;
assign x_28967 = v_1093 | ~v_16;
assign x_28968 = v_1093 | ~v_15;
assign x_28969 = v_1093 | ~v_10;
assign x_28970 = ~v_48 | ~v_141 | v_1092;
assign x_28971 = ~v_5 | ~v_141 | v_1091;
assign x_28972 = ~v_33 | v_141 | v_1090;
assign x_28973 = ~v_1 | v_141 | v_1089;
assign x_28974 = ~v_1087 | ~v_1072 | ~v_1057 | v_1088;
assign x_28975 = v_1087 | ~v_809;
assign x_28976 = v_1087 | ~v_810;
assign x_28977 = v_1087 | ~v_811;
assign x_28978 = v_1087 | ~v_812;
assign x_28979 = v_1087 | ~v_1073;
assign x_28980 = v_1087 | ~v_1074;
assign x_28981 = v_1087 | ~v_1075;
assign x_28982 = v_1087 | ~v_1076;
assign x_28983 = v_1087 | ~v_813;
assign x_28984 = v_1087 | ~v_814;
assign x_28985 = v_1087 | ~v_815;
assign x_28986 = v_1087 | ~v_816;
assign x_28987 = v_1087 | ~v_817;
assign x_28988 = v_1087 | ~v_820;
assign x_28989 = v_1087 | ~v_1077;
assign x_28990 = v_1087 | ~v_1078;
assign x_28991 = v_1087 | ~v_1079;
assign x_28992 = v_1087 | ~v_1080;
assign x_28993 = v_1087 | ~v_823;
assign x_28994 = v_1087 | ~v_824;
assign x_28995 = v_1087 | ~v_825;
assign x_28996 = v_1087 | ~v_826;
assign x_28997 = v_1087 | ~v_827;
assign x_28998 = v_1087 | ~v_830;
assign x_28999 = v_1087 | ~v_837;
assign x_29000 = v_1087 | ~v_838;
assign x_29001 = v_1087 | ~v_1081;
assign x_29002 = v_1087 | ~v_1082;
assign x_29003 = v_1087 | ~v_1083;
assign x_29004 = v_1087 | ~v_1084;
assign x_29005 = v_1087 | ~v_1085;
assign x_29006 = v_1087 | ~v_1086;
assign x_29007 = v_1087 | ~v_184;
assign x_29008 = v_1087 | ~v_171;
assign x_29009 = v_1087 | ~v_170;
assign x_29010 = v_1087 | ~v_169;
assign x_29011 = v_1087 | ~v_160;
assign x_29012 = v_1087 | ~v_150;
assign x_29013 = v_1087 | ~v_148;
assign x_29014 = v_1087 | ~v_147;
assign x_29015 = v_1087 | ~v_103;
assign x_29016 = v_1087 | ~v_102;
assign x_29017 = v_1087 | ~v_100;
assign x_29018 = v_1087 | ~v_97;
assign x_29019 = ~v_129 | ~v_141 | v_1086;
assign x_29020 = ~v_114 | v_141 | v_1085;
assign x_29021 = ~v_132 | ~v_176 | v_1084;
assign x_29022 = ~v_6 | ~v_175 | v_1083;
assign x_29023 = ~v_117 | v_176 | v_1082;
assign x_29024 = ~v_3 | v_175 | v_1081;
assign x_29025 = ~v_127 | ~v_173 | v_1080;
assign x_29026 = ~v_121 | ~v_174 | v_1079;
assign x_29027 = ~v_112 | v_173 | v_1078;
assign x_29028 = ~v_106 | v_174 | v_1077;
assign x_29029 = ~v_128 | ~v_175 | v_1076;
assign x_29030 = ~v_125 | ~v_176 | v_1075;
assign x_29031 = ~v_113 | v_175 | v_1074;
assign x_29032 = ~v_110 | v_176 | v_1073;
assign x_29033 = v_1072 | ~v_776;
assign x_29034 = v_1072 | ~v_777;
assign x_29035 = v_1072 | ~v_778;
assign x_29036 = v_1072 | ~v_779;
assign x_29037 = v_1072 | ~v_1058;
assign x_29038 = v_1072 | ~v_1059;
assign x_29039 = v_1072 | ~v_1060;
assign x_29040 = v_1072 | ~v_1061;
assign x_29041 = v_1072 | ~v_780;
assign x_29042 = v_1072 | ~v_781;
assign x_29043 = v_1072 | ~v_782;
assign x_29044 = v_1072 | ~v_783;
assign x_29045 = v_1072 | ~v_784;
assign x_29046 = v_1072 | ~v_787;
assign x_29047 = v_1072 | ~v_1062;
assign x_29048 = v_1072 | ~v_1063;
assign x_29049 = v_1072 | ~v_1064;
assign x_29050 = v_1072 | ~v_1065;
assign x_29051 = v_1072 | ~v_790;
assign x_29052 = v_1072 | ~v_791;
assign x_29053 = v_1072 | ~v_792;
assign x_29054 = v_1072 | ~v_793;
assign x_29055 = v_1072 | ~v_794;
assign x_29056 = v_1072 | ~v_797;
assign x_29057 = v_1072 | ~v_804;
assign x_29058 = v_1072 | ~v_805;
assign x_29059 = v_1072 | ~v_1066;
assign x_29060 = v_1072 | ~v_1067;
assign x_29061 = v_1072 | ~v_1068;
assign x_29062 = v_1072 | ~v_1069;
assign x_29063 = v_1072 | ~v_1070;
assign x_29064 = v_1072 | ~v_1071;
assign x_29065 = v_1072 | ~v_183;
assign x_29066 = v_1072 | ~v_167;
assign x_29067 = v_1072 | ~v_166;
assign x_29068 = v_1072 | ~v_165;
assign x_29069 = v_1072 | ~v_159;
assign x_29070 = v_1072 | ~v_145;
assign x_29071 = v_1072 | ~v_143;
assign x_29072 = v_1072 | ~v_142;
assign x_29073 = v_1072 | ~v_61;
assign x_29074 = v_1072 | ~v_60;
assign x_29075 = v_1072 | ~v_58;
assign x_29076 = v_1072 | ~v_55;
assign x_29077 = ~v_87 | ~v_141 | v_1071;
assign x_29078 = ~v_72 | v_141 | v_1070;
assign x_29079 = ~v_90 | ~v_176 | v_1069;
assign x_29080 = ~v_4 | ~v_175 | v_1068;
assign x_29081 = ~v_75 | v_176 | v_1067;
assign x_29082 = ~v_2 | v_175 | v_1066;
assign x_29083 = ~v_85 | ~v_173 | v_1065;
assign x_29084 = ~v_79 | ~v_174 | v_1064;
assign x_29085 = ~v_70 | v_173 | v_1063;
assign x_29086 = ~v_64 | v_174 | v_1062;
assign x_29087 = ~v_86 | ~v_175 | v_1061;
assign x_29088 = ~v_83 | ~v_176 | v_1060;
assign x_29089 = ~v_71 | v_175 | v_1059;
assign x_29090 = ~v_68 | v_176 | v_1058;
assign x_29091 = v_1057 | ~v_743;
assign x_29092 = v_1057 | ~v_744;
assign x_29093 = v_1057 | ~v_745;
assign x_29094 = v_1057 | ~v_746;
assign x_29095 = v_1057 | ~v_1043;
assign x_29096 = v_1057 | ~v_1044;
assign x_29097 = v_1057 | ~v_1045;
assign x_29098 = v_1057 | ~v_1046;
assign x_29099 = v_1057 | ~v_747;
assign x_29100 = v_1057 | ~v_748;
assign x_29101 = v_1057 | ~v_749;
assign x_29102 = v_1057 | ~v_750;
assign x_29103 = v_1057 | ~v_751;
assign x_29104 = v_1057 | ~v_754;
assign x_29105 = v_1057 | ~v_1047;
assign x_29106 = v_1057 | ~v_1048;
assign x_29107 = v_1057 | ~v_1049;
assign x_29108 = v_1057 | ~v_1050;
assign x_29109 = v_1057 | ~v_757;
assign x_29110 = v_1057 | ~v_758;
assign x_29111 = v_1057 | ~v_759;
assign x_29112 = v_1057 | ~v_760;
assign x_29113 = v_1057 | ~v_761;
assign x_29114 = v_1057 | ~v_764;
assign x_29115 = v_1057 | ~v_771;
assign x_29116 = v_1057 | ~v_772;
assign x_29117 = v_1057 | ~v_1051;
assign x_29118 = v_1057 | ~v_1052;
assign x_29119 = v_1057 | ~v_1053;
assign x_29120 = v_1057 | ~v_1054;
assign x_29121 = v_1057 | ~v_1055;
assign x_29122 = v_1057 | ~v_1056;
assign x_29123 = v_1057 | ~v_182;
assign x_29124 = v_1057 | ~v_163;
assign x_29125 = v_1057 | ~v_162;
assign x_29126 = v_1057 | ~v_161;
assign x_29127 = v_1057 | ~v_155;
assign x_29128 = v_1057 | ~v_137;
assign x_29129 = v_1057 | ~v_135;
assign x_29130 = v_1057 | ~v_134;
assign x_29131 = v_1057 | ~v_18;
assign x_29132 = v_1057 | ~v_17;
assign x_29133 = v_1057 | ~v_15;
assign x_29134 = v_1057 | ~v_12;
assign x_29135 = ~v_45 | ~v_141 | v_1056;
assign x_29136 = ~v_30 | v_141 | v_1055;
assign x_29137 = ~v_48 | ~v_176 | v_1054;
assign x_29138 = ~v_5 | ~v_175 | v_1053;
assign x_29139 = ~v_33 | v_176 | v_1052;
assign x_29140 = ~v_1 | v_175 | v_1051;
assign x_29141 = ~v_43 | ~v_173 | v_1050;
assign x_29142 = ~v_37 | ~v_174 | v_1049;
assign x_29143 = ~v_28 | v_173 | v_1048;
assign x_29144 = ~v_22 | v_174 | v_1047;
assign x_29145 = ~v_44 | ~v_175 | v_1046;
assign x_29146 = ~v_41 | ~v_176 | v_1045;
assign x_29147 = ~v_29 | v_175 | v_1044;
assign x_29148 = ~v_26 | v_176 | v_1043;
assign x_29149 = ~v_1041 | ~v_1036 | ~v_1031 | v_1042;
assign x_29150 = v_1041 | ~v_809;
assign x_29151 = v_1041 | ~v_810;
assign x_29152 = v_1041 | ~v_811;
assign x_29153 = v_1041 | ~v_812;
assign x_29154 = v_1041 | ~v_919;
assign x_29155 = v_1041 | ~v_920;
assign x_29156 = v_1041 | ~v_817;
assign x_29157 = v_1041 | ~v_818;
assign x_29158 = v_1041 | ~v_819;
assign x_29159 = v_1041 | ~v_820;
assign x_29160 = v_1041 | ~v_821;
assign x_29161 = v_1041 | ~v_822;
assign x_29162 = v_1041 | ~v_921;
assign x_29163 = v_1041 | ~v_922;
assign x_29164 = v_1041 | ~v_923;
assign x_29165 = v_1041 | ~v_924;
assign x_29166 = v_1041 | ~v_827;
assign x_29167 = v_1041 | ~v_828;
assign x_29168 = v_1041 | ~v_829;
assign x_29169 = v_1041 | ~v_830;
assign x_29170 = v_1041 | ~v_831;
assign x_29171 = v_1041 | ~v_832;
assign x_29172 = v_1041 | ~v_1037;
assign x_29173 = v_1041 | ~v_1038;
assign x_29174 = v_1041 | ~v_1039;
assign x_29175 = v_1041 | ~v_1040;
assign x_29176 = v_1041 | ~v_927;
assign x_29177 = v_1041 | ~v_928;
assign x_29178 = v_1041 | ~v_839;
assign x_29179 = v_1041 | ~v_840;
assign x_29180 = v_1041 | ~v_931;
assign x_29181 = v_1041 | ~v_932;
assign x_29182 = v_1041 | ~v_184;
assign x_29183 = v_1041 | ~v_170;
assign x_29184 = v_1041 | ~v_169;
assign x_29185 = v_1041 | ~v_151;
assign x_29186 = v_1041 | ~v_150;
assign x_29187 = v_1041 | ~v_149;
assign x_29188 = v_1041 | ~v_148;
assign x_29189 = v_1041 | ~v_147;
assign x_29190 = v_1041 | ~v_103;
assign x_29191 = v_1041 | ~v_101;
assign x_29192 = v_1041 | ~v_100;
assign x_29193 = v_1041 | ~v_98;
assign x_29194 = ~v_132 | ~v_140 | v_1040;
assign x_29195 = ~v_6 | ~v_139 | v_1039;
assign x_29196 = ~v_117 | v_140 | v_1038;
assign x_29197 = ~v_3 | v_139 | v_1037;
assign x_29198 = v_1036 | ~v_776;
assign x_29199 = v_1036 | ~v_777;
assign x_29200 = v_1036 | ~v_778;
assign x_29201 = v_1036 | ~v_779;
assign x_29202 = v_1036 | ~v_904;
assign x_29203 = v_1036 | ~v_905;
assign x_29204 = v_1036 | ~v_784;
assign x_29205 = v_1036 | ~v_785;
assign x_29206 = v_1036 | ~v_786;
assign x_29207 = v_1036 | ~v_787;
assign x_29208 = v_1036 | ~v_788;
assign x_29209 = v_1036 | ~v_789;
assign x_29210 = v_1036 | ~v_906;
assign x_29211 = v_1036 | ~v_907;
assign x_29212 = v_1036 | ~v_908;
assign x_29213 = v_1036 | ~v_909;
assign x_29214 = v_1036 | ~v_794;
assign x_29215 = v_1036 | ~v_795;
assign x_29216 = v_1036 | ~v_796;
assign x_29217 = v_1036 | ~v_797;
assign x_29218 = v_1036 | ~v_798;
assign x_29219 = v_1036 | ~v_799;
assign x_29220 = v_1036 | ~v_1032;
assign x_29221 = v_1036 | ~v_1033;
assign x_29222 = v_1036 | ~v_1034;
assign x_29223 = v_1036 | ~v_1035;
assign x_29224 = v_1036 | ~v_912;
assign x_29225 = v_1036 | ~v_913;
assign x_29226 = v_1036 | ~v_806;
assign x_29227 = v_1036 | ~v_807;
assign x_29228 = v_1036 | ~v_916;
assign x_29229 = v_1036 | ~v_917;
assign x_29230 = v_1036 | ~v_183;
assign x_29231 = v_1036 | ~v_166;
assign x_29232 = v_1036 | ~v_165;
assign x_29233 = v_1036 | ~v_146;
assign x_29234 = v_1036 | ~v_145;
assign x_29235 = v_1036 | ~v_144;
assign x_29236 = v_1036 | ~v_143;
assign x_29237 = v_1036 | ~v_142;
assign x_29238 = v_1036 | ~v_61;
assign x_29239 = v_1036 | ~v_59;
assign x_29240 = v_1036 | ~v_58;
assign x_29241 = v_1036 | ~v_56;
assign x_29242 = ~v_90 | ~v_140 | v_1035;
assign x_29243 = ~v_4 | ~v_139 | v_1034;
assign x_29244 = ~v_75 | v_140 | v_1033;
assign x_29245 = ~v_2 | v_139 | v_1032;
assign x_29246 = v_1031 | ~v_743;
assign x_29247 = v_1031 | ~v_744;
assign x_29248 = v_1031 | ~v_745;
assign x_29249 = v_1031 | ~v_746;
assign x_29250 = v_1031 | ~v_889;
assign x_29251 = v_1031 | ~v_890;
assign x_29252 = v_1031 | ~v_751;
assign x_29253 = v_1031 | ~v_752;
assign x_29254 = v_1031 | ~v_753;
assign x_29255 = v_1031 | ~v_754;
assign x_29256 = v_1031 | ~v_755;
assign x_29257 = v_1031 | ~v_756;
assign x_29258 = v_1031 | ~v_891;
assign x_29259 = v_1031 | ~v_892;
assign x_29260 = v_1031 | ~v_893;
assign x_29261 = v_1031 | ~v_894;
assign x_29262 = v_1031 | ~v_761;
assign x_29263 = v_1031 | ~v_762;
assign x_29264 = v_1031 | ~v_763;
assign x_29265 = v_1031 | ~v_764;
assign x_29266 = v_1031 | ~v_765;
assign x_29267 = v_1031 | ~v_766;
assign x_29268 = v_1031 | ~v_1027;
assign x_29269 = v_1031 | ~v_1028;
assign x_29270 = v_1031 | ~v_1029;
assign x_29271 = v_1031 | ~v_1030;
assign x_29272 = v_1031 | ~v_897;
assign x_29273 = v_1031 | ~v_898;
assign x_29274 = v_1031 | ~v_773;
assign x_29275 = v_1031 | ~v_774;
assign x_29276 = v_1031 | ~v_901;
assign x_29277 = v_1031 | ~v_902;
assign x_29278 = v_1031 | ~v_182;
assign x_29279 = v_1031 | ~v_162;
assign x_29280 = v_1031 | ~v_161;
assign x_29281 = v_1031 | ~v_138;
assign x_29282 = v_1031 | ~v_137;
assign x_29283 = v_1031 | ~v_136;
assign x_29284 = v_1031 | ~v_135;
assign x_29285 = v_1031 | ~v_134;
assign x_29286 = v_1031 | ~v_18;
assign x_29287 = v_1031 | ~v_16;
assign x_29288 = v_1031 | ~v_15;
assign x_29289 = v_1031 | ~v_13;
assign x_29290 = ~v_48 | ~v_140 | v_1030;
assign x_29291 = ~v_5 | ~v_139 | v_1029;
assign x_29292 = ~v_33 | v_140 | v_1028;
assign x_29293 = ~v_1 | v_139 | v_1027;
assign x_29294 = ~v_1025 | ~v_1010 | ~v_995 | v_1026;
assign x_29295 = v_1025 | ~v_809;
assign x_29296 = v_1025 | ~v_810;
assign x_29297 = v_1025 | ~v_811;
assign x_29298 = v_1025 | ~v_812;
assign x_29299 = v_1025 | ~v_873;
assign x_29300 = v_1025 | ~v_874;
assign x_29301 = v_1025 | ~v_875;
assign x_29302 = v_1025 | ~v_876;
assign x_29303 = v_1025 | ~v_817;
assign x_29304 = v_1025 | ~v_1011;
assign x_29305 = v_1025 | ~v_1012;
assign x_29306 = v_1025 | ~v_820;
assign x_29307 = v_1025 | ~v_1013;
assign x_29308 = v_1025 | ~v_1014;
assign x_29309 = v_1025 | ~v_877;
assign x_29310 = v_1025 | ~v_878;
assign x_29311 = v_1025 | ~v_879;
assign x_29312 = v_1025 | ~v_880;
assign x_29313 = v_1025 | ~v_827;
assign x_29314 = v_1025 | ~v_1015;
assign x_29315 = v_1025 | ~v_1016;
assign x_29316 = v_1025 | ~v_830;
assign x_29317 = v_1025 | ~v_1017;
assign x_29318 = v_1025 | ~v_1018;
assign x_29319 = v_1025 | ~v_885;
assign x_29320 = v_1025 | ~v_1019;
assign x_29321 = v_1025 | ~v_1020;
assign x_29322 = v_1025 | ~v_886;
assign x_29323 = v_1025 | ~v_1021;
assign x_29324 = v_1025 | ~v_1022;
assign x_29325 = v_1025 | ~v_1023;
assign x_29326 = v_1025 | ~v_1024;
assign x_29327 = v_1025 | ~v_184;
assign x_29328 = v_1025 | ~v_181;
assign x_29329 = v_1025 | ~v_171;
assign x_29330 = v_1025 | ~v_169;
assign x_29331 = v_1025 | ~v_149;
assign x_29332 = v_1025 | ~v_148;
assign x_29333 = v_1025 | ~v_147;
assign x_29334 = v_1025 | ~v_103;
assign x_29335 = v_1025 | ~v_102;
assign x_29336 = v_1025 | ~v_101;
assign x_29337 = v_1025 | ~v_99;
assign x_29338 = v_1025 | ~v_94;
assign x_29339 = ~v_19 | ~v_133 | v_1024;
assign x_29340 = v_19 | ~v_118 | v_1023;
assign x_29341 = ~v_132 | ~v_156 | v_1022;
assign x_29342 = ~v_6 | ~v_157 | v_1021;
assign x_29343 = ~v_117 | v_156 | v_1020;
assign x_29344 = ~v_3 | v_157 | v_1019;
assign x_29345 = ~v_130 | ~v_152 | v_1018;
assign x_29346 = ~v_122 | ~v_153 | v_1017;
assign x_29347 = ~v_115 | v_152 | v_1016;
assign x_29348 = ~v_107 | v_153 | v_1015;
assign x_29349 = ~v_131 | ~v_156 | v_1014;
assign x_29350 = ~v_126 | ~v_157 | v_1013;
assign x_29351 = ~v_116 | v_156 | v_1012;
assign x_29352 = ~v_111 | v_157 | v_1011;
assign x_29353 = v_1010 | ~v_776;
assign x_29354 = v_1010 | ~v_777;
assign x_29355 = v_1010 | ~v_778;
assign x_29356 = v_1010 | ~v_779;
assign x_29357 = v_1010 | ~v_858;
assign x_29358 = v_1010 | ~v_859;
assign x_29359 = v_1010 | ~v_860;
assign x_29360 = v_1010 | ~v_861;
assign x_29361 = v_1010 | ~v_784;
assign x_29362 = v_1010 | ~v_996;
assign x_29363 = v_1010 | ~v_997;
assign x_29364 = v_1010 | ~v_787;
assign x_29365 = v_1010 | ~v_998;
assign x_29366 = v_1010 | ~v_999;
assign x_29367 = v_1010 | ~v_862;
assign x_29368 = v_1010 | ~v_863;
assign x_29369 = v_1010 | ~v_864;
assign x_29370 = v_1010 | ~v_865;
assign x_29371 = v_1010 | ~v_794;
assign x_29372 = v_1010 | ~v_1000;
assign x_29373 = v_1010 | ~v_1001;
assign x_29374 = v_1010 | ~v_797;
assign x_29375 = v_1010 | ~v_1002;
assign x_29376 = v_1010 | ~v_1003;
assign x_29377 = v_1010 | ~v_870;
assign x_29378 = v_1010 | ~v_1004;
assign x_29379 = v_1010 | ~v_1005;
assign x_29380 = v_1010 | ~v_871;
assign x_29381 = v_1010 | ~v_1006;
assign x_29382 = v_1010 | ~v_1007;
assign x_29383 = v_1010 | ~v_1008;
assign x_29384 = v_1010 | ~v_1009;
assign x_29385 = v_1010 | ~v_183;
assign x_29386 = v_1010 | ~v_180;
assign x_29387 = v_1010 | ~v_167;
assign x_29388 = v_1010 | ~v_165;
assign x_29389 = v_1010 | ~v_144;
assign x_29390 = v_1010 | ~v_143;
assign x_29391 = v_1010 | ~v_142;
assign x_29392 = v_1010 | ~v_61;
assign x_29393 = v_1010 | ~v_60;
assign x_29394 = v_1010 | ~v_59;
assign x_29395 = v_1010 | ~v_57;
assign x_29396 = v_1010 | ~v_52;
assign x_29397 = ~v_19 | ~v_91 | v_1009;
assign x_29398 = v_19 | ~v_76 | v_1008;
assign x_29399 = ~v_90 | ~v_156 | v_1007;
assign x_29400 = ~v_4 | ~v_157 | v_1006;
assign x_29401 = ~v_75 | v_156 | v_1005;
assign x_29402 = ~v_2 | v_157 | v_1004;
assign x_29403 = ~v_88 | ~v_152 | v_1003;
assign x_29404 = ~v_80 | ~v_153 | v_1002;
assign x_29405 = ~v_73 | v_152 | v_1001;
assign x_29406 = ~v_65 | v_153 | v_1000;
assign x_29407 = ~v_89 | ~v_156 | v_999;
assign x_29408 = ~v_84 | ~v_157 | v_998;
assign x_29409 = ~v_74 | v_156 | v_997;
assign x_29410 = ~v_69 | v_157 | v_996;
assign x_29411 = v_995 | ~v_743;
assign x_29412 = v_995 | ~v_744;
assign x_29413 = v_995 | ~v_745;
assign x_29414 = v_995 | ~v_746;
assign x_29415 = v_995 | ~v_843;
assign x_29416 = v_995 | ~v_844;
assign x_29417 = v_995 | ~v_845;
assign x_29418 = v_995 | ~v_846;
assign x_29419 = v_995 | ~v_751;
assign x_29420 = v_995 | ~v_981;
assign x_29421 = v_995 | ~v_982;
assign x_29422 = v_995 | ~v_754;
assign x_29423 = v_995 | ~v_983;
assign x_29424 = v_995 | ~v_984;
assign x_29425 = v_995 | ~v_847;
assign x_29426 = v_995 | ~v_848;
assign x_29427 = v_995 | ~v_849;
assign x_29428 = v_995 | ~v_850;
assign x_29429 = v_995 | ~v_761;
assign x_29430 = v_995 | ~v_985;
assign x_29431 = v_995 | ~v_986;
assign x_29432 = v_995 | ~v_764;
assign x_29433 = v_995 | ~v_987;
assign x_29434 = v_995 | ~v_988;
assign x_29435 = v_995 | ~v_855;
assign x_29436 = v_995 | ~v_989;
assign x_29437 = v_995 | ~v_990;
assign x_29438 = v_995 | ~v_856;
assign x_29439 = v_995 | ~v_991;
assign x_29440 = v_995 | ~v_992;
assign x_29441 = v_995 | ~v_182;
assign x_29442 = v_995 | ~v_179;
assign x_29443 = v_995 | ~v_163;
assign x_29444 = v_995 | ~v_161;
assign x_29445 = v_995 | ~v_136;
assign x_29446 = v_995 | ~v_135;
assign x_29447 = v_995 | ~v_134;
assign x_29448 = v_995 | ~v_993;
assign x_29449 = v_995 | ~v_994;
assign x_29450 = v_995 | ~v_18;
assign x_29451 = v_995 | ~v_17;
assign x_29452 = v_995 | ~v_16;
assign x_29453 = v_995 | ~v_14;
assign x_29454 = v_995 | ~v_9;
assign x_29455 = ~v_19 | ~v_49 | v_994;
assign x_29456 = ~v_34 | v_19 | v_993;
assign x_29457 = ~v_48 | ~v_156 | v_992;
assign x_29458 = ~v_5 | ~v_157 | v_991;
assign x_29459 = ~v_33 | v_156 | v_990;
assign x_29460 = ~v_1 | v_157 | v_989;
assign x_29461 = ~v_46 | ~v_152 | v_988;
assign x_29462 = ~v_38 | ~v_153 | v_987;
assign x_29463 = ~v_31 | v_152 | v_986;
assign x_29464 = ~v_23 | v_153 | v_985;
assign x_29465 = ~v_47 | ~v_156 | v_984;
assign x_29466 = ~v_42 | ~v_157 | v_983;
assign x_29467 = ~v_32 | v_156 | v_982;
assign x_29468 = ~v_27 | v_157 | v_981;
assign x_29469 = ~v_979 | ~v_964 | ~v_949 | v_980;
assign x_29470 = v_979 | ~v_809;
assign x_29471 = v_979 | ~v_810;
assign x_29472 = v_979 | ~v_811;
assign x_29473 = v_979 | ~v_812;
assign x_29474 = v_979 | ~v_965;
assign x_29475 = v_979 | ~v_966;
assign x_29476 = v_979 | ~v_967;
assign x_29477 = v_979 | ~v_968;
assign x_29478 = v_979 | ~v_873;
assign x_29479 = v_979 | ~v_874;
assign x_29480 = v_979 | ~v_875;
assign x_29481 = v_979 | ~v_876;
assign x_29482 = v_979 | ~v_817;
assign x_29483 = v_979 | ~v_820;
assign x_29484 = v_979 | ~v_877;
assign x_29485 = v_979 | ~v_878;
assign x_29486 = v_979 | ~v_879;
assign x_29487 = v_979 | ~v_880;
assign x_29488 = v_979 | ~v_969;
assign x_29489 = v_979 | ~v_970;
assign x_29490 = v_979 | ~v_971;
assign x_29491 = v_979 | ~v_972;
assign x_29492 = v_979 | ~v_827;
assign x_29493 = v_979 | ~v_830;
assign x_29494 = v_979 | ~v_973;
assign x_29495 = v_979 | ~v_974;
assign x_29496 = v_979 | ~v_885;
assign x_29497 = v_979 | ~v_886;
assign x_29498 = v_979 | ~v_975;
assign x_29499 = v_979 | ~v_976;
assign x_29500 = v_979 | ~v_977;
assign x_29501 = v_979 | ~v_978;
assign x_29502 = v_979 | ~v_184;
assign x_29503 = v_979 | ~v_181;
assign x_29504 = v_979 | ~v_172;
assign x_29505 = v_979 | ~v_171;
assign x_29506 = v_979 | ~v_169;
assign x_29507 = v_979 | ~v_150;
assign x_29508 = v_979 | ~v_149;
assign x_29509 = v_979 | ~v_147;
assign x_29510 = v_979 | ~v_102;
assign x_29511 = v_979 | ~v_101;
assign x_29512 = v_979 | ~v_96;
assign x_29513 = v_979 | ~v_94;
assign x_29514 = ~v_132 | ~v_177 | v_978;
assign x_29515 = ~v_117 | v_177 | v_977;
assign x_29516 = ~v_133 | ~v_154 | v_976;
assign x_29517 = ~v_118 | v_154 | v_975;
assign x_29518 = ~v_6 | ~v_178 | v_974;
assign x_29519 = ~v_3 | v_178 | v_973;
assign x_29520 = ~v_130 | ~v_154 | v_972;
assign x_29521 = ~v_122 | ~v_154 | v_971;
assign x_29522 = ~v_115 | v_154 | v_970;
assign x_29523 = ~v_107 | v_154 | v_969;
assign x_29524 = ~v_131 | ~v_177 | v_968;
assign x_29525 = ~v_126 | ~v_178 | v_967;
assign x_29526 = ~v_116 | v_177 | v_966;
assign x_29527 = ~v_111 | v_178 | v_965;
assign x_29528 = v_964 | ~v_776;
assign x_29529 = v_964 | ~v_777;
assign x_29530 = v_964 | ~v_778;
assign x_29531 = v_964 | ~v_779;
assign x_29532 = v_964 | ~v_950;
assign x_29533 = v_964 | ~v_951;
assign x_29534 = v_964 | ~v_952;
assign x_29535 = v_964 | ~v_953;
assign x_29536 = v_964 | ~v_858;
assign x_29537 = v_964 | ~v_859;
assign x_29538 = v_964 | ~v_860;
assign x_29539 = v_964 | ~v_861;
assign x_29540 = v_964 | ~v_784;
assign x_29541 = v_964 | ~v_787;
assign x_29542 = v_964 | ~v_862;
assign x_29543 = v_964 | ~v_863;
assign x_29544 = v_964 | ~v_864;
assign x_29545 = v_964 | ~v_865;
assign x_29546 = v_964 | ~v_954;
assign x_29547 = v_964 | ~v_955;
assign x_29548 = v_964 | ~v_956;
assign x_29549 = v_964 | ~v_957;
assign x_29550 = v_964 | ~v_794;
assign x_29551 = v_964 | ~v_797;
assign x_29552 = v_964 | ~v_958;
assign x_29553 = v_964 | ~v_959;
assign x_29554 = v_964 | ~v_870;
assign x_29555 = v_964 | ~v_871;
assign x_29556 = v_964 | ~v_960;
assign x_29557 = v_964 | ~v_961;
assign x_29558 = v_964 | ~v_962;
assign x_29559 = v_964 | ~v_963;
assign x_29560 = v_964 | ~v_183;
assign x_29561 = v_964 | ~v_180;
assign x_29562 = v_964 | ~v_168;
assign x_29563 = v_964 | ~v_167;
assign x_29564 = v_964 | ~v_165;
assign x_29565 = v_964 | ~v_145;
assign x_29566 = v_964 | ~v_144;
assign x_29567 = v_964 | ~v_142;
assign x_29568 = v_964 | ~v_60;
assign x_29569 = v_964 | ~v_59;
assign x_29570 = v_964 | ~v_54;
assign x_29571 = v_964 | ~v_52;
assign x_29572 = ~v_90 | ~v_177 | v_963;
assign x_29573 = ~v_75 | v_177 | v_962;
assign x_29574 = ~v_91 | ~v_154 | v_961;
assign x_29575 = ~v_76 | v_154 | v_960;
assign x_29576 = ~v_4 | ~v_178 | v_959;
assign x_29577 = ~v_2 | v_178 | v_958;
assign x_29578 = ~v_88 | ~v_154 | v_957;
assign x_29579 = ~v_80 | ~v_154 | v_956;
assign x_29580 = ~v_73 | v_154 | v_955;
assign x_29581 = ~v_65 | v_154 | v_954;
assign x_29582 = ~v_89 | ~v_177 | v_953;
assign x_29583 = ~v_84 | ~v_178 | v_952;
assign x_29584 = ~v_74 | v_177 | v_951;
assign x_29585 = ~v_69 | v_178 | v_950;
assign x_29586 = v_949 | ~v_743;
assign x_29587 = v_949 | ~v_744;
assign x_29588 = v_949 | ~v_745;
assign x_29589 = v_949 | ~v_746;
assign x_29590 = v_949 | ~v_935;
assign x_29591 = v_949 | ~v_936;
assign x_29592 = v_949 | ~v_937;
assign x_29593 = v_949 | ~v_938;
assign x_29594 = v_949 | ~v_843;
assign x_29595 = v_949 | ~v_844;
assign x_29596 = v_949 | ~v_845;
assign x_29597 = v_949 | ~v_846;
assign x_29598 = v_949 | ~v_751;
assign x_29599 = v_949 | ~v_754;
assign x_29600 = v_949 | ~v_847;
assign x_29601 = v_949 | ~v_848;
assign x_29602 = v_949 | ~v_849;
assign x_29603 = v_949 | ~v_850;
assign x_29604 = v_949 | ~v_939;
assign x_29605 = v_949 | ~v_940;
assign x_29606 = v_949 | ~v_941;
assign x_29607 = v_949 | ~v_942;
assign x_29608 = v_949 | ~v_761;
assign x_29609 = v_949 | ~v_764;
assign x_29610 = v_949 | ~v_943;
assign x_29611 = v_949 | ~v_944;
assign x_29612 = v_949 | ~v_855;
assign x_29613 = v_949 | ~v_856;
assign x_29614 = v_949 | ~v_945;
assign x_29615 = v_949 | ~v_946;
assign x_29616 = v_949 | ~v_947;
assign x_29617 = v_949 | ~v_948;
assign x_29618 = v_949 | ~v_182;
assign x_29619 = v_949 | ~v_179;
assign x_29620 = v_949 | ~v_164;
assign x_29621 = v_949 | ~v_163;
assign x_29622 = v_949 | ~v_161;
assign x_29623 = v_949 | ~v_137;
assign x_29624 = v_949 | ~v_136;
assign x_29625 = v_949 | ~v_134;
assign x_29626 = v_949 | ~v_17;
assign x_29627 = v_949 | ~v_16;
assign x_29628 = v_949 | ~v_11;
assign x_29629 = v_949 | ~v_9;
assign x_29630 = ~v_48 | ~v_177 | v_948;
assign x_29631 = ~v_33 | v_177 | v_947;
assign x_29632 = ~v_49 | ~v_154 | v_946;
assign x_29633 = ~v_34 | v_154 | v_945;
assign x_29634 = ~v_5 | ~v_178 | v_944;
assign x_29635 = ~v_1 | v_178 | v_943;
assign x_29636 = ~v_46 | ~v_154 | v_942;
assign x_29637 = ~v_38 | ~v_154 | v_941;
assign x_29638 = ~v_31 | v_154 | v_940;
assign x_29639 = ~v_23 | v_154 | v_939;
assign x_29640 = ~v_47 | ~v_177 | v_938;
assign x_29641 = ~v_42 | ~v_178 | v_937;
assign x_29642 = ~v_32 | v_177 | v_936;
assign x_29643 = ~v_27 | v_178 | v_935;
assign x_29644 = ~v_933 | ~v_918 | ~v_903 | v_934;
assign x_29645 = v_933 | ~v_809;
assign x_29646 = v_933 | ~v_810;
assign x_29647 = v_933 | ~v_811;
assign x_29648 = v_933 | ~v_812;
assign x_29649 = v_933 | ~v_919;
assign x_29650 = v_933 | ~v_920;
assign x_29651 = v_933 | ~v_873;
assign x_29652 = v_933 | ~v_874;
assign x_29653 = v_933 | ~v_875;
assign x_29654 = v_933 | ~v_876;
assign x_29655 = v_933 | ~v_817;
assign x_29656 = v_933 | ~v_820;
assign x_29657 = v_933 | ~v_877;
assign x_29658 = v_933 | ~v_878;
assign x_29659 = v_933 | ~v_879;
assign x_29660 = v_933 | ~v_880;
assign x_29661 = v_933 | ~v_921;
assign x_29662 = v_933 | ~v_922;
assign x_29663 = v_933 | ~v_923;
assign x_29664 = v_933 | ~v_924;
assign x_29665 = v_933 | ~v_827;
assign x_29666 = v_933 | ~v_830;
assign x_29667 = v_933 | ~v_925;
assign x_29668 = v_933 | ~v_926;
assign x_29669 = v_933 | ~v_885;
assign x_29670 = v_933 | ~v_886;
assign x_29671 = v_933 | ~v_927;
assign x_29672 = v_933 | ~v_928;
assign x_29673 = v_933 | ~v_929;
assign x_29674 = v_933 | ~v_930;
assign x_29675 = v_933 | ~v_931;
assign x_29676 = v_933 | ~v_932;
assign x_29677 = v_933 | ~v_184;
assign x_29678 = v_933 | ~v_181;
assign x_29679 = v_933 | ~v_171;
assign x_29680 = v_933 | ~v_169;
assign x_29681 = v_933 | ~v_150;
assign x_29682 = v_933 | ~v_149;
assign x_29683 = v_933 | ~v_148;
assign x_29684 = v_933 | ~v_147;
assign x_29685 = v_933 | ~v_103;
assign x_29686 = v_933 | ~v_102;
assign x_29687 = v_933 | ~v_101;
assign x_29688 = v_933 | ~v_94;
assign x_29689 = ~v_131 | ~v_175 | v_932;
assign x_29690 = ~v_116 | v_175 | v_931;
assign x_29691 = ~v_117 | v_175 | v_930;
assign x_29692 = ~v_132 | ~v_175 | v_929;
assign x_29693 = ~v_133 | ~v_141 | v_928;
assign x_29694 = ~v_118 | v_141 | v_927;
assign x_29695 = ~v_6 | ~v_176 | v_926;
assign x_29696 = ~v_3 | v_176 | v_925;
assign x_29697 = ~v_130 | ~v_173 | v_924;
assign x_29698 = ~v_122 | ~v_174 | v_923;
assign x_29699 = ~v_115 | v_173 | v_922;
assign x_29700 = ~v_107 | v_174 | v_921;
assign x_29701 = ~v_126 | ~v_176 | v_920;
assign x_29702 = ~v_111 | v_176 | v_919;
assign x_29703 = v_918 | ~v_776;
assign x_29704 = v_918 | ~v_777;
assign x_29705 = v_918 | ~v_778;
assign x_29706 = v_918 | ~v_779;
assign x_29707 = v_918 | ~v_904;
assign x_29708 = v_918 | ~v_905;
assign x_29709 = v_918 | ~v_858;
assign x_29710 = v_918 | ~v_859;
assign x_29711 = v_918 | ~v_860;
assign x_29712 = v_918 | ~v_861;
assign x_29713 = v_918 | ~v_784;
assign x_29714 = v_918 | ~v_787;
assign x_29715 = v_918 | ~v_862;
assign x_29716 = v_918 | ~v_863;
assign x_29717 = v_918 | ~v_864;
assign x_29718 = v_918 | ~v_865;
assign x_29719 = v_918 | ~v_906;
assign x_29720 = v_918 | ~v_907;
assign x_29721 = v_918 | ~v_908;
assign x_29722 = v_918 | ~v_909;
assign x_29723 = v_918 | ~v_794;
assign x_29724 = v_918 | ~v_797;
assign x_29725 = v_918 | ~v_910;
assign x_29726 = v_918 | ~v_911;
assign x_29727 = v_918 | ~v_870;
assign x_29728 = v_918 | ~v_871;
assign x_29729 = v_918 | ~v_912;
assign x_29730 = v_918 | ~v_913;
assign x_29731 = v_918 | ~v_914;
assign x_29732 = v_918 | ~v_915;
assign x_29733 = v_918 | ~v_916;
assign x_29734 = v_918 | ~v_917;
assign x_29735 = v_918 | ~v_183;
assign x_29736 = v_918 | ~v_180;
assign x_29737 = v_918 | ~v_167;
assign x_29738 = v_918 | ~v_165;
assign x_29739 = v_918 | ~v_145;
assign x_29740 = v_918 | ~v_144;
assign x_29741 = v_918 | ~v_143;
assign x_29742 = v_918 | ~v_142;
assign x_29743 = v_918 | ~v_61;
assign x_29744 = v_918 | ~v_60;
assign x_29745 = v_918 | ~v_59;
assign x_29746 = v_918 | ~v_52;
assign x_29747 = ~v_89 | ~v_175 | v_917;
assign x_29748 = ~v_74 | v_175 | v_916;
assign x_29749 = ~v_75 | v_175 | v_915;
assign x_29750 = ~v_90 | ~v_175 | v_914;
assign x_29751 = ~v_91 | ~v_141 | v_913;
assign x_29752 = ~v_76 | v_141 | v_912;
assign x_29753 = ~v_4 | ~v_176 | v_911;
assign x_29754 = ~v_2 | v_176 | v_910;
assign x_29755 = ~v_88 | ~v_173 | v_909;
assign x_29756 = ~v_80 | ~v_174 | v_908;
assign x_29757 = ~v_73 | v_173 | v_907;
assign x_29758 = ~v_65 | v_174 | v_906;
assign x_29759 = ~v_84 | ~v_176 | v_905;
assign x_29760 = ~v_69 | v_176 | v_904;
assign x_29761 = v_903 | ~v_743;
assign x_29762 = v_903 | ~v_744;
assign x_29763 = v_903 | ~v_745;
assign x_29764 = v_903 | ~v_746;
assign x_29765 = v_903 | ~v_889;
assign x_29766 = v_903 | ~v_890;
assign x_29767 = v_903 | ~v_843;
assign x_29768 = v_903 | ~v_844;
assign x_29769 = v_903 | ~v_845;
assign x_29770 = v_903 | ~v_846;
assign x_29771 = v_903 | ~v_751;
assign x_29772 = v_903 | ~v_754;
assign x_29773 = v_903 | ~v_847;
assign x_29774 = v_903 | ~v_848;
assign x_29775 = v_903 | ~v_849;
assign x_29776 = v_903 | ~v_850;
assign x_29777 = v_903 | ~v_891;
assign x_29778 = v_903 | ~v_892;
assign x_29779 = v_903 | ~v_893;
assign x_29780 = v_903 | ~v_894;
assign x_29781 = v_903 | ~v_761;
assign x_29782 = v_903 | ~v_764;
assign x_29783 = v_903 | ~v_895;
assign x_29784 = v_903 | ~v_896;
assign x_29785 = v_903 | ~v_855;
assign x_29786 = v_903 | ~v_856;
assign x_29787 = v_903 | ~v_897;
assign x_29788 = v_903 | ~v_898;
assign x_29789 = v_903 | ~v_899;
assign x_29790 = v_903 | ~v_900;
assign x_29791 = v_903 | ~v_901;
assign x_29792 = v_903 | ~v_902;
assign x_29793 = v_903 | ~v_182;
assign x_29794 = v_903 | ~v_179;
assign x_29795 = v_903 | ~v_163;
assign x_29796 = v_903 | ~v_161;
assign x_29797 = v_903 | ~v_137;
assign x_29798 = v_903 | ~v_136;
assign x_29799 = v_903 | ~v_135;
assign x_29800 = v_903 | ~v_134;
assign x_29801 = v_903 | ~v_18;
assign x_29802 = v_903 | ~v_17;
assign x_29803 = v_903 | ~v_16;
assign x_29804 = v_903 | ~v_9;
assign x_29805 = ~v_47 | ~v_175 | v_902;
assign x_29806 = ~v_32 | v_175 | v_901;
assign x_29807 = ~v_33 | v_175 | v_900;
assign x_29808 = ~v_48 | ~v_175 | v_899;
assign x_29809 = ~v_49 | ~v_141 | v_898;
assign x_29810 = ~v_34 | v_141 | v_897;
assign x_29811 = ~v_5 | ~v_176 | v_896;
assign x_29812 = ~v_1 | v_176 | v_895;
assign x_29813 = ~v_46 | ~v_173 | v_894;
assign x_29814 = ~v_38 | ~v_174 | v_893;
assign x_29815 = ~v_31 | v_173 | v_892;
assign x_29816 = ~v_23 | v_174 | v_891;
assign x_29817 = ~v_42 | ~v_176 | v_890;
assign x_29818 = ~v_27 | v_176 | v_889;
assign x_29819 = ~v_887 | ~v_872 | ~v_857 | v_888;
assign x_29820 = v_887 | ~v_809;
assign x_29821 = v_887 | ~v_810;
assign x_29822 = v_887 | ~v_811;
assign x_29823 = v_887 | ~v_812;
assign x_29824 = v_887 | ~v_813;
assign x_29825 = v_887 | ~v_814;
assign x_29826 = v_887 | ~v_815;
assign x_29827 = v_887 | ~v_816;
assign x_29828 = v_887 | ~v_873;
assign x_29829 = v_887 | ~v_874;
assign x_29830 = v_887 | ~v_875;
assign x_29831 = v_887 | ~v_876;
assign x_29832 = v_887 | ~v_817;
assign x_29833 = v_887 | ~v_820;
assign x_29834 = v_887 | ~v_877;
assign x_29835 = v_887 | ~v_878;
assign x_29836 = v_887 | ~v_879;
assign x_29837 = v_887 | ~v_880;
assign x_29838 = v_887 | ~v_823;
assign x_29839 = v_887 | ~v_824;
assign x_29840 = v_887 | ~v_825;
assign x_29841 = v_887 | ~v_826;
assign x_29842 = v_887 | ~v_827;
assign x_29843 = v_887 | ~v_830;
assign x_29844 = v_887 | ~v_881;
assign x_29845 = v_887 | ~v_882;
assign x_29846 = v_887 | ~v_883;
assign x_29847 = v_887 | ~v_884;
assign x_29848 = v_887 | ~v_885;
assign x_29849 = v_887 | ~v_886;
assign x_29850 = v_887 | ~v_837;
assign x_29851 = v_887 | ~v_838;
assign x_29852 = v_887 | ~v_184;
assign x_29853 = v_887 | ~v_181;
assign x_29854 = v_887 | ~v_171;
assign x_29855 = v_887 | ~v_169;
assign x_29856 = v_887 | ~v_160;
assign x_29857 = v_887 | ~v_150;
assign x_29858 = v_887 | ~v_148;
assign x_29859 = v_887 | ~v_103;
assign x_29860 = v_887 | ~v_102;
assign x_29861 = v_887 | ~v_97;
assign x_29862 = v_887 | ~v_95;
assign x_29863 = v_887 | ~v_94;
assign x_29864 = ~v_129 | ~v_158 | v_886;
assign x_29865 = ~v_114 | v_158 | v_885;
assign x_29866 = ~v_132 | ~v_158 | v_884;
assign x_29867 = ~v_6 | ~v_158 | v_883;
assign x_29868 = ~v_117 | v_158 | v_882;
assign x_29869 = ~v_3 | v_158 | v_881;
assign x_29870 = ~v_127 | ~v_178 | v_880;
assign x_29871 = ~v_121 | ~v_177 | v_879;
assign x_29872 = ~v_112 | v_178 | v_878;
assign x_29873 = ~v_106 | v_177 | v_877;
assign x_29874 = ~v_128 | ~v_158 | v_876;
assign x_29875 = ~v_125 | ~v_158 | v_875;
assign x_29876 = ~v_113 | v_158 | v_874;
assign x_29877 = ~v_110 | v_158 | v_873;
assign x_29878 = v_872 | ~v_776;
assign x_29879 = v_872 | ~v_777;
assign x_29880 = v_872 | ~v_778;
assign x_29881 = v_872 | ~v_779;
assign x_29882 = v_872 | ~v_780;
assign x_29883 = v_872 | ~v_781;
assign x_29884 = v_872 | ~v_782;
assign x_29885 = v_872 | ~v_783;
assign x_29886 = v_872 | ~v_858;
assign x_29887 = v_872 | ~v_859;
assign x_29888 = v_872 | ~v_860;
assign x_29889 = v_872 | ~v_861;
assign x_29890 = v_872 | ~v_784;
assign x_29891 = v_872 | ~v_787;
assign x_29892 = v_872 | ~v_862;
assign x_29893 = v_872 | ~v_863;
assign x_29894 = v_872 | ~v_864;
assign x_29895 = v_872 | ~v_865;
assign x_29896 = v_872 | ~v_790;
assign x_29897 = v_872 | ~v_791;
assign x_29898 = v_872 | ~v_792;
assign x_29899 = v_872 | ~v_793;
assign x_29900 = v_872 | ~v_794;
assign x_29901 = v_872 | ~v_797;
assign x_29902 = v_872 | ~v_866;
assign x_29903 = v_872 | ~v_867;
assign x_29904 = v_872 | ~v_868;
assign x_29905 = v_872 | ~v_869;
assign x_29906 = v_872 | ~v_870;
assign x_29907 = v_872 | ~v_871;
assign x_29908 = v_872 | ~v_804;
assign x_29909 = v_872 | ~v_805;
assign x_29910 = v_872 | ~v_183;
assign x_29911 = v_872 | ~v_180;
assign x_29912 = v_872 | ~v_167;
assign x_29913 = v_872 | ~v_165;
assign x_29914 = v_872 | ~v_159;
assign x_29915 = v_872 | ~v_145;
assign x_29916 = v_872 | ~v_143;
assign x_29917 = v_872 | ~v_61;
assign x_29918 = v_872 | ~v_60;
assign x_29919 = v_872 | ~v_55;
assign x_29920 = v_872 | ~v_53;
assign x_29921 = v_872 | ~v_52;
assign x_29922 = ~v_87 | ~v_158 | v_871;
assign x_29923 = ~v_72 | v_158 | v_870;
assign x_29924 = ~v_90 | ~v_158 | v_869;
assign x_29925 = ~v_4 | ~v_158 | v_868;
assign x_29926 = ~v_75 | v_158 | v_867;
assign x_29927 = ~v_2 | v_158 | v_866;
assign x_29928 = ~v_85 | ~v_178 | v_865;
assign x_29929 = ~v_79 | ~v_177 | v_864;
assign x_29930 = ~v_70 | v_178 | v_863;
assign x_29931 = ~v_64 | v_177 | v_862;
assign x_29932 = ~v_86 | ~v_158 | v_861;
assign x_29933 = ~v_83 | ~v_158 | v_860;
assign x_29934 = ~v_71 | v_158 | v_859;
assign x_29935 = ~v_68 | v_158 | v_858;
assign x_29936 = v_857 | ~v_743;
assign x_29937 = v_857 | ~v_744;
assign x_29938 = v_857 | ~v_745;
assign x_29939 = v_857 | ~v_746;
assign x_29940 = v_857 | ~v_747;
assign x_29941 = v_857 | ~v_748;
assign x_29942 = v_857 | ~v_749;
assign x_29943 = v_857 | ~v_750;
assign x_29944 = v_857 | ~v_843;
assign x_29945 = v_857 | ~v_844;
assign x_29946 = v_857 | ~v_845;
assign x_29947 = v_857 | ~v_846;
assign x_29948 = v_857 | ~v_751;
assign x_29949 = v_857 | ~v_754;
assign x_29950 = v_857 | ~v_847;
assign x_29951 = v_857 | ~v_848;
assign x_29952 = v_857 | ~v_849;
assign x_29953 = v_857 | ~v_850;
assign x_29954 = v_857 | ~v_757;
assign x_29955 = v_857 | ~v_758;
assign x_29956 = v_857 | ~v_759;
assign x_29957 = v_857 | ~v_760;
assign x_29958 = v_857 | ~v_761;
assign x_29959 = v_857 | ~v_764;
assign x_29960 = v_857 | ~v_851;
assign x_29961 = v_857 | ~v_852;
assign x_29962 = v_857 | ~v_853;
assign x_29963 = v_857 | ~v_854;
assign x_29964 = v_857 | ~v_855;
assign x_29965 = v_857 | ~v_856;
assign x_29966 = v_857 | ~v_771;
assign x_29967 = v_857 | ~v_772;
assign x_29968 = v_857 | ~v_182;
assign x_29969 = v_857 | ~v_179;
assign x_29970 = v_857 | ~v_163;
assign x_29971 = v_857 | ~v_161;
assign x_29972 = v_857 | ~v_155;
assign x_29973 = v_857 | ~v_137;
assign x_29974 = v_857 | ~v_135;
assign x_29975 = v_857 | ~v_18;
assign x_29976 = v_857 | ~v_17;
assign x_29977 = v_857 | ~v_12;
assign x_29978 = v_857 | ~v_10;
assign x_29979 = v_857 | ~v_9;
assign x_29980 = ~v_45 | ~v_158 | v_856;
assign x_29981 = ~v_30 | v_158 | v_855;
assign x_29982 = ~v_48 | ~v_158 | v_854;
assign x_29983 = ~v_5 | ~v_158 | v_853;
assign x_29984 = ~v_33 | v_158 | v_852;
assign x_29985 = ~v_1 | v_158 | v_851;
assign x_29986 = ~v_43 | ~v_178 | v_850;
assign x_29987 = ~v_37 | ~v_177 | v_849;
assign x_29988 = ~v_28 | v_178 | v_848;
assign x_29989 = ~v_22 | v_177 | v_847;
assign x_29990 = ~v_44 | ~v_158 | v_846;
assign x_29991 = ~v_41 | ~v_158 | v_845;
assign x_29992 = ~v_29 | v_158 | v_844;
assign x_29993 = ~v_26 | v_158 | v_843;
assign x_29994 = ~v_841 | ~v_808 | ~v_775 | v_842;
assign x_29995 = v_841 | ~v_809;
assign x_29996 = v_841 | ~v_810;
assign x_29997 = v_841 | ~v_811;
assign x_29998 = v_841 | ~v_812;
assign x_29999 = v_841 | ~v_813;
assign x_30000 = v_841 | ~v_814;
assign x_30001 = v_841 | ~v_815;
assign x_30002 = v_841 | ~v_816;
assign x_30003 = v_841 | ~v_817;
assign x_30004 = v_841 | ~v_818;
assign x_30005 = v_841 | ~v_819;
assign x_30006 = v_841 | ~v_820;
assign x_30007 = v_841 | ~v_821;
assign x_30008 = v_841 | ~v_822;
assign x_30009 = v_841 | ~v_823;
assign x_30010 = v_841 | ~v_824;
assign x_30011 = v_841 | ~v_825;
assign x_30012 = v_841 | ~v_826;
assign x_30013 = v_841 | ~v_827;
assign x_30014 = v_841 | ~v_828;
assign x_30015 = v_841 | ~v_829;
assign x_30016 = v_841 | ~v_830;
assign x_30017 = v_841 | ~v_831;
assign x_30018 = v_841 | ~v_832;
assign x_30019 = v_841 | ~v_833;
assign x_30020 = v_841 | ~v_834;
assign x_30021 = v_841 | ~v_835;
assign x_30022 = v_841 | ~v_836;
assign x_30023 = v_841 | ~v_837;
assign x_30024 = v_841 | ~v_838;
assign x_30025 = v_841 | ~v_839;
assign x_30026 = v_841 | ~v_840;
assign x_30027 = v_841 | ~v_184;
assign x_30028 = v_841 | ~v_170;
assign x_30029 = v_841 | ~v_169;
assign x_30030 = v_841 | ~v_160;
assign x_30031 = v_841 | ~v_150;
assign x_30032 = v_841 | ~v_148;
assign x_30033 = v_841 | ~v_147;
assign x_30034 = v_841 | ~v_103;
assign x_30035 = v_841 | ~v_102;
assign x_30036 = v_841 | ~v_100;
assign x_30037 = v_841 | ~v_98;
assign x_30038 = v_841 | ~v_97;
assign x_30039 = ~v_19 | ~v_129 | v_840;
assign x_30040 = v_19 | ~v_114 | v_839;
assign x_30041 = ~v_133 | ~v_158 | v_838;
assign x_30042 = ~v_118 | v_158 | v_837;
assign x_30043 = ~v_132 | ~v_157 | v_836;
assign x_30044 = ~v_6 | ~v_156 | v_835;
assign x_30045 = ~v_117 | v_157 | v_834;
assign x_30046 = ~v_3 | v_156 | v_833;
assign x_30047 = ~v_127 | ~v_152 | v_832;
assign x_30048 = ~v_121 | ~v_153 | v_831;
assign x_30049 = ~v_119 | ~v_154 | v_830;
assign x_30050 = ~v_112 | v_152 | v_829;
assign x_30051 = ~v_106 | v_153 | v_828;
assign x_30052 = ~v_104 | v_154 | v_827;
assign x_30053 = ~v_130 | ~v_178 | v_826;
assign x_30054 = ~v_122 | ~v_177 | v_825;
assign x_30055 = ~v_115 | v_178 | v_824;
assign x_30056 = ~v_107 | v_177 | v_823;
assign x_30057 = ~v_128 | ~v_156 | v_822;
assign x_30058 = ~v_125 | ~v_157 | v_821;
assign x_30059 = ~v_124 | ~v_158 | v_820;
assign x_30060 = ~v_113 | v_156 | v_819;
assign x_30061 = ~v_110 | v_157 | v_818;
assign x_30062 = ~v_109 | v_158 | v_817;
assign x_30063 = ~v_131 | ~v_158 | v_816;
assign x_30064 = ~v_126 | ~v_158 | v_815;
assign x_30065 = ~v_116 | v_158 | v_814;
assign x_30066 = ~v_111 | v_158 | v_813;
assign x_30067 = ~v_123 | ~v_178 | v_812;
assign x_30068 = ~v_120 | ~v_177 | v_811;
assign x_30069 = ~v_108 | v_178 | v_810;
assign x_30070 = ~v_105 | v_177 | v_809;
assign x_30071 = v_808 | ~v_776;
assign x_30072 = v_808 | ~v_777;
assign x_30073 = v_808 | ~v_778;
assign x_30074 = v_808 | ~v_779;
assign x_30075 = v_808 | ~v_780;
assign x_30076 = v_808 | ~v_781;
assign x_30077 = v_808 | ~v_782;
assign x_30078 = v_808 | ~v_783;
assign x_30079 = v_808 | ~v_784;
assign x_30080 = v_808 | ~v_785;
assign x_30081 = v_808 | ~v_786;
assign x_30082 = v_808 | ~v_787;
assign x_30083 = v_808 | ~v_788;
assign x_30084 = v_808 | ~v_789;
assign x_30085 = v_808 | ~v_790;
assign x_30086 = v_808 | ~v_791;
assign x_30087 = v_808 | ~v_792;
assign x_30088 = v_808 | ~v_793;
assign x_30089 = v_808 | ~v_794;
assign x_30090 = v_808 | ~v_795;
assign x_30091 = v_808 | ~v_796;
assign x_30092 = v_808 | ~v_797;
assign x_30093 = v_808 | ~v_798;
assign x_30094 = v_808 | ~v_799;
assign x_30095 = v_808 | ~v_800;
assign x_30096 = v_808 | ~v_801;
assign x_30097 = v_808 | ~v_802;
assign x_30098 = v_808 | ~v_803;
assign x_30099 = v_808 | ~v_804;
assign x_30100 = v_808 | ~v_805;
assign x_30101 = v_808 | ~v_806;
assign x_30102 = v_808 | ~v_807;
assign x_30103 = v_808 | ~v_183;
assign x_30104 = v_808 | ~v_166;
assign x_30105 = v_808 | ~v_165;
assign x_30106 = v_808 | ~v_159;
assign x_30107 = v_808 | ~v_145;
assign x_30108 = v_808 | ~v_143;
assign x_30109 = v_808 | ~v_142;
assign x_30110 = v_808 | ~v_61;
assign x_30111 = v_808 | ~v_60;
assign x_30112 = v_808 | ~v_58;
assign x_30113 = v_808 | ~v_56;
assign x_30114 = v_808 | ~v_55;
assign x_30115 = ~v_19 | ~v_87 | v_807;
assign x_30116 = v_19 | ~v_72 | v_806;
assign x_30117 = ~v_91 | ~v_158 | v_805;
assign x_30118 = ~v_76 | v_158 | v_804;
assign x_30119 = ~v_90 | ~v_157 | v_803;
assign x_30120 = ~v_4 | ~v_156 | v_802;
assign x_30121 = ~v_75 | v_157 | v_801;
assign x_30122 = ~v_2 | v_156 | v_800;
assign x_30123 = ~v_85 | ~v_152 | v_799;
assign x_30124 = ~v_79 | ~v_153 | v_798;
assign x_30125 = ~v_77 | ~v_154 | v_797;
assign x_30126 = ~v_70 | v_152 | v_796;
assign x_30127 = ~v_64 | v_153 | v_795;
assign x_30128 = ~v_62 | v_154 | v_794;
assign x_30129 = ~v_88 | ~v_178 | v_793;
assign x_30130 = ~v_80 | ~v_177 | v_792;
assign x_30131 = ~v_73 | v_178 | v_791;
assign x_30132 = ~v_65 | v_177 | v_790;
assign x_30133 = ~v_86 | ~v_156 | v_789;
assign x_30134 = ~v_83 | ~v_157 | v_788;
assign x_30135 = ~v_82 | ~v_158 | v_787;
assign x_30136 = ~v_71 | v_156 | v_786;
assign x_30137 = ~v_68 | v_157 | v_785;
assign x_30138 = ~v_67 | v_158 | v_784;
assign x_30139 = ~v_89 | ~v_158 | v_783;
assign x_30140 = ~v_84 | ~v_158 | v_782;
assign x_30141 = ~v_74 | v_158 | v_781;
assign x_30142 = ~v_69 | v_158 | v_780;
assign x_30143 = ~v_81 | ~v_178 | v_779;
assign x_30144 = ~v_78 | ~v_177 | v_778;
assign x_30145 = ~v_66 | v_178 | v_777;
assign x_30146 = ~v_63 | v_177 | v_776;
assign x_30147 = v_775 | ~v_743;
assign x_30148 = v_775 | ~v_744;
assign x_30149 = v_775 | ~v_745;
assign x_30150 = v_775 | ~v_746;
assign x_30151 = v_775 | ~v_747;
assign x_30152 = v_775 | ~v_748;
assign x_30153 = v_775 | ~v_749;
assign x_30154 = v_775 | ~v_750;
assign x_30155 = v_775 | ~v_751;
assign x_30156 = v_775 | ~v_752;
assign x_30157 = v_775 | ~v_753;
assign x_30158 = v_775 | ~v_754;
assign x_30159 = v_775 | ~v_755;
assign x_30160 = v_775 | ~v_756;
assign x_30161 = v_775 | ~v_757;
assign x_30162 = v_775 | ~v_758;
assign x_30163 = v_775 | ~v_759;
assign x_30164 = v_775 | ~v_760;
assign x_30165 = v_775 | ~v_761;
assign x_30166 = v_775 | ~v_762;
assign x_30167 = v_775 | ~v_763;
assign x_30168 = v_775 | ~v_764;
assign x_30169 = v_775 | ~v_765;
assign x_30170 = v_775 | ~v_766;
assign x_30171 = v_775 | ~v_767;
assign x_30172 = v_775 | ~v_768;
assign x_30173 = v_775 | ~v_769;
assign x_30174 = v_775 | ~v_770;
assign x_30175 = v_775 | ~v_771;
assign x_30176 = v_775 | ~v_772;
assign x_30177 = v_775 | ~v_773;
assign x_30178 = v_775 | ~v_774;
assign x_30179 = v_775 | ~v_182;
assign x_30180 = v_775 | ~v_162;
assign x_30181 = v_775 | ~v_161;
assign x_30182 = v_775 | ~v_155;
assign x_30183 = v_775 | ~v_137;
assign x_30184 = v_775 | ~v_135;
assign x_30185 = v_775 | ~v_134;
assign x_30186 = v_775 | ~v_18;
assign x_30187 = v_775 | ~v_17;
assign x_30188 = v_775 | ~v_15;
assign x_30189 = v_775 | ~v_13;
assign x_30190 = v_775 | ~v_12;
assign x_30191 = ~v_19 | ~v_45 | v_774;
assign x_30192 = ~v_30 | v_19 | v_773;
assign x_30193 = ~v_49 | ~v_158 | v_772;
assign x_30194 = ~v_34 | v_158 | v_771;
assign x_30195 = ~v_48 | ~v_157 | v_770;
assign x_30196 = ~v_5 | ~v_156 | v_769;
assign x_30197 = ~v_33 | v_157 | v_768;
assign x_30198 = ~v_1 | v_156 | v_767;
assign x_30199 = ~v_43 | ~v_152 | v_766;
assign x_30200 = ~v_37 | ~v_153 | v_765;
assign x_30201 = ~v_35 | ~v_154 | v_764;
assign x_30202 = ~v_28 | v_152 | v_763;
assign x_30203 = ~v_22 | v_153 | v_762;
assign x_30204 = ~v_20 | v_154 | v_761;
assign x_30205 = ~v_46 | ~v_178 | v_760;
assign x_30206 = ~v_38 | ~v_177 | v_759;
assign x_30207 = ~v_31 | v_178 | v_758;
assign x_30208 = ~v_23 | v_177 | v_757;
assign x_30209 = ~v_44 | ~v_156 | v_756;
assign x_30210 = ~v_41 | ~v_157 | v_755;
assign x_30211 = ~v_40 | ~v_158 | v_754;
assign x_30212 = ~v_29 | v_156 | v_753;
assign x_30213 = ~v_26 | v_157 | v_752;
assign x_30214 = ~v_25 | v_158 | v_751;
assign x_30215 = ~v_47 | ~v_158 | v_750;
assign x_30216 = ~v_42 | ~v_158 | v_749;
assign x_30217 = ~v_32 | v_158 | v_748;
assign x_30218 = ~v_27 | v_158 | v_747;
assign x_30219 = ~v_39 | ~v_178 | v_746;
assign x_30220 = ~v_36 | ~v_177 | v_745;
assign x_30221 = ~v_24 | v_178 | v_744;
assign x_30222 = ~v_21 | v_177 | v_743;
assign x_30223 = v_742 | ~v_727;
assign x_30224 = v_742 | ~v_737;
assign x_30225 = v_741 | ~v_735;
assign x_30226 = v_741 | ~v_731;
assign x_30227 = v_740 | ~v_739;
assign x_30228 = v_740 | ~v_737;
assign x_30229 = v_157 | v_156 | ~v_738 | ~v_736 | v_739;
assign x_30230 = v_738 | ~v_737;
assign x_30231 = v_738 | ~v_730;
assign x_30232 = v_152 | v_153 | v_737;
assign x_30233 = v_736 | ~v_735;
assign x_30234 = v_736 | ~v_728;
assign x_30235 = v_176 | v_175 | v_735;
assign x_30236 = v_734 | ~v_733;
assign x_30237 = v_734 | ~v_731;
assign x_30238 = v_176 | v_175 | ~v_732 | ~v_729 | v_733;
assign x_30239 = v_732 | ~v_730;
assign x_30240 = v_732 | ~v_731;
assign x_30241 = v_174 | v_173 | v_731;
assign x_30242 = v_177 | v_178 | v_730;
assign x_30243 = v_729 | ~v_727;
assign x_30244 = v_729 | ~v_728;
assign x_30245 = v_140 | v_139 | v_728;
assign x_30246 = v_157 | v_156 | v_727;
assign x_30247 = ~v_725 | ~v_724 | ~v_723 | ~v_722 | ~v_721 | ~v_705 | ~v_689 | ~v_673 | ~v_657 | ~v_611 | ~v_595 | ~v_579 | ~v_563 | ~v_547 | ~v_501 | ~v_485 | ~v_439 | ~v_393 | ~v_347 | ~v_301 | ~v_201 | v_726;
assign x_30248 = v_725 | v_5;
assign x_30249 = v_725 | ~v_4;
assign x_30250 = v_724 | v_4;
assign x_30251 = v_724 | ~v_6;
assign x_30252 = v_723 | v_3;
assign x_30253 = v_723 | ~v_2;
assign x_30254 = v_722 | v_2;
assign x_30255 = v_722 | ~v_1;
assign x_30256 = v_721 | ~v_710;
assign x_30257 = v_721 | ~v_715;
assign x_30258 = v_721 | ~v_720;
assign x_30259 = v_98 | v_103 | v_101 | v_100 | v_95 | v_99 | v_102 | ~v_719 | ~v_718 | v_170 | v_169 | v_149 | v_148 | v_184 | ~v_483 | ~v_717 | ~v_299 | ~v_482 | ~v_716 | ~v_298 | ~v_477 | ~v_291 | ~v_476 | ~v_290 | ~v_289 | ~v_475 | ~v_288 | ~v_474 | ~v_287 | ~v_286 | ~v_473 | ~v_281 | ~v_472 | ~v_280 | ~v_279 | ~v_471 | ~v_278 | ~v_470 | ~v_277 | ~v_276 | ~v_271 | ~v_270 | ~v_269 | ~v_268 | v_720;
assign x_30260 = v_719 | v_3;
assign x_30261 = v_719 | ~v_19;
assign x_30262 = v_718 | v_19;
assign x_30263 = v_718 | v_6;
assign x_30264 = v_717 | v_132;
assign x_30265 = v_717 | v_19;
assign x_30266 = v_716 | v_117;
assign x_30267 = v_716 | ~v_19;
assign x_30268 = v_53 | v_56 | v_61 | v_60 | v_59 | v_58 | v_57 | ~v_714 | ~v_713 | v_144 | v_143 | v_166 | v_165 | v_183 | ~v_266 | ~v_468 | ~v_712 | ~v_467 | ~v_711 | ~v_265 | ~v_462 | ~v_258 | ~v_461 | ~v_257 | ~v_256 | ~v_460 | ~v_255 | ~v_459 | ~v_254 | ~v_253 | ~v_458 | ~v_248 | ~v_457 | ~v_247 | ~v_246 | ~v_456 | ~v_245 | ~v_455 | ~v_244 | ~v_243 | ~v_238 | ~v_237 | ~v_236 | ~v_235 | v_715;
assign x_30269 = v_714 | v_2;
assign x_30270 = v_714 | ~v_19;
assign x_30271 = v_713 | v_19;
assign x_30272 = v_713 | v_4;
assign x_30273 = v_712 | v_90;
assign x_30274 = v_712 | v_19;
assign x_30275 = v_711 | v_75;
assign x_30276 = v_711 | ~v_19;
assign x_30277 = v_13 | v_18 | v_17 | v_16 | v_15 | v_14 | v_10 | ~v_453 | ~v_709 | ~v_452 | ~v_708 | v_136 | v_135 | ~v_707 | ~v_706 | v_162 | v_161 | v_182 | ~v_233 | ~v_232 | ~v_447 | ~v_225 | ~v_446 | ~v_224 | ~v_223 | ~v_445 | ~v_222 | ~v_444 | ~v_221 | ~v_220 | ~v_443 | ~v_215 | ~v_442 | ~v_214 | ~v_213 | ~v_441 | ~v_212 | ~v_440 | ~v_211 | ~v_210 | ~v_205 | ~v_204 | ~v_203 | ~v_202 | v_710;
assign x_30278 = v_709 | v_48;
assign x_30279 = v_709 | v_19;
assign x_30280 = v_708 | v_33;
assign x_30281 = v_708 | ~v_19;
assign x_30282 = v_707 | v_1;
assign x_30283 = v_707 | ~v_19;
assign x_30284 = v_706 | v_19;
assign x_30285 = v_706 | v_5;
assign x_30286 = v_705 | ~v_694;
assign x_30287 = v_705 | ~v_699;
assign x_30288 = v_705 | ~v_704;
assign x_30289 = v_103 | v_101 | v_100 | v_99 | v_93 | v_102 | v_171 | v_170 | v_149 | v_148 | v_147 | v_184 | ~v_703 | ~v_702 | ~v_483 | ~v_482 | ~v_701 | ~v_653 | ~v_700 | ~v_652 | ~v_477 | ~v_476 | ~v_289 | ~v_475 | ~v_474 | ~v_286 | ~v_649 | ~v_648 | ~v_647 | ~v_646 | ~v_473 | ~v_472 | ~v_279 | ~v_471 | ~v_470 | ~v_276 | ~v_645 | ~v_644 | ~v_643 | ~v_642 | ~v_271 | ~v_270 | ~v_269 | ~v_268 | v_704;
assign x_30290 = v_703 | v_152;
assign x_30291 = v_703 | v_132;
assign x_30292 = v_702 | ~v_152;
assign x_30293 = v_702 | v_117;
assign x_30294 = v_701 | v_153;
assign x_30295 = v_701 | v_6;
assign x_30296 = v_700 | ~v_153;
assign x_30297 = v_700 | v_3;
assign x_30298 = v_61 | v_51 | v_60 | v_59 | v_58 | v_57 | v_144 | v_143 | v_142 | v_167 | v_166 | v_183 | ~v_698 | ~v_697 | ~v_468 | ~v_467 | ~v_696 | ~v_638 | ~v_695 | ~v_637 | ~v_462 | ~v_461 | ~v_256 | ~v_460 | ~v_459 | ~v_253 | ~v_634 | ~v_633 | ~v_632 | ~v_631 | ~v_458 | ~v_457 | ~v_246 | ~v_456 | ~v_455 | ~v_243 | ~v_630 | ~v_629 | ~v_628 | ~v_627 | ~v_238 | ~v_237 | ~v_236 | ~v_235 | v_699;
assign x_30299 = v_698 | v_152;
assign x_30300 = v_698 | v_90;
assign x_30301 = v_697 | ~v_152;
assign x_30302 = v_697 | v_75;
assign x_30303 = v_696 | v_153;
assign x_30304 = v_696 | v_4;
assign x_30305 = v_695 | ~v_153;
assign x_30306 = v_695 | v_2;
assign x_30307 = v_18 | v_17 | v_16 | v_8 | v_15 | v_14 | ~v_453 | ~v_452 | v_136 | v_135 | v_134 | v_163 | v_162 | v_182 | ~v_693 | ~v_692 | ~v_691 | ~v_623 | ~v_690 | ~v_622 | ~v_447 | ~v_446 | ~v_223 | ~v_445 | ~v_444 | ~v_220 | ~v_619 | ~v_618 | ~v_617 | ~v_616 | ~v_443 | ~v_442 | ~v_213 | ~v_441 | ~v_440 | ~v_210 | ~v_615 | ~v_614 | ~v_613 | ~v_612 | ~v_205 | ~v_204 | ~v_203 | ~v_202 | v_694;
assign x_30308 = v_693 | v_152;
assign x_30309 = v_693 | v_48;
assign x_30310 = v_692 | ~v_152;
assign x_30311 = v_692 | v_33;
assign x_30312 = v_691 | v_153;
assign x_30313 = v_691 | v_5;
assign x_30314 = v_690 | ~v_153;
assign x_30315 = v_690 | v_1;
assign x_30316 = v_689 | ~v_678;
assign x_30317 = v_689 | ~v_683;
assign x_30318 = v_689 | ~v_688;
assign x_30319 = v_103 | v_101 | v_96 | v_100 | v_95 | v_93 | v_102 | v_171 | v_170 | v_150 | v_149 | v_184 | ~v_435 | ~v_434 | ~v_653 | ~v_652 | ~v_687 | ~v_686 | ~v_685 | ~v_684 | ~v_289 | ~v_286 | ~v_649 | ~v_648 | ~v_647 | ~v_646 | ~v_431 | ~v_430 | ~v_429 | ~v_428 | ~v_279 | ~v_276 | ~v_427 | ~v_426 | ~v_425 | ~v_424 | ~v_645 | ~v_644 | ~v_643 | ~v_642 | ~v_271 | ~v_270 | ~v_269 | ~v_268 | v_688;
assign x_30320 = v_687 | v_154;
assign x_30321 = v_687 | v_132;
assign x_30322 = v_686 | v_154;
assign x_30323 = v_686 | v_6;
assign x_30324 = v_685 | ~v_154;
assign x_30325 = v_685 | v_117;
assign x_30326 = v_684 | ~v_154;
assign x_30327 = v_684 | v_3;
assign x_30328 = v_54 | v_53 | v_61 | v_51 | v_60 | v_59 | v_58 | v_144 | v_145 | v_167 | v_166 | v_183 | ~v_420 | ~v_419 | ~v_638 | ~v_637 | ~v_682 | ~v_681 | ~v_680 | ~v_679 | ~v_256 | ~v_253 | ~v_634 | ~v_633 | ~v_632 | ~v_631 | ~v_416 | ~v_415 | ~v_414 | ~v_413 | ~v_246 | ~v_243 | ~v_412 | ~v_411 | ~v_410 | ~v_409 | ~v_630 | ~v_629 | ~v_628 | ~v_627 | ~v_238 | ~v_237 | ~v_236 | ~v_235 | v_683;
assign x_30329 = v_682 | v_154;
assign x_30330 = v_682 | v_90;
assign x_30331 = v_681 | v_154;
assign x_30332 = v_681 | v_4;
assign x_30333 = v_680 | ~v_154;
assign x_30334 = v_680 | v_75;
assign x_30335 = v_679 | ~v_154;
assign x_30336 = v_679 | v_2;
assign x_30337 = v_18 | v_17 | v_16 | v_8 | v_15 | v_11 | v_10 | v_136 | v_137 | v_163 | v_162 | v_182 | ~v_405 | ~v_404 | ~v_623 | ~v_622 | ~v_677 | ~v_676 | ~v_675 | ~v_674 | ~v_223 | ~v_220 | ~v_619 | ~v_618 | ~v_617 | ~v_616 | ~v_401 | ~v_400 | ~v_399 | ~v_398 | ~v_213 | ~v_210 | ~v_397 | ~v_396 | ~v_395 | ~v_394 | ~v_615 | ~v_614 | ~v_613 | ~v_612 | ~v_205 | ~v_204 | ~v_203 | ~v_202 | v_678;
assign x_30338 = v_677 | v_154;
assign x_30339 = v_677 | v_48;
assign x_30340 = v_676 | v_154;
assign x_30341 = v_676 | v_5;
assign x_30342 = v_675 | ~v_154;
assign x_30343 = v_675 | v_33;
assign x_30344 = v_674 | ~v_154;
assign x_30345 = v_674 | v_1;
assign x_30346 = v_673 | ~v_662;
assign x_30347 = v_673 | ~v_667;
assign x_30348 = v_673 | ~v_672;
assign x_30349 = v_101 | v_100 | v_93 | v_102 | v_172 | v_171 | v_170 | v_150 | v_149 | v_148 | v_147 | v_184 | ~v_389 | ~v_388 | ~v_671 | ~v_670 | ~v_387 | ~v_386 | ~v_653 | ~v_652 | ~v_669 | ~v_668 | ~v_289 | ~v_286 | ~v_649 | ~v_648 | ~v_647 | ~v_646 | ~v_383 | ~v_382 | ~v_381 | ~v_380 | ~v_279 | ~v_276 | ~v_379 | ~v_378 | ~v_645 | ~v_644 | ~v_643 | ~v_642 | ~v_271 | ~v_270 | ~v_269 | ~v_268 | v_672;
assign x_30350 = v_671 | v_173;
assign x_30351 = v_671 | v_132;
assign x_30352 = v_670 | ~v_173;
assign x_30353 = v_670 | v_117;
assign x_30354 = v_669 | v_174;
assign x_30355 = v_669 | v_6;
assign x_30356 = v_668 | ~v_174;
assign x_30357 = v_668 | v_3;
assign x_30358 = v_51 | v_60 | v_59 | v_58 | v_144 | v_145 | v_143 | v_142 | v_168 | v_167 | v_166 | v_183 | ~v_374 | ~v_373 | ~v_666 | ~v_665 | ~v_372 | ~v_371 | ~v_638 | ~v_637 | ~v_664 | ~v_663 | ~v_256 | ~v_253 | ~v_634 | ~v_633 | ~v_632 | ~v_631 | ~v_368 | ~v_367 | ~v_366 | ~v_365 | ~v_246 | ~v_243 | ~v_364 | ~v_363 | ~v_630 | ~v_629 | ~v_628 | ~v_627 | ~v_238 | ~v_237 | ~v_236 | ~v_235 | v_667;
assign x_30359 = v_666 | v_173;
assign x_30360 = v_666 | v_90;
assign x_30361 = v_665 | ~v_173;
assign x_30362 = v_665 | v_75;
assign x_30363 = v_664 | v_174;
assign x_30364 = v_664 | v_4;
assign x_30365 = v_663 | ~v_174;
assign x_30366 = v_663 | v_2;
assign x_30367 = v_17 | v_16 | v_8 | v_15 | v_136 | v_135 | v_134 | v_137 | v_164 | v_163 | v_162 | v_182 | ~v_359 | ~v_358 | ~v_661 | ~v_660 | ~v_357 | ~v_356 | ~v_623 | ~v_622 | ~v_659 | ~v_658 | ~v_223 | ~v_220 | ~v_619 | ~v_618 | ~v_617 | ~v_616 | ~v_353 | ~v_352 | ~v_351 | ~v_350 | ~v_213 | ~v_210 | ~v_349 | ~v_348 | ~v_615 | ~v_614 | ~v_613 | ~v_612 | ~v_205 | ~v_204 | ~v_203 | ~v_202 | v_662;
assign x_30368 = v_661 | v_173;
assign x_30369 = v_661 | v_48;
assign x_30370 = v_660 | ~v_173;
assign x_30371 = v_660 | v_33;
assign x_30372 = v_659 | v_174;
assign x_30373 = v_659 | v_5;
assign x_30374 = v_658 | ~v_174;
assign x_30375 = v_658 | v_1;
assign x_30376 = v_657 | ~v_626;
assign x_30377 = v_657 | ~v_641;
assign x_30378 = v_657 | ~v_656;
assign x_30379 = v_103 | v_97 | v_100 | v_93 | v_151 | v_171 | v_170 | v_160 | v_150 | v_148 | v_147 | v_184 | ~v_655 | ~v_654 | ~v_297 | ~v_296 | ~v_653 | ~v_652 | ~v_651 | ~v_650 | ~v_289 | ~v_286 | ~v_649 | ~v_648 | ~v_647 | ~v_646 | ~v_285 | ~v_284 | ~v_283 | ~v_282 | ~v_279 | ~v_276 | ~v_275 | ~v_274 | ~v_273 | ~v_272 | ~v_645 | ~v_644 | ~v_643 | ~v_642 | ~v_271 | ~v_270 | ~v_269 | ~v_268 | v_656;
assign x_30380 = v_655 | v_178;
assign x_30381 = v_655 | v_132;
assign x_30382 = v_654 | ~v_178;
assign x_30383 = v_654 | v_117;
assign x_30384 = v_653 | v_154;
assign x_30385 = v_653 | v_129;
assign x_30386 = v_652 | ~v_154;
assign x_30387 = v_652 | v_114;
assign x_30388 = v_651 | v_177;
assign x_30389 = v_651 | v_6;
assign x_30390 = v_650 | ~v_177;
assign x_30391 = v_650 | v_3;
assign x_30392 = v_649 | v_154;
assign x_30393 = v_649 | v_127;
assign x_30394 = v_648 | v_154;
assign x_30395 = v_648 | v_121;
assign x_30396 = v_647 | ~v_154;
assign x_30397 = v_647 | v_112;
assign x_30398 = v_646 | ~v_154;
assign x_30399 = v_646 | v_106;
assign x_30400 = v_645 | v_177;
assign x_30401 = v_645 | v_128;
assign x_30402 = v_644 | v_178;
assign x_30403 = v_644 | v_125;
assign x_30404 = v_643 | ~v_177;
assign x_30405 = v_643 | v_113;
assign x_30406 = v_642 | ~v_178;
assign x_30407 = v_642 | v_110;
assign x_30408 = v_55 | v_61 | v_51 | v_58 | v_159 | v_145 | v_143 | v_142 | v_167 | v_166 | v_146 | v_183 | ~v_640 | ~v_639 | ~v_264 | ~v_263 | ~v_638 | ~v_637 | ~v_636 | ~v_635 | ~v_256 | ~v_253 | ~v_634 | ~v_633 | ~v_632 | ~v_631 | ~v_252 | ~v_251 | ~v_250 | ~v_249 | ~v_246 | ~v_243 | ~v_242 | ~v_241 | ~v_240 | ~v_239 | ~v_630 | ~v_629 | ~v_628 | ~v_627 | ~v_238 | ~v_237 | ~v_236 | ~v_235 | v_641;
assign x_30409 = v_640 | v_178;
assign x_30410 = v_640 | v_90;
assign x_30411 = v_639 | ~v_178;
assign x_30412 = v_639 | v_75;
assign x_30413 = v_638 | v_154;
assign x_30414 = v_638 | v_87;
assign x_30415 = v_637 | ~v_154;
assign x_30416 = v_637 | v_72;
assign x_30417 = v_636 | v_177;
assign x_30418 = v_636 | v_4;
assign x_30419 = v_635 | ~v_177;
assign x_30420 = v_635 | v_2;
assign x_30421 = v_634 | v_154;
assign x_30422 = v_634 | v_85;
assign x_30423 = v_633 | v_154;
assign x_30424 = v_633 | v_79;
assign x_30425 = v_632 | ~v_154;
assign x_30426 = v_632 | v_70;
assign x_30427 = v_631 | ~v_154;
assign x_30428 = v_631 | v_64;
assign x_30429 = v_630 | v_177;
assign x_30430 = v_630 | v_86;
assign x_30431 = v_629 | v_178;
assign x_30432 = v_629 | v_83;
assign x_30433 = v_628 | ~v_177;
assign x_30434 = v_628 | v_71;
assign x_30435 = v_627 | ~v_178;
assign x_30436 = v_627 | v_68;
assign x_30437 = v_18 | v_8 | v_15 | v_12 | v_135 | v_134 | v_137 | v_138 | v_163 | v_162 | v_155 | v_182 | ~v_625 | ~v_624 | ~v_231 | ~v_230 | ~v_623 | ~v_622 | ~v_621 | ~v_620 | ~v_223 | ~v_220 | ~v_619 | ~v_618 | ~v_617 | ~v_616 | ~v_219 | ~v_218 | ~v_217 | ~v_216 | ~v_213 | ~v_210 | ~v_209 | ~v_208 | ~v_207 | ~v_206 | ~v_615 | ~v_614 | ~v_613 | ~v_612 | ~v_205 | ~v_204 | ~v_203 | ~v_202 | v_626;
assign x_30438 = v_625 | v_178;
assign x_30439 = v_625 | v_48;
assign x_30440 = v_624 | ~v_178;
assign x_30441 = v_624 | v_33;
assign x_30442 = v_623 | v_154;
assign x_30443 = v_623 | v_45;
assign x_30444 = v_622 | ~v_154;
assign x_30445 = v_622 | v_30;
assign x_30446 = v_621 | v_177;
assign x_30447 = v_621 | v_5;
assign x_30448 = v_620 | ~v_177;
assign x_30449 = v_620 | v_1;
assign x_30450 = v_619 | v_154;
assign x_30451 = v_619 | v_43;
assign x_30452 = v_618 | v_154;
assign x_30453 = v_618 | v_37;
assign x_30454 = v_617 | ~v_154;
assign x_30455 = v_617 | v_28;
assign x_30456 = v_616 | ~v_154;
assign x_30457 = v_616 | v_22;
assign x_30458 = v_615 | v_177;
assign x_30459 = v_615 | v_44;
assign x_30460 = v_614 | v_178;
assign x_30461 = v_614 | v_41;
assign x_30462 = v_613 | ~v_177;
assign x_30463 = v_613 | v_29;
assign x_30464 = v_612 | ~v_178;
assign x_30465 = v_612 | v_26;
assign x_30466 = v_611 | ~v_600;
assign x_30467 = v_611 | ~v_605;
assign x_30468 = v_611 | ~v_610;
assign x_30469 = v_98 | v_103 | v_101 | v_96 | v_100 | v_102 | v_170 | v_169 | v_150 | v_149 | v_147 | v_184 | ~v_609 | ~v_608 | ~v_299 | ~v_298 | ~v_435 | ~v_434 | ~v_607 | ~v_606 | ~v_291 | ~v_290 | ~v_289 | ~v_288 | ~v_287 | ~v_286 | ~v_431 | ~v_430 | ~v_429 | ~v_428 | ~v_281 | ~v_280 | ~v_279 | ~v_278 | ~v_277 | ~v_276 | ~v_427 | ~v_426 | ~v_425 | ~v_424 | ~v_271 | ~v_270 | ~v_269 | ~v_268 | v_610;
assign x_30470 = v_609 | v_153;
assign x_30471 = v_609 | v_132;
assign x_30472 = v_608 | ~v_153;
assign x_30473 = v_608 | v_117;
assign x_30474 = v_607 | v_152;
assign x_30475 = v_607 | v_6;
assign x_30476 = v_606 | ~v_152;
assign x_30477 = v_606 | v_3;
assign x_30478 = v_54 | v_56 | v_61 | v_60 | v_59 | v_58 | v_144 | v_145 | v_142 | v_166 | v_165 | v_183 | ~v_604 | ~v_603 | ~v_266 | ~v_265 | ~v_420 | ~v_419 | ~v_602 | ~v_601 | ~v_258 | ~v_257 | ~v_256 | ~v_255 | ~v_254 | ~v_253 | ~v_416 | ~v_415 | ~v_414 | ~v_413 | ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_244 | ~v_243 | ~v_412 | ~v_411 | ~v_410 | ~v_409 | ~v_238 | ~v_237 | ~v_236 | ~v_235 | v_605;
assign x_30479 = v_604 | v_153;
assign x_30480 = v_604 | v_90;
assign x_30481 = v_603 | ~v_153;
assign x_30482 = v_603 | v_75;
assign x_30483 = v_602 | v_152;
assign x_30484 = v_602 | v_4;
assign x_30485 = v_601 | ~v_152;
assign x_30486 = v_601 | v_2;
assign x_30487 = v_13 | v_18 | v_17 | v_16 | v_15 | v_11 | v_136 | v_134 | v_137 | v_162 | v_161 | v_182 | ~v_599 | ~v_598 | ~v_233 | ~v_232 | ~v_405 | ~v_404 | ~v_597 | ~v_596 | ~v_225 | ~v_224 | ~v_223 | ~v_222 | ~v_221 | ~v_220 | ~v_401 | ~v_400 | ~v_399 | ~v_398 | ~v_215 | ~v_214 | ~v_213 | ~v_212 | ~v_211 | ~v_210 | ~v_397 | ~v_396 | ~v_395 | ~v_394 | ~v_205 | ~v_204 | ~v_203 | ~v_202 | v_600;
assign x_30488 = v_599 | v_153;
assign x_30489 = v_599 | v_48;
assign x_30490 = v_598 | ~v_153;
assign x_30491 = v_598 | v_33;
assign x_30492 = v_597 | v_152;
assign x_30493 = v_597 | v_5;
assign x_30494 = v_596 | ~v_152;
assign x_30495 = v_596 | v_1;
assign x_30496 = v_595 | ~v_584;
assign x_30497 = v_595 | ~v_589;
assign x_30498 = v_595 | ~v_594;
assign x_30499 = v_101 | v_100 | v_99 | v_102 | v_172 | v_171 | v_170 | v_169 | v_149 | v_148 | v_147 | v_184 | ~v_483 | ~v_482 | ~v_593 | ~v_592 | ~v_545 | ~v_591 | ~v_590 | ~v_544 | ~v_477 | ~v_476 | ~v_289 | ~v_475 | ~v_474 | ~v_286 | ~v_539 | ~v_538 | ~v_537 | ~v_536 | ~v_473 | ~v_472 | ~v_279 | ~v_471 | ~v_470 | ~v_276 | ~v_535 | ~v_534 | ~v_533 | ~v_532 | ~v_271 | ~v_270 | ~v_269 | ~v_268 | v_594;
assign x_30500 = v_593 | v_139;
assign x_30501 = v_593 | v_132;
assign x_30502 = v_592 | v_140;
assign x_30503 = v_592 | v_6;
assign x_30504 = v_591 | ~v_139;
assign x_30505 = v_591 | v_117;
assign x_30506 = v_590 | ~v_140;
assign x_30507 = v_590 | v_3;
assign x_30508 = v_60 | v_59 | v_58 | v_57 | v_144 | v_143 | v_142 | v_168 | v_167 | v_166 | v_165 | v_183 | ~v_468 | ~v_467 | ~v_588 | ~v_587 | ~v_530 | ~v_586 | ~v_585 | ~v_529 | ~v_462 | ~v_461 | ~v_256 | ~v_460 | ~v_459 | ~v_253 | ~v_524 | ~v_523 | ~v_522 | ~v_521 | ~v_458 | ~v_457 | ~v_246 | ~v_456 | ~v_455 | ~v_243 | ~v_520 | ~v_519 | ~v_518 | ~v_517 | ~v_238 | ~v_237 | ~v_236 | ~v_235 | v_589;
assign x_30509 = v_588 | v_139;
assign x_30510 = v_588 | v_90;
assign x_30511 = v_587 | v_140;
assign x_30512 = v_587 | v_4;
assign x_30513 = v_586 | ~v_139;
assign x_30514 = v_586 | v_75;
assign x_30515 = v_585 | ~v_140;
assign x_30516 = v_585 | v_2;
assign x_30517 = v_17 | v_16 | v_15 | v_14 | ~v_453 | ~v_452 | v_136 | v_135 | v_134 | v_164 | v_163 | v_162 | v_161 | v_182 | ~v_583 | ~v_582 | ~v_515 | ~v_581 | ~v_580 | ~v_514 | ~v_447 | ~v_446 | ~v_223 | ~v_445 | ~v_444 | ~v_220 | ~v_509 | ~v_508 | ~v_507 | ~v_506 | ~v_443 | ~v_442 | ~v_213 | ~v_441 | ~v_440 | ~v_210 | ~v_505 | ~v_504 | ~v_503 | ~v_502 | ~v_205 | ~v_204 | ~v_203 | ~v_202 | v_584;
assign x_30518 = v_583 | v_139;
assign x_30519 = v_583 | v_48;
assign x_30520 = v_582 | v_140;
assign x_30521 = v_582 | v_5;
assign x_30522 = v_581 | ~v_139;
assign x_30523 = v_581 | v_33;
assign x_30524 = v_580 | ~v_140;
assign x_30525 = v_580 | v_1;
assign x_30526 = v_579 | ~v_568;
assign x_30527 = v_579 | ~v_573;
assign x_30528 = v_579 | ~v_578;
assign x_30529 = v_103 | v_101 | v_96 | v_100 | v_151 | v_171 | v_170 | v_169 | v_150 | v_149 | v_147 | v_184 | ~v_577 | ~v_576 | ~v_545 | ~v_544 | ~v_575 | ~v_574 | ~v_435 | ~v_434 | ~v_289 | ~v_286 | ~v_431 | ~v_430 | ~v_429 | ~v_428 | ~v_539 | ~v_538 | ~v_537 | ~v_536 | ~v_279 | ~v_276 | ~v_427 | ~v_426 | ~v_425 | ~v_424 | ~v_535 | ~v_534 | ~v_533 | ~v_532 | ~v_271 | ~v_270 | ~v_269 | ~v_268 | v_578;
assign x_30530 = v_577 | v_174;
assign x_30531 = v_577 | v_132;
assign x_30532 = v_576 | ~v_174;
assign x_30533 = v_576 | v_117;
assign x_30534 = v_575 | v_173;
assign x_30535 = v_575 | v_6;
assign x_30536 = v_574 | ~v_173;
assign x_30537 = v_574 | v_3;
assign x_30538 = v_54 | v_61 | v_59 | v_58 | v_144 | v_145 | v_142 | v_167 | v_166 | v_165 | v_146 | v_183 | ~v_572 | ~v_571 | ~v_530 | ~v_529 | ~v_570 | ~v_569 | ~v_420 | ~v_419 | ~v_256 | ~v_253 | ~v_416 | ~v_415 | ~v_414 | ~v_413 | ~v_524 | ~v_523 | ~v_522 | ~v_521 | ~v_246 | ~v_243 | ~v_412 | ~v_411 | ~v_410 | ~v_409 | ~v_520 | ~v_519 | ~v_518 | ~v_517 | ~v_238 | ~v_237 | ~v_236 | ~v_235 | v_573;
assign x_30539 = v_572 | v_174;
assign x_30540 = v_572 | v_90;
assign x_30541 = v_571 | ~v_174;
assign x_30542 = v_571 | v_75;
assign x_30543 = v_570 | v_173;
assign x_30544 = v_570 | v_4;
assign x_30545 = v_569 | ~v_173;
assign x_30546 = v_569 | v_2;
assign x_30547 = v_18 | v_16 | v_15 | v_11 | v_136 | v_134 | v_137 | v_138 | v_163 | v_162 | v_161 | v_182 | ~v_567 | ~v_566 | ~v_515 | ~v_514 | ~v_565 | ~v_564 | ~v_405 | ~v_404 | ~v_223 | ~v_220 | ~v_401 | ~v_400 | ~v_399 | ~v_398 | ~v_509 | ~v_508 | ~v_507 | ~v_506 | ~v_213 | ~v_210 | ~v_397 | ~v_396 | ~v_395 | ~v_394 | ~v_505 | ~v_504 | ~v_503 | ~v_502 | ~v_205 | ~v_204 | ~v_203 | ~v_202 | v_568;
assign x_30548 = v_567 | v_174;
assign x_30549 = v_567 | v_48;
assign x_30550 = v_566 | ~v_174;
assign x_30551 = v_566 | v_33;
assign x_30552 = v_565 | v_173;
assign x_30553 = v_565 | v_5;
assign x_30554 = v_564 | ~v_173;
assign x_30555 = v_564 | v_1;
assign x_30556 = v_563 | ~v_552;
assign x_30557 = v_563 | ~v_557;
assign x_30558 = v_563 | ~v_562;
assign x_30559 = v_103 | v_101 | v_100 | v_95 | v_102 | v_171 | v_170 | v_169 | v_150 | v_149 | v_148 | v_184 | ~v_389 | ~v_388 | ~v_545 | ~v_544 | ~v_561 | ~v_560 | ~v_559 | ~v_558 | ~v_387 | ~v_386 | ~v_289 | ~v_286 | ~v_383 | ~v_382 | ~v_381 | ~v_380 | ~v_539 | ~v_538 | ~v_537 | ~v_536 | ~v_279 | ~v_276 | ~v_379 | ~v_378 | ~v_535 | ~v_534 | ~v_533 | ~v_532 | ~v_271 | ~v_270 | ~v_269 | ~v_268 | v_562;
assign x_30560 = v_561 | v_141;
assign x_30561 = v_561 | v_132;
assign x_30562 = v_560 | v_141;
assign x_30563 = v_560 | v_6;
assign x_30564 = v_559 | ~v_141;
assign x_30565 = v_559 | v_117;
assign x_30566 = v_558 | ~v_141;
assign x_30567 = v_558 | v_3;
assign x_30568 = v_53 | v_61 | v_60 | v_59 | v_58 | v_144 | v_145 | v_143 | v_167 | v_166 | v_165 | v_183 | ~v_374 | ~v_373 | ~v_530 | ~v_529 | ~v_556 | ~v_555 | ~v_554 | ~v_553 | ~v_372 | ~v_371 | ~v_256 | ~v_253 | ~v_368 | ~v_367 | ~v_366 | ~v_365 | ~v_524 | ~v_523 | ~v_522 | ~v_521 | ~v_246 | ~v_243 | ~v_364 | ~v_363 | ~v_520 | ~v_519 | ~v_518 | ~v_517 | ~v_238 | ~v_237 | ~v_236 | ~v_235 | v_557;
assign x_30569 = v_556 | v_141;
assign x_30570 = v_556 | v_90;
assign x_30571 = v_555 | v_141;
assign x_30572 = v_555 | v_4;
assign x_30573 = v_554 | ~v_141;
assign x_30574 = v_554 | v_75;
assign x_30575 = v_553 | ~v_141;
assign x_30576 = v_553 | v_2;
assign x_30577 = v_18 | v_17 | v_16 | v_15 | v_10 | v_136 | v_135 | v_137 | v_163 | v_162 | v_161 | v_182 | ~v_359 | ~v_358 | ~v_515 | ~v_514 | ~v_551 | ~v_550 | ~v_549 | ~v_548 | ~v_357 | ~v_356 | ~v_223 | ~v_220 | ~v_353 | ~v_352 | ~v_351 | ~v_350 | ~v_509 | ~v_508 | ~v_507 | ~v_506 | ~v_213 | ~v_210 | ~v_349 | ~v_348 | ~v_505 | ~v_504 | ~v_503 | ~v_502 | ~v_205 | ~v_204 | ~v_203 | ~v_202 | v_552;
assign x_30578 = v_551 | v_141;
assign x_30579 = v_551 | v_48;
assign x_30580 = v_550 | v_141;
assign x_30581 = v_550 | v_5;
assign x_30582 = v_549 | ~v_141;
assign x_30583 = v_549 | v_33;
assign x_30584 = v_548 | ~v_141;
assign x_30585 = v_548 | v_1;
assign x_30586 = v_547 | ~v_516;
assign x_30587 = v_547 | ~v_531;
assign x_30588 = v_547 | ~v_546;
assign x_30589 = v_103 | v_97 | v_100 | v_102 | v_171 | v_170 | v_169 | v_160 | v_150 | v_148 | v_147 | v_184 | ~v_545 | ~v_544 | ~v_543 | ~v_542 | ~v_541 | ~v_540 | ~v_297 | ~v_296 | ~v_289 | ~v_286 | ~v_285 | ~v_284 | ~v_283 | ~v_282 | ~v_539 | ~v_538 | ~v_537 | ~v_536 | ~v_279 | ~v_276 | ~v_275 | ~v_274 | ~v_273 | ~v_272 | ~v_535 | ~v_534 | ~v_533 | ~v_532 | ~v_271 | ~v_270 | ~v_269 | ~v_268 | v_546;
assign x_30590 = v_545 | v_141;
assign x_30591 = v_545 | v_129;
assign x_30592 = v_544 | ~v_141;
assign x_30593 = v_544 | v_114;
assign x_30594 = v_543 | v_176;
assign x_30595 = v_543 | v_132;
assign x_30596 = v_542 | v_175;
assign x_30597 = v_542 | v_6;
assign x_30598 = v_541 | ~v_176;
assign x_30599 = v_541 | v_117;
assign x_30600 = v_540 | ~v_175;
assign x_30601 = v_540 | v_3;
assign x_30602 = v_539 | v_173;
assign x_30603 = v_539 | v_127;
assign x_30604 = v_538 | v_174;
assign x_30605 = v_538 | v_121;
assign x_30606 = v_537 | ~v_173;
assign x_30607 = v_537 | v_112;
assign x_30608 = v_536 | ~v_174;
assign x_30609 = v_536 | v_106;
assign x_30610 = v_535 | v_175;
assign x_30611 = v_535 | v_128;
assign x_30612 = v_534 | v_176;
assign x_30613 = v_534 | v_125;
assign x_30614 = v_533 | ~v_175;
assign x_30615 = v_533 | v_113;
assign x_30616 = v_532 | ~v_176;
assign x_30617 = v_532 | v_110;
assign x_30618 = v_55 | v_61 | v_60 | v_58 | v_159 | v_145 | v_143 | v_142 | v_167 | v_166 | v_165 | v_183 | ~v_530 | ~v_529 | ~v_528 | ~v_527 | ~v_526 | ~v_525 | ~v_264 | ~v_263 | ~v_256 | ~v_253 | ~v_252 | ~v_251 | ~v_250 | ~v_249 | ~v_524 | ~v_523 | ~v_522 | ~v_521 | ~v_246 | ~v_243 | ~v_242 | ~v_241 | ~v_240 | ~v_239 | ~v_520 | ~v_519 | ~v_518 | ~v_517 | ~v_238 | ~v_237 | ~v_236 | ~v_235 | v_531;
assign x_30619 = v_530 | v_141;
assign x_30620 = v_530 | v_87;
assign x_30621 = v_529 | ~v_141;
assign x_30622 = v_529 | v_72;
assign x_30623 = v_528 | v_176;
assign x_30624 = v_528 | v_90;
assign x_30625 = v_527 | v_175;
assign x_30626 = v_527 | v_4;
assign x_30627 = v_526 | ~v_176;
assign x_30628 = v_526 | v_75;
assign x_30629 = v_525 | ~v_175;
assign x_30630 = v_525 | v_2;
assign x_30631 = v_524 | v_173;
assign x_30632 = v_524 | v_85;
assign x_30633 = v_523 | v_174;
assign x_30634 = v_523 | v_79;
assign x_30635 = v_522 | ~v_173;
assign x_30636 = v_522 | v_70;
assign x_30637 = v_521 | ~v_174;
assign x_30638 = v_521 | v_64;
assign x_30639 = v_520 | v_175;
assign x_30640 = v_520 | v_86;
assign x_30641 = v_519 | v_176;
assign x_30642 = v_519 | v_83;
assign x_30643 = v_518 | ~v_175;
assign x_30644 = v_518 | v_71;
assign x_30645 = v_517 | ~v_176;
assign x_30646 = v_517 | v_68;
assign x_30647 = v_18 | v_17 | v_15 | v_12 | v_135 | v_134 | v_137 | v_163 | v_162 | v_161 | v_155 | v_182 | ~v_515 | ~v_514 | ~v_513 | ~v_512 | ~v_511 | ~v_510 | ~v_231 | ~v_230 | ~v_223 | ~v_220 | ~v_219 | ~v_218 | ~v_217 | ~v_216 | ~v_509 | ~v_508 | ~v_507 | ~v_506 | ~v_213 | ~v_210 | ~v_209 | ~v_208 | ~v_207 | ~v_206 | ~v_505 | ~v_504 | ~v_503 | ~v_502 | ~v_205 | ~v_204 | ~v_203 | ~v_202 | v_516;
assign x_30648 = v_515 | v_141;
assign x_30649 = v_515 | v_45;
assign x_30650 = v_514 | ~v_141;
assign x_30651 = v_514 | v_30;
assign x_30652 = v_513 | v_176;
assign x_30653 = v_513 | v_48;
assign x_30654 = v_512 | v_175;
assign x_30655 = v_512 | v_5;
assign x_30656 = v_511 | ~v_176;
assign x_30657 = v_511 | v_33;
assign x_30658 = v_510 | ~v_175;
assign x_30659 = v_510 | v_1;
assign x_30660 = v_509 | v_173;
assign x_30661 = v_509 | v_43;
assign x_30662 = v_508 | v_174;
assign x_30663 = v_508 | v_37;
assign x_30664 = v_507 | ~v_173;
assign x_30665 = v_507 | v_28;
assign x_30666 = v_506 | ~v_174;
assign x_30667 = v_506 | v_22;
assign x_30668 = v_505 | v_175;
assign x_30669 = v_505 | v_44;
assign x_30670 = v_504 | v_176;
assign x_30671 = v_504 | v_41;
assign x_30672 = v_503 | ~v_175;
assign x_30673 = v_503 | v_29;
assign x_30674 = v_502 | ~v_176;
assign x_30675 = v_502 | v_26;
assign x_30676 = v_501 | ~v_490;
assign x_30677 = v_501 | ~v_495;
assign x_30678 = v_501 | ~v_500;
assign x_30679 = v_98 | v_103 | v_101 | v_100 | v_151 | v_170 | v_169 | v_150 | v_149 | v_148 | v_147 | v_184 | ~v_389 | ~v_388 | ~v_299 | ~v_298 | ~v_387 | ~v_386 | ~v_499 | ~v_498 | ~v_497 | ~v_496 | ~v_291 | ~v_290 | ~v_289 | ~v_288 | ~v_287 | ~v_286 | ~v_383 | ~v_382 | ~v_381 | ~v_380 | ~v_281 | ~v_280 | ~v_279 | ~v_278 | ~v_277 | ~v_276 | ~v_379 | ~v_378 | ~v_271 | ~v_270 | ~v_269 | ~v_268 | v_500;
assign x_30680 = v_499 | v_140;
assign x_30681 = v_499 | v_132;
assign x_30682 = v_498 | v_139;
assign x_30683 = v_498 | v_6;
assign x_30684 = v_497 | ~v_140;
assign x_30685 = v_497 | v_117;
assign x_30686 = v_496 | ~v_139;
assign x_30687 = v_496 | v_3;
assign x_30688 = v_56 | v_61 | v_59 | v_58 | v_144 | v_145 | v_143 | v_142 | v_166 | v_165 | v_146 | v_183 | ~v_374 | ~v_373 | ~v_266 | ~v_265 | ~v_372 | ~v_371 | ~v_494 | ~v_493 | ~v_492 | ~v_491 | ~v_258 | ~v_257 | ~v_256 | ~v_255 | ~v_254 | ~v_253 | ~v_368 | ~v_367 | ~v_366 | ~v_365 | ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_244 | ~v_243 | ~v_364 | ~v_363 | ~v_238 | ~v_237 | ~v_236 | ~v_235 | v_495;
assign x_30689 = v_494 | v_140;
assign x_30690 = v_494 | v_90;
assign x_30691 = v_493 | v_139;
assign x_30692 = v_493 | v_4;
assign x_30693 = v_492 | ~v_140;
assign x_30694 = v_492 | v_75;
assign x_30695 = v_491 | ~v_139;
assign x_30696 = v_491 | v_2;
assign x_30697 = v_13 | v_18 | v_16 | v_15 | v_136 | v_135 | v_134 | v_137 | v_138 | v_162 | v_161 | v_182 | ~v_359 | ~v_358 | ~v_233 | ~v_232 | ~v_357 | ~v_356 | ~v_489 | ~v_488 | ~v_487 | ~v_486 | ~v_225 | ~v_224 | ~v_223 | ~v_222 | ~v_221 | ~v_220 | ~v_353 | ~v_352 | ~v_351 | ~v_350 | ~v_215 | ~v_214 | ~v_213 | ~v_212 | ~v_211 | ~v_210 | ~v_349 | ~v_348 | ~v_205 | ~v_204 | ~v_203 | ~v_202 | v_490;
assign x_30698 = v_489 | v_140;
assign x_30699 = v_489 | v_48;
assign x_30700 = v_488 | v_139;
assign x_30701 = v_488 | v_5;
assign x_30702 = v_487 | ~v_140;
assign x_30703 = v_487 | v_33;
assign x_30704 = v_486 | ~v_139;
assign x_30705 = v_486 | v_1;
assign x_30706 = v_485 | ~v_454;
assign x_30707 = v_485 | ~v_469;
assign x_30708 = v_485 | ~v_484;
assign x_30709 = v_103 | v_101 | v_94 | v_99 | v_102 | v_171 | v_169 | v_149 | v_148 | v_147 | v_184 | v_181 | ~v_483 | ~v_482 | ~v_481 | ~v_480 | ~v_345 | ~v_479 | ~v_478 | ~v_344 | ~v_477 | ~v_476 | ~v_289 | ~v_475 | ~v_474 | ~v_286 | ~v_339 | ~v_338 | ~v_337 | ~v_336 | ~v_473 | ~v_472 | ~v_279 | ~v_471 | ~v_470 | ~v_276 | ~v_335 | ~v_334 | ~v_333 | ~v_332 | ~v_271 | ~v_270 | ~v_269 | ~v_268 | v_484;
assign x_30710 = v_483 | v_133;
assign x_30711 = v_483 | v_19;
assign x_30712 = v_482 | v_118;
assign x_30713 = v_482 | ~v_19;
assign x_30714 = v_481 | v_156;
assign x_30715 = v_481 | v_132;
assign x_30716 = v_480 | v_157;
assign x_30717 = v_480 | v_6;
assign x_30718 = v_479 | ~v_156;
assign x_30719 = v_479 | v_117;
assign x_30720 = v_478 | ~v_157;
assign x_30721 = v_478 | v_3;
assign x_30722 = v_477 | v_152;
assign x_30723 = v_477 | v_130;
assign x_30724 = v_476 | v_153;
assign x_30725 = v_476 | v_122;
assign x_30726 = v_475 | ~v_152;
assign x_30727 = v_475 | v_115;
assign x_30728 = v_474 | ~v_153;
assign x_30729 = v_474 | v_107;
assign x_30730 = v_473 | v_156;
assign x_30731 = v_473 | v_131;
assign x_30732 = v_472 | v_157;
assign x_30733 = v_472 | v_126;
assign x_30734 = v_471 | ~v_156;
assign x_30735 = v_471 | v_116;
assign x_30736 = v_470 | ~v_157;
assign x_30737 = v_470 | v_111;
assign x_30738 = v_61 | v_52 | v_60 | v_59 | v_57 | v_144 | v_180 | v_143 | v_142 | v_167 | v_165 | v_183 | ~v_468 | ~v_467 | ~v_466 | ~v_465 | ~v_330 | ~v_464 | ~v_463 | ~v_329 | ~v_462 | ~v_461 | ~v_256 | ~v_460 | ~v_459 | ~v_253 | ~v_324 | ~v_323 | ~v_322 | ~v_321 | ~v_458 | ~v_457 | ~v_246 | ~v_456 | ~v_455 | ~v_243 | ~v_320 | ~v_319 | ~v_318 | ~v_317 | ~v_238 | ~v_237 | ~v_236 | ~v_235 | v_469;
assign x_30739 = v_468 | v_91;
assign x_30740 = v_468 | v_19;
assign x_30741 = v_467 | v_76;
assign x_30742 = v_467 | ~v_19;
assign x_30743 = v_466 | v_156;
assign x_30744 = v_466 | v_90;
assign x_30745 = v_465 | v_157;
assign x_30746 = v_465 | v_4;
assign x_30747 = v_464 | ~v_156;
assign x_30748 = v_464 | v_75;
assign x_30749 = v_463 | ~v_157;
assign x_30750 = v_463 | v_2;
assign x_30751 = v_462 | v_152;
assign x_30752 = v_462 | v_88;
assign x_30753 = v_461 | v_153;
assign x_30754 = v_461 | v_80;
assign x_30755 = v_460 | ~v_152;
assign x_30756 = v_460 | v_73;
assign x_30757 = v_459 | ~v_153;
assign x_30758 = v_459 | v_65;
assign x_30759 = v_458 | v_156;
assign x_30760 = v_458 | v_89;
assign x_30761 = v_457 | v_157;
assign x_30762 = v_457 | v_84;
assign x_30763 = v_456 | ~v_156;
assign x_30764 = v_456 | v_74;
assign x_30765 = v_455 | ~v_157;
assign x_30766 = v_455 | v_69;
assign x_30767 = v_9 | v_18 | v_17 | v_16 | v_14 | ~v_453 | ~v_452 | v_136 | v_135 | v_134 | v_179 | v_163 | v_161 | v_182 | ~v_451 | ~v_450 | ~v_315 | ~v_449 | ~v_448 | ~v_314 | ~v_447 | ~v_446 | ~v_223 | ~v_445 | ~v_444 | ~v_220 | ~v_309 | ~v_308 | ~v_307 | ~v_306 | ~v_443 | ~v_442 | ~v_213 | ~v_441 | ~v_440 | ~v_210 | ~v_305 | ~v_304 | ~v_303 | ~v_302 | ~v_205 | ~v_204 | ~v_203 | ~v_202 | v_454;
assign x_30768 = v_453 | v_49;
assign x_30769 = v_453 | v_19;
assign x_30770 = v_452 | v_34;
assign x_30771 = v_452 | ~v_19;
assign x_30772 = v_451 | v_156;
assign x_30773 = v_451 | v_48;
assign x_30774 = v_450 | v_157;
assign x_30775 = v_450 | v_5;
assign x_30776 = v_449 | ~v_156;
assign x_30777 = v_449 | v_33;
assign x_30778 = v_448 | ~v_157;
assign x_30779 = v_448 | v_1;
assign x_30780 = v_447 | v_152;
assign x_30781 = v_447 | v_46;
assign x_30782 = v_446 | v_153;
assign x_30783 = v_446 | v_38;
assign x_30784 = v_445 | ~v_152;
assign x_30785 = v_445 | v_31;
assign x_30786 = v_444 | ~v_153;
assign x_30787 = v_444 | v_23;
assign x_30788 = v_443 | v_156;
assign x_30789 = v_443 | v_47;
assign x_30790 = v_442 | v_157;
assign x_30791 = v_442 | v_42;
assign x_30792 = v_441 | ~v_156;
assign x_30793 = v_441 | v_32;
assign x_30794 = v_440 | ~v_157;
assign x_30795 = v_440 | v_27;
assign x_30796 = v_439 | ~v_408;
assign x_30797 = v_439 | ~v_423;
assign x_30798 = v_439 | ~v_438;
assign x_30799 = v_101 | v_96 | v_94 | v_102 | v_172 | v_171 | v_169 | v_150 | v_149 | v_147 | v_184 | v_181 | ~v_437 | ~v_436 | ~v_435 | ~v_434 | ~v_345 | ~v_344 | ~v_433 | ~v_432 | ~v_289 | ~v_286 | ~v_431 | ~v_430 | ~v_429 | ~v_428 | ~v_339 | ~v_338 | ~v_337 | ~v_336 | ~v_279 | ~v_276 | ~v_335 | ~v_334 | ~v_333 | ~v_332 | ~v_427 | ~v_426 | ~v_425 | ~v_424 | ~v_271 | ~v_270 | ~v_269 | ~v_268 | v_438;
assign x_30800 = v_437 | v_177;
assign x_30801 = v_437 | v_132;
assign x_30802 = v_436 | ~v_177;
assign x_30803 = v_436 | v_117;
assign x_30804 = v_435 | v_154;
assign x_30805 = v_435 | v_133;
assign x_30806 = v_434 | ~v_154;
assign x_30807 = v_434 | v_118;
assign x_30808 = v_433 | v_178;
assign x_30809 = v_433 | v_6;
assign x_30810 = v_432 | ~v_178;
assign x_30811 = v_432 | v_3;
assign x_30812 = v_431 | v_154;
assign x_30813 = v_431 | v_130;
assign x_30814 = v_430 | v_154;
assign x_30815 = v_430 | v_122;
assign x_30816 = v_429 | ~v_154;
assign x_30817 = v_429 | v_115;
assign x_30818 = v_428 | ~v_154;
assign x_30819 = v_428 | v_107;
assign x_30820 = v_427 | v_177;
assign x_30821 = v_427 | v_131;
assign x_30822 = v_426 | v_178;
assign x_30823 = v_426 | v_126;
assign x_30824 = v_425 | ~v_177;
assign x_30825 = v_425 | v_116;
assign x_30826 = v_424 | ~v_178;
assign x_30827 = v_424 | v_111;
assign x_30828 = v_54 | v_52 | v_60 | v_59 | v_144 | v_180 | v_145 | v_142 | v_168 | v_167 | v_165 | v_183 | ~v_422 | ~v_421 | ~v_420 | ~v_419 | ~v_330 | ~v_329 | ~v_418 | ~v_417 | ~v_256 | ~v_253 | ~v_416 | ~v_415 | ~v_414 | ~v_413 | ~v_324 | ~v_323 | ~v_322 | ~v_321 | ~v_246 | ~v_243 | ~v_320 | ~v_319 | ~v_318 | ~v_317 | ~v_412 | ~v_411 | ~v_410 | ~v_409 | ~v_238 | ~v_237 | ~v_236 | ~v_235 | v_423;
assign x_30829 = v_422 | v_177;
assign x_30830 = v_422 | v_90;
assign x_30831 = v_421 | ~v_177;
assign x_30832 = v_421 | v_75;
assign x_30833 = v_420 | v_154;
assign x_30834 = v_420 | v_91;
assign x_30835 = v_419 | ~v_154;
assign x_30836 = v_419 | v_76;
assign x_30837 = v_418 | v_178;
assign x_30838 = v_418 | v_4;
assign x_30839 = v_417 | ~v_178;
assign x_30840 = v_417 | v_2;
assign x_30841 = v_416 | v_154;
assign x_30842 = v_416 | v_88;
assign x_30843 = v_415 | v_154;
assign x_30844 = v_415 | v_80;
assign x_30845 = v_414 | ~v_154;
assign x_30846 = v_414 | v_73;
assign x_30847 = v_413 | ~v_154;
assign x_30848 = v_413 | v_65;
assign x_30849 = v_412 | v_177;
assign x_30850 = v_412 | v_89;
assign x_30851 = v_411 | v_178;
assign x_30852 = v_411 | v_84;
assign x_30853 = v_410 | ~v_177;
assign x_30854 = v_410 | v_74;
assign x_30855 = v_409 | ~v_178;
assign x_30856 = v_409 | v_69;
assign x_30857 = v_9 | v_17 | v_16 | v_11 | v_136 | v_134 | v_137 | v_179 | v_164 | v_163 | v_161 | v_182 | ~v_407 | ~v_406 | ~v_405 | ~v_404 | ~v_315 | ~v_314 | ~v_403 | ~v_402 | ~v_223 | ~v_220 | ~v_401 | ~v_400 | ~v_399 | ~v_398 | ~v_309 | ~v_308 | ~v_307 | ~v_306 | ~v_213 | ~v_210 | ~v_305 | ~v_304 | ~v_303 | ~v_302 | ~v_397 | ~v_396 | ~v_395 | ~v_394 | ~v_205 | ~v_204 | ~v_203 | ~v_202 | v_408;
assign x_30858 = v_407 | v_177;
assign x_30859 = v_407 | v_48;
assign x_30860 = v_406 | ~v_177;
assign x_30861 = v_406 | v_33;
assign x_30862 = v_405 | v_154;
assign x_30863 = v_405 | v_49;
assign x_30864 = v_404 | ~v_154;
assign x_30865 = v_404 | v_34;
assign x_30866 = v_403 | v_178;
assign x_30867 = v_403 | v_5;
assign x_30868 = v_402 | ~v_178;
assign x_30869 = v_402 | v_1;
assign x_30870 = v_401 | v_154;
assign x_30871 = v_401 | v_46;
assign x_30872 = v_400 | v_154;
assign x_30873 = v_400 | v_38;
assign x_30874 = v_399 | ~v_154;
assign x_30875 = v_399 | v_31;
assign x_30876 = v_398 | ~v_154;
assign x_30877 = v_398 | v_23;
assign x_30878 = v_397 | v_177;
assign x_30879 = v_397 | v_47;
assign x_30880 = v_396 | v_178;
assign x_30881 = v_396 | v_42;
assign x_30882 = v_395 | ~v_177;
assign x_30883 = v_395 | v_32;
assign x_30884 = v_394 | ~v_178;
assign x_30885 = v_394 | v_27;
assign x_30886 = v_393 | ~v_362;
assign x_30887 = v_393 | ~v_377;
assign x_30888 = v_393 | ~v_392;
assign x_30889 = v_103 | v_101 | v_94 | v_102 | v_171 | v_169 | v_150 | v_149 | v_148 | v_147 | v_184 | v_181 | ~v_391 | ~v_390 | ~v_389 | ~v_388 | ~v_387 | ~v_386 | ~v_345 | ~v_344 | ~v_385 | ~v_384 | ~v_289 | ~v_286 | ~v_383 | ~v_382 | ~v_381 | ~v_380 | ~v_339 | ~v_338 | ~v_337 | ~v_336 | ~v_279 | ~v_276 | ~v_335 | ~v_334 | ~v_333 | ~v_332 | ~v_379 | ~v_378 | ~v_271 | ~v_270 | ~v_269 | ~v_268 | v_392;
assign x_30890 = v_391 | v_175;
assign x_30891 = v_391 | v_132;
assign x_30892 = v_390 | ~v_175;
assign x_30893 = v_390 | v_117;
assign x_30894 = v_389 | v_175;
assign x_30895 = v_389 | v_131;
assign x_30896 = v_388 | ~v_175;
assign x_30897 = v_388 | v_116;
assign x_30898 = v_387 | v_141;
assign x_30899 = v_387 | v_133;
assign x_30900 = v_386 | ~v_141;
assign x_30901 = v_386 | v_118;
assign x_30902 = v_385 | v_176;
assign x_30903 = v_385 | v_6;
assign x_30904 = v_384 | ~v_176;
assign x_30905 = v_384 | v_3;
assign x_30906 = v_383 | v_173;
assign x_30907 = v_383 | v_130;
assign x_30908 = v_382 | v_174;
assign x_30909 = v_382 | v_122;
assign x_30910 = v_381 | ~v_173;
assign x_30911 = v_381 | v_115;
assign x_30912 = v_380 | ~v_174;
assign x_30913 = v_380 | v_107;
assign x_30914 = v_379 | v_176;
assign x_30915 = v_379 | v_126;
assign x_30916 = v_378 | ~v_176;
assign x_30917 = v_378 | v_111;
assign x_30918 = v_61 | v_52 | v_60 | v_59 | v_144 | v_180 | v_145 | v_143 | v_142 | v_167 | v_165 | v_183 | ~v_376 | ~v_375 | ~v_374 | ~v_373 | ~v_372 | ~v_371 | ~v_330 | ~v_329 | ~v_370 | ~v_369 | ~v_256 | ~v_253 | ~v_368 | ~v_367 | ~v_366 | ~v_365 | ~v_324 | ~v_323 | ~v_322 | ~v_321 | ~v_246 | ~v_243 | ~v_320 | ~v_319 | ~v_318 | ~v_317 | ~v_364 | ~v_363 | ~v_238 | ~v_237 | ~v_236 | ~v_235 | v_377;
assign x_30919 = v_376 | v_175;
assign x_30920 = v_376 | v_90;
assign x_30921 = v_375 | ~v_175;
assign x_30922 = v_375 | v_75;
assign x_30923 = v_374 | v_175;
assign x_30924 = v_374 | v_89;
assign x_30925 = v_373 | ~v_175;
assign x_30926 = v_373 | v_74;
assign x_30927 = v_372 | v_141;
assign x_30928 = v_372 | v_91;
assign x_30929 = v_371 | ~v_141;
assign x_30930 = v_371 | v_76;
assign x_30931 = v_370 | v_176;
assign x_30932 = v_370 | v_4;
assign x_30933 = v_369 | ~v_176;
assign x_30934 = v_369 | v_2;
assign x_30935 = v_368 | v_173;
assign x_30936 = v_368 | v_88;
assign x_30937 = v_367 | v_174;
assign x_30938 = v_367 | v_80;
assign x_30939 = v_366 | ~v_173;
assign x_30940 = v_366 | v_73;
assign x_30941 = v_365 | ~v_174;
assign x_30942 = v_365 | v_65;
assign x_30943 = v_364 | v_176;
assign x_30944 = v_364 | v_84;
assign x_30945 = v_363 | ~v_176;
assign x_30946 = v_363 | v_69;
assign x_30947 = v_9 | v_18 | v_17 | v_16 | v_136 | v_135 | v_134 | v_137 | v_179 | v_163 | v_161 | v_182 | ~v_361 | ~v_360 | ~v_359 | ~v_358 | ~v_357 | ~v_356 | ~v_315 | ~v_314 | ~v_355 | ~v_354 | ~v_223 | ~v_220 | ~v_353 | ~v_352 | ~v_351 | ~v_350 | ~v_309 | ~v_308 | ~v_307 | ~v_306 | ~v_213 | ~v_210 | ~v_305 | ~v_304 | ~v_303 | ~v_302 | ~v_349 | ~v_348 | ~v_205 | ~v_204 | ~v_203 | ~v_202 | v_362;
assign x_30948 = v_361 | v_175;
assign x_30949 = v_361 | v_48;
assign x_30950 = v_360 | ~v_175;
assign x_30951 = v_360 | v_33;
assign x_30952 = v_359 | v_175;
assign x_30953 = v_359 | v_47;
assign x_30954 = v_358 | ~v_175;
assign x_30955 = v_358 | v_32;
assign x_30956 = v_357 | v_141;
assign x_30957 = v_357 | v_49;
assign x_30958 = v_356 | ~v_141;
assign x_30959 = v_356 | v_34;
assign x_30960 = v_355 | v_176;
assign x_30961 = v_355 | v_5;
assign x_30962 = v_354 | ~v_176;
assign x_30963 = v_354 | v_1;
assign x_30964 = v_353 | v_173;
assign x_30965 = v_353 | v_46;
assign x_30966 = v_352 | v_174;
assign x_30967 = v_352 | v_38;
assign x_30968 = v_351 | ~v_173;
assign x_30969 = v_351 | v_31;
assign x_30970 = v_350 | ~v_174;
assign x_30971 = v_350 | v_23;
assign x_30972 = v_349 | v_176;
assign x_30973 = v_349 | v_42;
assign x_30974 = v_348 | ~v_176;
assign x_30975 = v_348 | v_27;
assign x_30976 = v_347 | ~v_316;
assign x_30977 = v_347 | ~v_331;
assign x_30978 = v_347 | ~v_346;
assign x_30979 = v_103 | v_97 | v_95 | v_94 | v_102 | v_171 | v_169 | v_160 | v_150 | v_148 | v_184 | v_181 | ~v_297 | ~v_296 | ~v_345 | ~v_344 | ~v_343 | ~v_342 | ~v_341 | ~v_340 | ~v_289 | ~v_286 | ~v_285 | ~v_284 | ~v_283 | ~v_282 | ~v_339 | ~v_338 | ~v_337 | ~v_336 | ~v_279 | ~v_276 | ~v_335 | ~v_334 | ~v_333 | ~v_332 | ~v_275 | ~v_274 | ~v_273 | ~v_272 | ~v_271 | ~v_270 | ~v_269 | ~v_268 | v_346;
assign x_30980 = v_345 | v_158;
assign x_30981 = v_345 | v_129;
assign x_30982 = v_344 | ~v_158;
assign x_30983 = v_344 | v_114;
assign x_30984 = v_343 | v_158;
assign x_30985 = v_343 | v_132;
assign x_30986 = v_342 | v_158;
assign x_30987 = v_342 | v_6;
assign x_30988 = v_341 | ~v_158;
assign x_30989 = v_341 | v_117;
assign x_30990 = v_340 | ~v_158;
assign x_30991 = v_340 | v_3;
assign x_30992 = v_339 | v_178;
assign x_30993 = v_339 | v_127;
assign x_30994 = v_338 | v_177;
assign x_30995 = v_338 | v_121;
assign x_30996 = v_337 | ~v_178;
assign x_30997 = v_337 | v_112;
assign x_30998 = v_336 | ~v_177;
assign x_30999 = v_336 | v_106;
assign x_31000 = v_335 | v_158;
assign x_31001 = v_335 | v_128;
assign x_31002 = v_334 | v_158;
assign x_31003 = v_334 | v_125;
assign x_31004 = v_333 | ~v_158;
assign x_31005 = v_333 | v_113;
assign x_31006 = v_332 | ~v_158;
assign x_31007 = v_332 | v_110;
assign x_31008 = v_53 | v_55 | v_61 | v_52 | v_60 | v_180 | v_159 | v_145 | v_143 | v_167 | v_165 | v_183 | ~v_264 | ~v_263 | ~v_330 | ~v_329 | ~v_328 | ~v_327 | ~v_326 | ~v_325 | ~v_256 | ~v_253 | ~v_252 | ~v_251 | ~v_250 | ~v_249 | ~v_324 | ~v_323 | ~v_322 | ~v_321 | ~v_246 | ~v_243 | ~v_320 | ~v_319 | ~v_318 | ~v_317 | ~v_242 | ~v_241 | ~v_240 | ~v_239 | ~v_238 | ~v_237 | ~v_236 | ~v_235 | v_331;
assign x_31009 = v_330 | v_158;
assign x_31010 = v_330 | v_87;
assign x_31011 = v_329 | ~v_158;
assign x_31012 = v_329 | v_72;
assign x_31013 = v_328 | v_158;
assign x_31014 = v_328 | v_90;
assign x_31015 = v_327 | v_158;
assign x_31016 = v_327 | v_4;
assign x_31017 = v_326 | ~v_158;
assign x_31018 = v_326 | v_75;
assign x_31019 = v_325 | ~v_158;
assign x_31020 = v_325 | v_2;
assign x_31021 = v_324 | v_178;
assign x_31022 = v_324 | v_85;
assign x_31023 = v_323 | v_177;
assign x_31024 = v_323 | v_79;
assign x_31025 = v_322 | ~v_178;
assign x_31026 = v_322 | v_70;
assign x_31027 = v_321 | ~v_177;
assign x_31028 = v_321 | v_64;
assign x_31029 = v_320 | v_158;
assign x_31030 = v_320 | v_86;
assign x_31031 = v_319 | v_158;
assign x_31032 = v_319 | v_83;
assign x_31033 = v_318 | ~v_158;
assign x_31034 = v_318 | v_71;
assign x_31035 = v_317 | ~v_158;
assign x_31036 = v_317 | v_68;
assign x_31037 = v_9 | v_18 | v_17 | v_12 | v_10 | v_135 | v_137 | v_179 | v_163 | v_161 | v_155 | v_182 | ~v_231 | ~v_230 | ~v_315 | ~v_314 | ~v_313 | ~v_312 | ~v_311 | ~v_310 | ~v_223 | ~v_220 | ~v_219 | ~v_218 | ~v_217 | ~v_216 | ~v_309 | ~v_308 | ~v_307 | ~v_306 | ~v_213 | ~v_210 | ~v_305 | ~v_304 | ~v_303 | ~v_302 | ~v_209 | ~v_208 | ~v_207 | ~v_206 | ~v_205 | ~v_204 | ~v_203 | ~v_202 | v_316;
assign x_31038 = v_315 | v_158;
assign x_31039 = v_315 | v_45;
assign x_31040 = v_314 | ~v_158;
assign x_31041 = v_314 | v_30;
assign x_31042 = v_313 | v_158;
assign x_31043 = v_313 | v_48;
assign x_31044 = v_312 | v_158;
assign x_31045 = v_312 | v_5;
assign x_31046 = v_311 | ~v_158;
assign x_31047 = v_311 | v_33;
assign x_31048 = v_310 | ~v_158;
assign x_31049 = v_310 | v_1;
assign x_31050 = v_309 | v_178;
assign x_31051 = v_309 | v_43;
assign x_31052 = v_308 | v_177;
assign x_31053 = v_308 | v_37;
assign x_31054 = v_307 | ~v_178;
assign x_31055 = v_307 | v_28;
assign x_31056 = v_306 | ~v_177;
assign x_31057 = v_306 | v_22;
assign x_31058 = v_305 | v_158;
assign x_31059 = v_305 | v_44;
assign x_31060 = v_304 | v_158;
assign x_31061 = v_304 | v_41;
assign x_31062 = v_303 | ~v_158;
assign x_31063 = v_303 | v_29;
assign x_31064 = v_302 | ~v_158;
assign x_31065 = v_302 | v_26;
assign x_31066 = v_301 | ~v_234;
assign x_31067 = v_301 | ~v_267;
assign x_31068 = v_301 | ~v_300;
assign x_31069 = v_98 | v_103 | v_97 | v_100 | v_102 | v_170 | v_169 | v_160 | v_150 | v_148 | v_147 | v_184 | ~v_299 | ~v_298 | ~v_297 | ~v_296 | ~v_295 | ~v_294 | ~v_293 | ~v_292 | ~v_291 | ~v_290 | ~v_289 | ~v_288 | ~v_287 | ~v_286 | ~v_285 | ~v_284 | ~v_283 | ~v_282 | ~v_281 | ~v_280 | ~v_279 | ~v_278 | ~v_277 | ~v_276 | ~v_275 | ~v_274 | ~v_273 | ~v_272 | ~v_271 | ~v_270 | ~v_269 | ~v_268 | v_300;
assign x_31070 = v_299 | v_129;
assign x_31071 = v_299 | v_19;
assign x_31072 = v_298 | v_114;
assign x_31073 = v_298 | ~v_19;
assign x_31074 = v_297 | v_158;
assign x_31075 = v_297 | v_133;
assign x_31076 = v_296 | ~v_158;
assign x_31077 = v_296 | v_118;
assign x_31078 = v_295 | v_157;
assign x_31079 = v_295 | v_132;
assign x_31080 = v_294 | v_156;
assign x_31081 = v_294 | v_6;
assign x_31082 = v_293 | ~v_157;
assign x_31083 = v_293 | v_117;
assign x_31084 = v_292 | ~v_156;
assign x_31085 = v_292 | v_3;
assign x_31086 = v_291 | v_152;
assign x_31087 = v_291 | v_127;
assign x_31088 = v_290 | v_153;
assign x_31089 = v_290 | v_121;
assign x_31090 = v_289 | v_154;
assign x_31091 = v_289 | v_119;
assign x_31092 = v_288 | ~v_152;
assign x_31093 = v_288 | v_112;
assign x_31094 = v_287 | ~v_153;
assign x_31095 = v_287 | v_106;
assign x_31096 = v_286 | ~v_154;
assign x_31097 = v_286 | v_104;
assign x_31098 = v_285 | v_178;
assign x_31099 = v_285 | v_130;
assign x_31100 = v_284 | v_177;
assign x_31101 = v_284 | v_122;
assign x_31102 = v_283 | ~v_178;
assign x_31103 = v_283 | v_115;
assign x_31104 = v_282 | ~v_177;
assign x_31105 = v_282 | v_107;
assign x_31106 = v_281 | v_156;
assign x_31107 = v_281 | v_128;
assign x_31108 = v_280 | v_157;
assign x_31109 = v_280 | v_125;
assign x_31110 = v_279 | v_158;
assign x_31111 = v_279 | v_124;
assign x_31112 = v_278 | ~v_156;
assign x_31113 = v_278 | v_113;
assign x_31114 = v_277 | ~v_157;
assign x_31115 = v_277 | v_110;
assign x_31116 = v_276 | ~v_158;
assign x_31117 = v_276 | v_109;
assign x_31118 = v_275 | v_158;
assign x_31119 = v_275 | v_131;
assign x_31120 = v_274 | v_158;
assign x_31121 = v_274 | v_126;
assign x_31122 = v_273 | ~v_158;
assign x_31123 = v_273 | v_116;
assign x_31124 = v_272 | ~v_158;
assign x_31125 = v_272 | v_111;
assign x_31126 = v_271 | v_178;
assign x_31127 = v_271 | v_123;
assign x_31128 = v_270 | v_177;
assign x_31129 = v_270 | v_120;
assign x_31130 = v_269 | ~v_178;
assign x_31131 = v_269 | v_108;
assign x_31132 = v_268 | ~v_177;
assign x_31133 = v_268 | v_105;
assign x_31134 = v_56 | v_55 | v_61 | v_60 | v_58 | v_159 | v_145 | v_143 | v_142 | v_166 | v_165 | v_183 | ~v_266 | ~v_265 | ~v_264 | ~v_263 | ~v_262 | ~v_261 | ~v_260 | ~v_259 | ~v_258 | ~v_257 | ~v_256 | ~v_255 | ~v_254 | ~v_253 | ~v_252 | ~v_251 | ~v_250 | ~v_249 | ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_244 | ~v_243 | ~v_242 | ~v_241 | ~v_240 | ~v_239 | ~v_238 | ~v_237 | ~v_236 | ~v_235 | v_267;
assign x_31135 = v_266 | v_87;
assign x_31136 = v_266 | v_19;
assign x_31137 = v_265 | v_72;
assign x_31138 = v_265 | ~v_19;
assign x_31139 = v_264 | v_158;
assign x_31140 = v_264 | v_91;
assign x_31141 = v_263 | ~v_158;
assign x_31142 = v_263 | v_76;
assign x_31143 = v_262 | v_157;
assign x_31144 = v_262 | v_90;
assign x_31145 = v_261 | v_156;
assign x_31146 = v_261 | v_4;
assign x_31147 = v_260 | ~v_157;
assign x_31148 = v_260 | v_75;
assign x_31149 = v_259 | ~v_156;
assign x_31150 = v_259 | v_2;
assign x_31151 = v_258 | v_152;
assign x_31152 = v_258 | v_85;
assign x_31153 = v_257 | v_153;
assign x_31154 = v_257 | v_79;
assign x_31155 = v_256 | v_154;
assign x_31156 = v_256 | v_77;
assign x_31157 = v_255 | ~v_152;
assign x_31158 = v_255 | v_70;
assign x_31159 = v_254 | ~v_153;
assign x_31160 = v_254 | v_64;
assign x_31161 = v_253 | ~v_154;
assign x_31162 = v_253 | v_62;
assign x_31163 = v_252 | v_178;
assign x_31164 = v_252 | v_88;
assign x_31165 = v_251 | v_177;
assign x_31166 = v_251 | v_80;
assign x_31167 = v_250 | ~v_178;
assign x_31168 = v_250 | v_73;
assign x_31169 = v_249 | ~v_177;
assign x_31170 = v_249 | v_65;
assign x_31171 = v_248 | v_156;
assign x_31172 = v_248 | v_86;
assign x_31173 = v_247 | v_157;
assign x_31174 = v_247 | v_83;
assign x_31175 = v_246 | v_158;
assign x_31176 = v_246 | v_82;
assign x_31177 = v_245 | ~v_156;
assign x_31178 = v_245 | v_71;
assign x_31179 = v_244 | ~v_157;
assign x_31180 = v_244 | v_68;
assign x_31181 = v_243 | ~v_158;
assign x_31182 = v_243 | v_67;
assign x_31183 = v_242 | v_158;
assign x_31184 = v_242 | v_89;
assign x_31185 = v_241 | v_158;
assign x_31186 = v_241 | v_84;
assign x_31187 = v_240 | ~v_158;
assign x_31188 = v_240 | v_74;
assign x_31189 = v_239 | ~v_158;
assign x_31190 = v_239 | v_69;
assign x_31191 = v_238 | v_178;
assign x_31192 = v_238 | v_81;
assign x_31193 = v_237 | v_177;
assign x_31194 = v_237 | v_78;
assign x_31195 = v_236 | ~v_178;
assign x_31196 = v_236 | v_66;
assign x_31197 = v_235 | ~v_177;
assign x_31198 = v_235 | v_63;
assign x_31199 = v_13 | v_18 | v_17 | v_15 | v_12 | v_135 | v_134 | v_137 | v_162 | v_161 | v_155 | v_182 | ~v_233 | ~v_232 | ~v_231 | ~v_230 | ~v_229 | ~v_228 | ~v_227 | ~v_226 | ~v_225 | ~v_224 | ~v_223 | ~v_222 | ~v_221 | ~v_220 | ~v_219 | ~v_218 | ~v_217 | ~v_216 | ~v_215 | ~v_214 | ~v_213 | ~v_212 | ~v_211 | ~v_210 | ~v_209 | ~v_208 | ~v_207 | ~v_206 | ~v_205 | ~v_204 | ~v_203 | ~v_202 | v_234;
assign x_31200 = v_233 | v_45;
assign x_31201 = v_233 | v_19;
assign x_31202 = v_232 | v_30;
assign x_31203 = v_232 | ~v_19;
assign x_31204 = v_231 | v_158;
assign x_31205 = v_231 | v_49;
assign x_31206 = v_230 | ~v_158;
assign x_31207 = v_230 | v_34;
assign x_31208 = v_229 | v_157;
assign x_31209 = v_229 | v_48;
assign x_31210 = v_228 | v_156;
assign x_31211 = v_228 | v_5;
assign x_31212 = v_227 | ~v_157;
assign x_31213 = v_227 | v_33;
assign x_31214 = v_226 | ~v_156;
assign x_31215 = v_226 | v_1;
assign x_31216 = v_225 | v_152;
assign x_31217 = v_225 | v_43;
assign x_31218 = v_224 | v_153;
assign x_31219 = v_224 | v_37;
assign x_31220 = v_223 | v_154;
assign x_31221 = v_223 | v_35;
assign x_31222 = v_222 | ~v_152;
assign x_31223 = v_222 | v_28;
assign x_31224 = v_221 | ~v_153;
assign x_31225 = v_221 | v_22;
assign x_31226 = v_220 | ~v_154;
assign x_31227 = v_220 | v_20;
assign x_31228 = v_219 | v_178;
assign x_31229 = v_219 | v_46;
assign x_31230 = v_218 | v_177;
assign x_31231 = v_218 | v_38;
assign x_31232 = v_217 | ~v_178;
assign x_31233 = v_217 | v_31;
assign x_31234 = v_216 | ~v_177;
assign x_31235 = v_216 | v_23;
assign x_31236 = v_215 | v_156;
assign x_31237 = v_215 | v_44;
assign x_31238 = v_214 | v_157;
assign x_31239 = v_214 | v_41;
assign x_31240 = v_213 | v_158;
assign x_31241 = v_213 | v_40;
assign x_31242 = v_212 | ~v_156;
assign x_31243 = v_212 | v_29;
assign x_31244 = v_211 | ~v_157;
assign x_31245 = v_211 | v_26;
assign x_31246 = v_210 | ~v_158;
assign x_31247 = v_210 | v_25;
assign x_31248 = v_209 | v_158;
assign x_31249 = v_209 | v_47;
assign x_31250 = v_208 | v_158;
assign x_31251 = v_208 | v_42;
assign x_31252 = v_207 | ~v_158;
assign x_31253 = v_207 | v_32;
assign x_31254 = v_206 | ~v_158;
assign x_31255 = v_206 | v_27;
assign x_31256 = v_205 | v_178;
assign x_31257 = v_205 | v_39;
assign x_31258 = v_204 | v_177;
assign x_31259 = v_204 | v_36;
assign x_31260 = v_203 | ~v_178;
assign x_31261 = v_203 | v_24;
assign x_31262 = v_202 | ~v_177;
assign x_31263 = v_202 | v_21;
assign x_31264 = v_201 | ~v_192;
assign x_31265 = v_201 | ~v_198;
assign x_31266 = v_201 | ~v_199;
assign x_31267 = v_201 | ~v_200;
assign x_31268 = v_201 | ~v_178;
assign x_31269 = v_201 | ~v_177;
assign x_31270 = ~v_193 | ~v_185 | v_200;
assign x_31271 = ~v_189 | ~v_195 | v_199;
assign x_31272 = ~v_193 | ~v_197 | v_198;
assign x_31273 = v_197 | ~v_194;
assign x_31274 = v_197 | ~v_196;
assign x_31275 = v_197 | ~v_157;
assign x_31276 = v_197 | ~v_156;
assign x_31277 = ~v_186 | ~v_195 | v_196;
assign x_31278 = v_195 | ~v_176;
assign x_31279 = v_195 | ~v_175;
assign x_31280 = ~v_188 | ~v_193 | v_194;
assign x_31281 = v_193 | ~v_153;
assign x_31282 = v_193 | ~v_152;
assign x_31283 = ~v_189 | ~v_191 | v_192;
assign x_31284 = v_191 | ~v_187;
assign x_31285 = v_191 | ~v_190;
assign x_31286 = v_191 | ~v_176;
assign x_31287 = v_191 | ~v_175;
assign x_31288 = ~v_189 | ~v_188 | v_190;
assign x_31289 = v_189 | ~v_174;
assign x_31290 = v_189 | ~v_173;
assign x_31291 = v_188 | ~v_178;
assign x_31292 = v_188 | ~v_177;
assign x_31293 = ~v_186 | ~v_185 | v_187;
assign x_31294 = v_186 | ~v_140;
assign x_31295 = v_186 | ~v_139;
assign x_31296 = v_185 | ~v_157;
assign x_31297 = v_185 | ~v_156;
assign x_31298 = x_2 & x_3;
assign x_31299 = x_1 & x_31298;
assign x_31300 = x_4 & x_5;
assign x_31301 = x_6 & x_7;
assign x_31302 = x_31300 & x_31301;
assign x_31303 = x_31299 & x_31302;
assign x_31304 = x_8 & x_9;
assign x_31305 = x_10 & x_11;
assign x_31306 = x_31304 & x_31305;
assign x_31307 = x_12 & x_13;
assign x_31308 = x_14 & x_15;
assign x_31309 = x_31307 & x_31308;
assign x_31310 = x_31306 & x_31309;
assign x_31311 = x_31303 & x_31310;
assign x_31312 = x_17 & x_18;
assign x_31313 = x_16 & x_31312;
assign x_31314 = x_19 & x_20;
assign x_31315 = x_21 & x_22;
assign x_31316 = x_31314 & x_31315;
assign x_31317 = x_31313 & x_31316;
assign x_31318 = x_23 & x_24;
assign x_31319 = x_25 & x_26;
assign x_31320 = x_31318 & x_31319;
assign x_31321 = x_27 & x_28;
assign x_31322 = x_29 & x_30;
assign x_31323 = x_31321 & x_31322;
assign x_31324 = x_31320 & x_31323;
assign x_31325 = x_31317 & x_31324;
assign x_31326 = x_31311 & x_31325;
assign x_31327 = x_32 & x_33;
assign x_31328 = x_31 & x_31327;
assign x_31329 = x_34 & x_35;
assign x_31330 = x_36 & x_37;
assign x_31331 = x_31329 & x_31330;
assign x_31332 = x_31328 & x_31331;
assign x_31333 = x_38 & x_39;
assign x_31334 = x_40 & x_41;
assign x_31335 = x_31333 & x_31334;
assign x_31336 = x_42 & x_43;
assign x_31337 = x_44 & x_45;
assign x_31338 = x_31336 & x_31337;
assign x_31339 = x_31335 & x_31338;
assign x_31340 = x_31332 & x_31339;
assign x_31341 = x_46 & x_47;
assign x_31342 = x_48 & x_49;
assign x_31343 = x_31341 & x_31342;
assign x_31344 = x_50 & x_51;
assign x_31345 = x_52 & x_53;
assign x_31346 = x_31344 & x_31345;
assign x_31347 = x_31343 & x_31346;
assign x_31348 = x_54 & x_55;
assign x_31349 = x_56 & x_57;
assign x_31350 = x_31348 & x_31349;
assign x_31351 = x_58 & x_59;
assign x_31352 = x_60 & x_61;
assign x_31353 = x_31351 & x_31352;
assign x_31354 = x_31350 & x_31353;
assign x_31355 = x_31347 & x_31354;
assign x_31356 = x_31340 & x_31355;
assign x_31357 = x_31326 & x_31356;
assign x_31358 = x_63 & x_64;
assign x_31359 = x_62 & x_31358;
assign x_31360 = x_65 & x_66;
assign x_31361 = x_67 & x_68;
assign x_31362 = x_31360 & x_31361;
assign x_31363 = x_31359 & x_31362;
assign x_31364 = x_69 & x_70;
assign x_31365 = x_71 & x_72;
assign x_31366 = x_31364 & x_31365;
assign x_31367 = x_73 & x_74;
assign x_31368 = x_75 & x_76;
assign x_31369 = x_31367 & x_31368;
assign x_31370 = x_31366 & x_31369;
assign x_31371 = x_31363 & x_31370;
assign x_31372 = x_78 & x_79;
assign x_31373 = x_77 & x_31372;
assign x_31374 = x_80 & x_81;
assign x_31375 = x_82 & x_83;
assign x_31376 = x_31374 & x_31375;
assign x_31377 = x_31373 & x_31376;
assign x_31378 = x_84 & x_85;
assign x_31379 = x_86 & x_87;
assign x_31380 = x_31378 & x_31379;
assign x_31381 = x_88 & x_89;
assign x_31382 = x_90 & x_91;
assign x_31383 = x_31381 & x_31382;
assign x_31384 = x_31380 & x_31383;
assign x_31385 = x_31377 & x_31384;
assign x_31386 = x_31371 & x_31385;
assign x_31387 = x_93 & x_94;
assign x_31388 = x_92 & x_31387;
assign x_31389 = x_95 & x_96;
assign x_31390 = x_97 & x_98;
assign x_31391 = x_31389 & x_31390;
assign x_31392 = x_31388 & x_31391;
assign x_31393 = x_99 & x_100;
assign x_31394 = x_101 & x_102;
assign x_31395 = x_31393 & x_31394;
assign x_31396 = x_103 & x_104;
assign x_31397 = x_105 & x_106;
assign x_31398 = x_31396 & x_31397;
assign x_31399 = x_31395 & x_31398;
assign x_31400 = x_31392 & x_31399;
assign x_31401 = x_107 & x_108;
assign x_31402 = x_109 & x_110;
assign x_31403 = x_31401 & x_31402;
assign x_31404 = x_111 & x_112;
assign x_31405 = x_113 & x_114;
assign x_31406 = x_31404 & x_31405;
assign x_31407 = x_31403 & x_31406;
assign x_31408 = x_115 & x_116;
assign x_31409 = x_117 & x_118;
assign x_31410 = x_31408 & x_31409;
assign x_31411 = x_119 & x_120;
assign x_31412 = x_121 & x_122;
assign x_31413 = x_31411 & x_31412;
assign x_31414 = x_31410 & x_31413;
assign x_31415 = x_31407 & x_31414;
assign x_31416 = x_31400 & x_31415;
assign x_31417 = x_31386 & x_31416;
assign x_31418 = x_31357 & x_31417;
assign x_31419 = x_124 & x_125;
assign x_31420 = x_123 & x_31419;
assign x_31421 = x_126 & x_127;
assign x_31422 = x_128 & x_129;
assign x_31423 = x_31421 & x_31422;
assign x_31424 = x_31420 & x_31423;
assign x_31425 = x_130 & x_131;
assign x_31426 = x_132 & x_133;
assign x_31427 = x_31425 & x_31426;
assign x_31428 = x_134 & x_135;
assign x_31429 = x_136 & x_137;
assign x_31430 = x_31428 & x_31429;
assign x_31431 = x_31427 & x_31430;
assign x_31432 = x_31424 & x_31431;
assign x_31433 = x_139 & x_140;
assign x_31434 = x_138 & x_31433;
assign x_31435 = x_141 & x_142;
assign x_31436 = x_143 & x_144;
assign x_31437 = x_31435 & x_31436;
assign x_31438 = x_31434 & x_31437;
assign x_31439 = x_145 & x_146;
assign x_31440 = x_147 & x_148;
assign x_31441 = x_31439 & x_31440;
assign x_31442 = x_149 & x_150;
assign x_31443 = x_151 & x_152;
assign x_31444 = x_31442 & x_31443;
assign x_31445 = x_31441 & x_31444;
assign x_31446 = x_31438 & x_31445;
assign x_31447 = x_31432 & x_31446;
assign x_31448 = x_154 & x_155;
assign x_31449 = x_153 & x_31448;
assign x_31450 = x_156 & x_157;
assign x_31451 = x_158 & x_159;
assign x_31452 = x_31450 & x_31451;
assign x_31453 = x_31449 & x_31452;
assign x_31454 = x_160 & x_161;
assign x_31455 = x_162 & x_163;
assign x_31456 = x_31454 & x_31455;
assign x_31457 = x_164 & x_165;
assign x_31458 = x_166 & x_167;
assign x_31459 = x_31457 & x_31458;
assign x_31460 = x_31456 & x_31459;
assign x_31461 = x_31453 & x_31460;
assign x_31462 = x_168 & x_169;
assign x_31463 = x_170 & x_171;
assign x_31464 = x_31462 & x_31463;
assign x_31465 = x_172 & x_173;
assign x_31466 = x_174 & x_175;
assign x_31467 = x_31465 & x_31466;
assign x_31468 = x_31464 & x_31467;
assign x_31469 = x_176 & x_177;
assign x_31470 = x_178 & x_179;
assign x_31471 = x_31469 & x_31470;
assign x_31472 = x_180 & x_181;
assign x_31473 = x_182 & x_183;
assign x_31474 = x_31472 & x_31473;
assign x_31475 = x_31471 & x_31474;
assign x_31476 = x_31468 & x_31475;
assign x_31477 = x_31461 & x_31476;
assign x_31478 = x_31447 & x_31477;
assign x_31479 = x_185 & x_186;
assign x_31480 = x_184 & x_31479;
assign x_31481 = x_187 & x_188;
assign x_31482 = x_189 & x_190;
assign x_31483 = x_31481 & x_31482;
assign x_31484 = x_31480 & x_31483;
assign x_31485 = x_191 & x_192;
assign x_31486 = x_193 & x_194;
assign x_31487 = x_31485 & x_31486;
assign x_31488 = x_195 & x_196;
assign x_31489 = x_197 & x_198;
assign x_31490 = x_31488 & x_31489;
assign x_31491 = x_31487 & x_31490;
assign x_31492 = x_31484 & x_31491;
assign x_31493 = x_200 & x_201;
assign x_31494 = x_199 & x_31493;
assign x_31495 = x_202 & x_203;
assign x_31496 = x_204 & x_205;
assign x_31497 = x_31495 & x_31496;
assign x_31498 = x_31494 & x_31497;
assign x_31499 = x_206 & x_207;
assign x_31500 = x_208 & x_209;
assign x_31501 = x_31499 & x_31500;
assign x_31502 = x_210 & x_211;
assign x_31503 = x_212 & x_213;
assign x_31504 = x_31502 & x_31503;
assign x_31505 = x_31501 & x_31504;
assign x_31506 = x_31498 & x_31505;
assign x_31507 = x_31492 & x_31506;
assign x_31508 = x_215 & x_216;
assign x_31509 = x_214 & x_31508;
assign x_31510 = x_217 & x_218;
assign x_31511 = x_219 & x_220;
assign x_31512 = x_31510 & x_31511;
assign x_31513 = x_31509 & x_31512;
assign x_31514 = x_221 & x_222;
assign x_31515 = x_223 & x_224;
assign x_31516 = x_31514 & x_31515;
assign x_31517 = x_225 & x_226;
assign x_31518 = x_227 & x_228;
assign x_31519 = x_31517 & x_31518;
assign x_31520 = x_31516 & x_31519;
assign x_31521 = x_31513 & x_31520;
assign x_31522 = x_229 & x_230;
assign x_31523 = x_231 & x_232;
assign x_31524 = x_31522 & x_31523;
assign x_31525 = x_233 & x_234;
assign x_31526 = x_235 & x_236;
assign x_31527 = x_31525 & x_31526;
assign x_31528 = x_31524 & x_31527;
assign x_31529 = x_237 & x_238;
assign x_31530 = x_239 & x_240;
assign x_31531 = x_31529 & x_31530;
assign x_31532 = x_241 & x_242;
assign x_31533 = x_243 & x_244;
assign x_31534 = x_31532 & x_31533;
assign x_31535 = x_31531 & x_31534;
assign x_31536 = x_31528 & x_31535;
assign x_31537 = x_31521 & x_31536;
assign x_31538 = x_31507 & x_31537;
assign x_31539 = x_31478 & x_31538;
assign x_31540 = x_31418 & x_31539;
assign x_31541 = x_246 & x_247;
assign x_31542 = x_245 & x_31541;
assign x_31543 = x_248 & x_249;
assign x_31544 = x_250 & x_251;
assign x_31545 = x_31543 & x_31544;
assign x_31546 = x_31542 & x_31545;
assign x_31547 = x_252 & x_253;
assign x_31548 = x_254 & x_255;
assign x_31549 = x_31547 & x_31548;
assign x_31550 = x_256 & x_257;
assign x_31551 = x_258 & x_259;
assign x_31552 = x_31550 & x_31551;
assign x_31553 = x_31549 & x_31552;
assign x_31554 = x_31546 & x_31553;
assign x_31555 = x_261 & x_262;
assign x_31556 = x_260 & x_31555;
assign x_31557 = x_263 & x_264;
assign x_31558 = x_265 & x_266;
assign x_31559 = x_31557 & x_31558;
assign x_31560 = x_31556 & x_31559;
assign x_31561 = x_267 & x_268;
assign x_31562 = x_269 & x_270;
assign x_31563 = x_31561 & x_31562;
assign x_31564 = x_271 & x_272;
assign x_31565 = x_273 & x_274;
assign x_31566 = x_31564 & x_31565;
assign x_31567 = x_31563 & x_31566;
assign x_31568 = x_31560 & x_31567;
assign x_31569 = x_31554 & x_31568;
assign x_31570 = x_276 & x_277;
assign x_31571 = x_275 & x_31570;
assign x_31572 = x_278 & x_279;
assign x_31573 = x_280 & x_281;
assign x_31574 = x_31572 & x_31573;
assign x_31575 = x_31571 & x_31574;
assign x_31576 = x_282 & x_283;
assign x_31577 = x_284 & x_285;
assign x_31578 = x_31576 & x_31577;
assign x_31579 = x_286 & x_287;
assign x_31580 = x_288 & x_289;
assign x_31581 = x_31579 & x_31580;
assign x_31582 = x_31578 & x_31581;
assign x_31583 = x_31575 & x_31582;
assign x_31584 = x_290 & x_291;
assign x_31585 = x_292 & x_293;
assign x_31586 = x_31584 & x_31585;
assign x_31587 = x_294 & x_295;
assign x_31588 = x_296 & x_297;
assign x_31589 = x_31587 & x_31588;
assign x_31590 = x_31586 & x_31589;
assign x_31591 = x_298 & x_299;
assign x_31592 = x_300 & x_301;
assign x_31593 = x_31591 & x_31592;
assign x_31594 = x_302 & x_303;
assign x_31595 = x_304 & x_305;
assign x_31596 = x_31594 & x_31595;
assign x_31597 = x_31593 & x_31596;
assign x_31598 = x_31590 & x_31597;
assign x_31599 = x_31583 & x_31598;
assign x_31600 = x_31569 & x_31599;
assign x_31601 = x_307 & x_308;
assign x_31602 = x_306 & x_31601;
assign x_31603 = x_309 & x_310;
assign x_31604 = x_311 & x_312;
assign x_31605 = x_31603 & x_31604;
assign x_31606 = x_31602 & x_31605;
assign x_31607 = x_313 & x_314;
assign x_31608 = x_315 & x_316;
assign x_31609 = x_31607 & x_31608;
assign x_31610 = x_317 & x_318;
assign x_31611 = x_319 & x_320;
assign x_31612 = x_31610 & x_31611;
assign x_31613 = x_31609 & x_31612;
assign x_31614 = x_31606 & x_31613;
assign x_31615 = x_322 & x_323;
assign x_31616 = x_321 & x_31615;
assign x_31617 = x_324 & x_325;
assign x_31618 = x_326 & x_327;
assign x_31619 = x_31617 & x_31618;
assign x_31620 = x_31616 & x_31619;
assign x_31621 = x_328 & x_329;
assign x_31622 = x_330 & x_331;
assign x_31623 = x_31621 & x_31622;
assign x_31624 = x_332 & x_333;
assign x_31625 = x_334 & x_335;
assign x_31626 = x_31624 & x_31625;
assign x_31627 = x_31623 & x_31626;
assign x_31628 = x_31620 & x_31627;
assign x_31629 = x_31614 & x_31628;
assign x_31630 = x_337 & x_338;
assign x_31631 = x_336 & x_31630;
assign x_31632 = x_339 & x_340;
assign x_31633 = x_341 & x_342;
assign x_31634 = x_31632 & x_31633;
assign x_31635 = x_31631 & x_31634;
assign x_31636 = x_343 & x_344;
assign x_31637 = x_345 & x_346;
assign x_31638 = x_31636 & x_31637;
assign x_31639 = x_347 & x_348;
assign x_31640 = x_349 & x_350;
assign x_31641 = x_31639 & x_31640;
assign x_31642 = x_31638 & x_31641;
assign x_31643 = x_31635 & x_31642;
assign x_31644 = x_351 & x_352;
assign x_31645 = x_353 & x_354;
assign x_31646 = x_31644 & x_31645;
assign x_31647 = x_355 & x_356;
assign x_31648 = x_357 & x_358;
assign x_31649 = x_31647 & x_31648;
assign x_31650 = x_31646 & x_31649;
assign x_31651 = x_359 & x_360;
assign x_31652 = x_361 & x_362;
assign x_31653 = x_31651 & x_31652;
assign x_31654 = x_363 & x_364;
assign x_31655 = x_365 & x_366;
assign x_31656 = x_31654 & x_31655;
assign x_31657 = x_31653 & x_31656;
assign x_31658 = x_31650 & x_31657;
assign x_31659 = x_31643 & x_31658;
assign x_31660 = x_31629 & x_31659;
assign x_31661 = x_31600 & x_31660;
assign x_31662 = x_368 & x_369;
assign x_31663 = x_367 & x_31662;
assign x_31664 = x_370 & x_371;
assign x_31665 = x_372 & x_373;
assign x_31666 = x_31664 & x_31665;
assign x_31667 = x_31663 & x_31666;
assign x_31668 = x_374 & x_375;
assign x_31669 = x_376 & x_377;
assign x_31670 = x_31668 & x_31669;
assign x_31671 = x_378 & x_379;
assign x_31672 = x_380 & x_381;
assign x_31673 = x_31671 & x_31672;
assign x_31674 = x_31670 & x_31673;
assign x_31675 = x_31667 & x_31674;
assign x_31676 = x_383 & x_384;
assign x_31677 = x_382 & x_31676;
assign x_31678 = x_385 & x_386;
assign x_31679 = x_387 & x_388;
assign x_31680 = x_31678 & x_31679;
assign x_31681 = x_31677 & x_31680;
assign x_31682 = x_389 & x_390;
assign x_31683 = x_391 & x_392;
assign x_31684 = x_31682 & x_31683;
assign x_31685 = x_393 & x_394;
assign x_31686 = x_395 & x_396;
assign x_31687 = x_31685 & x_31686;
assign x_31688 = x_31684 & x_31687;
assign x_31689 = x_31681 & x_31688;
assign x_31690 = x_31675 & x_31689;
assign x_31691 = x_398 & x_399;
assign x_31692 = x_397 & x_31691;
assign x_31693 = x_400 & x_401;
assign x_31694 = x_402 & x_403;
assign x_31695 = x_31693 & x_31694;
assign x_31696 = x_31692 & x_31695;
assign x_31697 = x_404 & x_405;
assign x_31698 = x_406 & x_407;
assign x_31699 = x_31697 & x_31698;
assign x_31700 = x_408 & x_409;
assign x_31701 = x_410 & x_411;
assign x_31702 = x_31700 & x_31701;
assign x_31703 = x_31699 & x_31702;
assign x_31704 = x_31696 & x_31703;
assign x_31705 = x_412 & x_413;
assign x_31706 = x_414 & x_415;
assign x_31707 = x_31705 & x_31706;
assign x_31708 = x_416 & x_417;
assign x_31709 = x_418 & x_419;
assign x_31710 = x_31708 & x_31709;
assign x_31711 = x_31707 & x_31710;
assign x_31712 = x_420 & x_421;
assign x_31713 = x_422 & x_423;
assign x_31714 = x_31712 & x_31713;
assign x_31715 = x_424 & x_425;
assign x_31716 = x_426 & x_427;
assign x_31717 = x_31715 & x_31716;
assign x_31718 = x_31714 & x_31717;
assign x_31719 = x_31711 & x_31718;
assign x_31720 = x_31704 & x_31719;
assign x_31721 = x_31690 & x_31720;
assign x_31722 = x_429 & x_430;
assign x_31723 = x_428 & x_31722;
assign x_31724 = x_431 & x_432;
assign x_31725 = x_433 & x_434;
assign x_31726 = x_31724 & x_31725;
assign x_31727 = x_31723 & x_31726;
assign x_31728 = x_435 & x_436;
assign x_31729 = x_437 & x_438;
assign x_31730 = x_31728 & x_31729;
assign x_31731 = x_439 & x_440;
assign x_31732 = x_441 & x_442;
assign x_31733 = x_31731 & x_31732;
assign x_31734 = x_31730 & x_31733;
assign x_31735 = x_31727 & x_31734;
assign x_31736 = x_443 & x_444;
assign x_31737 = x_445 & x_446;
assign x_31738 = x_31736 & x_31737;
assign x_31739 = x_447 & x_448;
assign x_31740 = x_449 & x_450;
assign x_31741 = x_31739 & x_31740;
assign x_31742 = x_31738 & x_31741;
assign x_31743 = x_451 & x_452;
assign x_31744 = x_453 & x_454;
assign x_31745 = x_31743 & x_31744;
assign x_31746 = x_455 & x_456;
assign x_31747 = x_457 & x_458;
assign x_31748 = x_31746 & x_31747;
assign x_31749 = x_31745 & x_31748;
assign x_31750 = x_31742 & x_31749;
assign x_31751 = x_31735 & x_31750;
assign x_31752 = x_460 & x_461;
assign x_31753 = x_459 & x_31752;
assign x_31754 = x_462 & x_463;
assign x_31755 = x_464 & x_465;
assign x_31756 = x_31754 & x_31755;
assign x_31757 = x_31753 & x_31756;
assign x_31758 = x_466 & x_467;
assign x_31759 = x_468 & x_469;
assign x_31760 = x_31758 & x_31759;
assign x_31761 = x_470 & x_471;
assign x_31762 = x_472 & x_473;
assign x_31763 = x_31761 & x_31762;
assign x_31764 = x_31760 & x_31763;
assign x_31765 = x_31757 & x_31764;
assign x_31766 = x_474 & x_475;
assign x_31767 = x_476 & x_477;
assign x_31768 = x_31766 & x_31767;
assign x_31769 = x_478 & x_479;
assign x_31770 = x_480 & x_481;
assign x_31771 = x_31769 & x_31770;
assign x_31772 = x_31768 & x_31771;
assign x_31773 = x_482 & x_483;
assign x_31774 = x_484 & x_485;
assign x_31775 = x_31773 & x_31774;
assign x_31776 = x_486 & x_487;
assign x_31777 = x_488 & x_489;
assign x_31778 = x_31776 & x_31777;
assign x_31779 = x_31775 & x_31778;
assign x_31780 = x_31772 & x_31779;
assign x_31781 = x_31765 & x_31780;
assign x_31782 = x_31751 & x_31781;
assign x_31783 = x_31721 & x_31782;
assign x_31784 = x_31661 & x_31783;
assign x_31785 = x_31540 & x_31784;
assign x_31786 = x_491 & x_492;
assign x_31787 = x_490 & x_31786;
assign x_31788 = x_493 & x_494;
assign x_31789 = x_495 & x_496;
assign x_31790 = x_31788 & x_31789;
assign x_31791 = x_31787 & x_31790;
assign x_31792 = x_497 & x_498;
assign x_31793 = x_499 & x_500;
assign x_31794 = x_31792 & x_31793;
assign x_31795 = x_501 & x_502;
assign x_31796 = x_503 & x_504;
assign x_31797 = x_31795 & x_31796;
assign x_31798 = x_31794 & x_31797;
assign x_31799 = x_31791 & x_31798;
assign x_31800 = x_506 & x_507;
assign x_31801 = x_505 & x_31800;
assign x_31802 = x_508 & x_509;
assign x_31803 = x_510 & x_511;
assign x_31804 = x_31802 & x_31803;
assign x_31805 = x_31801 & x_31804;
assign x_31806 = x_512 & x_513;
assign x_31807 = x_514 & x_515;
assign x_31808 = x_31806 & x_31807;
assign x_31809 = x_516 & x_517;
assign x_31810 = x_518 & x_519;
assign x_31811 = x_31809 & x_31810;
assign x_31812 = x_31808 & x_31811;
assign x_31813 = x_31805 & x_31812;
assign x_31814 = x_31799 & x_31813;
assign x_31815 = x_521 & x_522;
assign x_31816 = x_520 & x_31815;
assign x_31817 = x_523 & x_524;
assign x_31818 = x_525 & x_526;
assign x_31819 = x_31817 & x_31818;
assign x_31820 = x_31816 & x_31819;
assign x_31821 = x_527 & x_528;
assign x_31822 = x_529 & x_530;
assign x_31823 = x_31821 & x_31822;
assign x_31824 = x_531 & x_532;
assign x_31825 = x_533 & x_534;
assign x_31826 = x_31824 & x_31825;
assign x_31827 = x_31823 & x_31826;
assign x_31828 = x_31820 & x_31827;
assign x_31829 = x_535 & x_536;
assign x_31830 = x_537 & x_538;
assign x_31831 = x_31829 & x_31830;
assign x_31832 = x_539 & x_540;
assign x_31833 = x_541 & x_542;
assign x_31834 = x_31832 & x_31833;
assign x_31835 = x_31831 & x_31834;
assign x_31836 = x_543 & x_544;
assign x_31837 = x_545 & x_546;
assign x_31838 = x_31836 & x_31837;
assign x_31839 = x_547 & x_548;
assign x_31840 = x_549 & x_550;
assign x_31841 = x_31839 & x_31840;
assign x_31842 = x_31838 & x_31841;
assign x_31843 = x_31835 & x_31842;
assign x_31844 = x_31828 & x_31843;
assign x_31845 = x_31814 & x_31844;
assign x_31846 = x_552 & x_553;
assign x_31847 = x_551 & x_31846;
assign x_31848 = x_554 & x_555;
assign x_31849 = x_556 & x_557;
assign x_31850 = x_31848 & x_31849;
assign x_31851 = x_31847 & x_31850;
assign x_31852 = x_558 & x_559;
assign x_31853 = x_560 & x_561;
assign x_31854 = x_31852 & x_31853;
assign x_31855 = x_562 & x_563;
assign x_31856 = x_564 & x_565;
assign x_31857 = x_31855 & x_31856;
assign x_31858 = x_31854 & x_31857;
assign x_31859 = x_31851 & x_31858;
assign x_31860 = x_567 & x_568;
assign x_31861 = x_566 & x_31860;
assign x_31862 = x_569 & x_570;
assign x_31863 = x_571 & x_572;
assign x_31864 = x_31862 & x_31863;
assign x_31865 = x_31861 & x_31864;
assign x_31866 = x_573 & x_574;
assign x_31867 = x_575 & x_576;
assign x_31868 = x_31866 & x_31867;
assign x_31869 = x_577 & x_578;
assign x_31870 = x_579 & x_580;
assign x_31871 = x_31869 & x_31870;
assign x_31872 = x_31868 & x_31871;
assign x_31873 = x_31865 & x_31872;
assign x_31874 = x_31859 & x_31873;
assign x_31875 = x_582 & x_583;
assign x_31876 = x_581 & x_31875;
assign x_31877 = x_584 & x_585;
assign x_31878 = x_586 & x_587;
assign x_31879 = x_31877 & x_31878;
assign x_31880 = x_31876 & x_31879;
assign x_31881 = x_588 & x_589;
assign x_31882 = x_590 & x_591;
assign x_31883 = x_31881 & x_31882;
assign x_31884 = x_592 & x_593;
assign x_31885 = x_594 & x_595;
assign x_31886 = x_31884 & x_31885;
assign x_31887 = x_31883 & x_31886;
assign x_31888 = x_31880 & x_31887;
assign x_31889 = x_596 & x_597;
assign x_31890 = x_598 & x_599;
assign x_31891 = x_31889 & x_31890;
assign x_31892 = x_600 & x_601;
assign x_31893 = x_602 & x_603;
assign x_31894 = x_31892 & x_31893;
assign x_31895 = x_31891 & x_31894;
assign x_31896 = x_604 & x_605;
assign x_31897 = x_606 & x_607;
assign x_31898 = x_31896 & x_31897;
assign x_31899 = x_608 & x_609;
assign x_31900 = x_610 & x_611;
assign x_31901 = x_31899 & x_31900;
assign x_31902 = x_31898 & x_31901;
assign x_31903 = x_31895 & x_31902;
assign x_31904 = x_31888 & x_31903;
assign x_31905 = x_31874 & x_31904;
assign x_31906 = x_31845 & x_31905;
assign x_31907 = x_613 & x_614;
assign x_31908 = x_612 & x_31907;
assign x_31909 = x_615 & x_616;
assign x_31910 = x_617 & x_618;
assign x_31911 = x_31909 & x_31910;
assign x_31912 = x_31908 & x_31911;
assign x_31913 = x_619 & x_620;
assign x_31914 = x_621 & x_622;
assign x_31915 = x_31913 & x_31914;
assign x_31916 = x_623 & x_624;
assign x_31917 = x_625 & x_626;
assign x_31918 = x_31916 & x_31917;
assign x_31919 = x_31915 & x_31918;
assign x_31920 = x_31912 & x_31919;
assign x_31921 = x_628 & x_629;
assign x_31922 = x_627 & x_31921;
assign x_31923 = x_630 & x_631;
assign x_31924 = x_632 & x_633;
assign x_31925 = x_31923 & x_31924;
assign x_31926 = x_31922 & x_31925;
assign x_31927 = x_634 & x_635;
assign x_31928 = x_636 & x_637;
assign x_31929 = x_31927 & x_31928;
assign x_31930 = x_638 & x_639;
assign x_31931 = x_640 & x_641;
assign x_31932 = x_31930 & x_31931;
assign x_31933 = x_31929 & x_31932;
assign x_31934 = x_31926 & x_31933;
assign x_31935 = x_31920 & x_31934;
assign x_31936 = x_643 & x_644;
assign x_31937 = x_642 & x_31936;
assign x_31938 = x_645 & x_646;
assign x_31939 = x_647 & x_648;
assign x_31940 = x_31938 & x_31939;
assign x_31941 = x_31937 & x_31940;
assign x_31942 = x_649 & x_650;
assign x_31943 = x_651 & x_652;
assign x_31944 = x_31942 & x_31943;
assign x_31945 = x_653 & x_654;
assign x_31946 = x_655 & x_656;
assign x_31947 = x_31945 & x_31946;
assign x_31948 = x_31944 & x_31947;
assign x_31949 = x_31941 & x_31948;
assign x_31950 = x_657 & x_658;
assign x_31951 = x_659 & x_660;
assign x_31952 = x_31950 & x_31951;
assign x_31953 = x_661 & x_662;
assign x_31954 = x_663 & x_664;
assign x_31955 = x_31953 & x_31954;
assign x_31956 = x_31952 & x_31955;
assign x_31957 = x_665 & x_666;
assign x_31958 = x_667 & x_668;
assign x_31959 = x_31957 & x_31958;
assign x_31960 = x_669 & x_670;
assign x_31961 = x_671 & x_672;
assign x_31962 = x_31960 & x_31961;
assign x_31963 = x_31959 & x_31962;
assign x_31964 = x_31956 & x_31963;
assign x_31965 = x_31949 & x_31964;
assign x_31966 = x_31935 & x_31965;
assign x_31967 = x_674 & x_675;
assign x_31968 = x_673 & x_31967;
assign x_31969 = x_676 & x_677;
assign x_31970 = x_678 & x_679;
assign x_31971 = x_31969 & x_31970;
assign x_31972 = x_31968 & x_31971;
assign x_31973 = x_680 & x_681;
assign x_31974 = x_682 & x_683;
assign x_31975 = x_31973 & x_31974;
assign x_31976 = x_684 & x_685;
assign x_31977 = x_686 & x_687;
assign x_31978 = x_31976 & x_31977;
assign x_31979 = x_31975 & x_31978;
assign x_31980 = x_31972 & x_31979;
assign x_31981 = x_689 & x_690;
assign x_31982 = x_688 & x_31981;
assign x_31983 = x_691 & x_692;
assign x_31984 = x_693 & x_694;
assign x_31985 = x_31983 & x_31984;
assign x_31986 = x_31982 & x_31985;
assign x_31987 = x_695 & x_696;
assign x_31988 = x_697 & x_698;
assign x_31989 = x_31987 & x_31988;
assign x_31990 = x_699 & x_700;
assign x_31991 = x_701 & x_702;
assign x_31992 = x_31990 & x_31991;
assign x_31993 = x_31989 & x_31992;
assign x_31994 = x_31986 & x_31993;
assign x_31995 = x_31980 & x_31994;
assign x_31996 = x_704 & x_705;
assign x_31997 = x_703 & x_31996;
assign x_31998 = x_706 & x_707;
assign x_31999 = x_708 & x_709;
assign x_32000 = x_31998 & x_31999;
assign x_32001 = x_31997 & x_32000;
assign x_32002 = x_710 & x_711;
assign x_32003 = x_712 & x_713;
assign x_32004 = x_32002 & x_32003;
assign x_32005 = x_714 & x_715;
assign x_32006 = x_716 & x_717;
assign x_32007 = x_32005 & x_32006;
assign x_32008 = x_32004 & x_32007;
assign x_32009 = x_32001 & x_32008;
assign x_32010 = x_718 & x_719;
assign x_32011 = x_720 & x_721;
assign x_32012 = x_32010 & x_32011;
assign x_32013 = x_722 & x_723;
assign x_32014 = x_724 & x_725;
assign x_32015 = x_32013 & x_32014;
assign x_32016 = x_32012 & x_32015;
assign x_32017 = x_726 & x_727;
assign x_32018 = x_728 & x_729;
assign x_32019 = x_32017 & x_32018;
assign x_32020 = x_730 & x_731;
assign x_32021 = x_732 & x_733;
assign x_32022 = x_32020 & x_32021;
assign x_32023 = x_32019 & x_32022;
assign x_32024 = x_32016 & x_32023;
assign x_32025 = x_32009 & x_32024;
assign x_32026 = x_31995 & x_32025;
assign x_32027 = x_31966 & x_32026;
assign x_32028 = x_31906 & x_32027;
assign x_32029 = x_735 & x_736;
assign x_32030 = x_734 & x_32029;
assign x_32031 = x_737 & x_738;
assign x_32032 = x_739 & x_740;
assign x_32033 = x_32031 & x_32032;
assign x_32034 = x_32030 & x_32033;
assign x_32035 = x_741 & x_742;
assign x_32036 = x_743 & x_744;
assign x_32037 = x_32035 & x_32036;
assign x_32038 = x_745 & x_746;
assign x_32039 = x_747 & x_748;
assign x_32040 = x_32038 & x_32039;
assign x_32041 = x_32037 & x_32040;
assign x_32042 = x_32034 & x_32041;
assign x_32043 = x_750 & x_751;
assign x_32044 = x_749 & x_32043;
assign x_32045 = x_752 & x_753;
assign x_32046 = x_754 & x_755;
assign x_32047 = x_32045 & x_32046;
assign x_32048 = x_32044 & x_32047;
assign x_32049 = x_756 & x_757;
assign x_32050 = x_758 & x_759;
assign x_32051 = x_32049 & x_32050;
assign x_32052 = x_760 & x_761;
assign x_32053 = x_762 & x_763;
assign x_32054 = x_32052 & x_32053;
assign x_32055 = x_32051 & x_32054;
assign x_32056 = x_32048 & x_32055;
assign x_32057 = x_32042 & x_32056;
assign x_32058 = x_765 & x_766;
assign x_32059 = x_764 & x_32058;
assign x_32060 = x_767 & x_768;
assign x_32061 = x_769 & x_770;
assign x_32062 = x_32060 & x_32061;
assign x_32063 = x_32059 & x_32062;
assign x_32064 = x_771 & x_772;
assign x_32065 = x_773 & x_774;
assign x_32066 = x_32064 & x_32065;
assign x_32067 = x_775 & x_776;
assign x_32068 = x_777 & x_778;
assign x_32069 = x_32067 & x_32068;
assign x_32070 = x_32066 & x_32069;
assign x_32071 = x_32063 & x_32070;
assign x_32072 = x_779 & x_780;
assign x_32073 = x_781 & x_782;
assign x_32074 = x_32072 & x_32073;
assign x_32075 = x_783 & x_784;
assign x_32076 = x_785 & x_786;
assign x_32077 = x_32075 & x_32076;
assign x_32078 = x_32074 & x_32077;
assign x_32079 = x_787 & x_788;
assign x_32080 = x_789 & x_790;
assign x_32081 = x_32079 & x_32080;
assign x_32082 = x_791 & x_792;
assign x_32083 = x_793 & x_794;
assign x_32084 = x_32082 & x_32083;
assign x_32085 = x_32081 & x_32084;
assign x_32086 = x_32078 & x_32085;
assign x_32087 = x_32071 & x_32086;
assign x_32088 = x_32057 & x_32087;
assign x_32089 = x_796 & x_797;
assign x_32090 = x_795 & x_32089;
assign x_32091 = x_798 & x_799;
assign x_32092 = x_800 & x_801;
assign x_32093 = x_32091 & x_32092;
assign x_32094 = x_32090 & x_32093;
assign x_32095 = x_802 & x_803;
assign x_32096 = x_804 & x_805;
assign x_32097 = x_32095 & x_32096;
assign x_32098 = x_806 & x_807;
assign x_32099 = x_808 & x_809;
assign x_32100 = x_32098 & x_32099;
assign x_32101 = x_32097 & x_32100;
assign x_32102 = x_32094 & x_32101;
assign x_32103 = x_811 & x_812;
assign x_32104 = x_810 & x_32103;
assign x_32105 = x_813 & x_814;
assign x_32106 = x_815 & x_816;
assign x_32107 = x_32105 & x_32106;
assign x_32108 = x_32104 & x_32107;
assign x_32109 = x_817 & x_818;
assign x_32110 = x_819 & x_820;
assign x_32111 = x_32109 & x_32110;
assign x_32112 = x_821 & x_822;
assign x_32113 = x_823 & x_824;
assign x_32114 = x_32112 & x_32113;
assign x_32115 = x_32111 & x_32114;
assign x_32116 = x_32108 & x_32115;
assign x_32117 = x_32102 & x_32116;
assign x_32118 = x_826 & x_827;
assign x_32119 = x_825 & x_32118;
assign x_32120 = x_828 & x_829;
assign x_32121 = x_830 & x_831;
assign x_32122 = x_32120 & x_32121;
assign x_32123 = x_32119 & x_32122;
assign x_32124 = x_832 & x_833;
assign x_32125 = x_834 & x_835;
assign x_32126 = x_32124 & x_32125;
assign x_32127 = x_836 & x_837;
assign x_32128 = x_838 & x_839;
assign x_32129 = x_32127 & x_32128;
assign x_32130 = x_32126 & x_32129;
assign x_32131 = x_32123 & x_32130;
assign x_32132 = x_840 & x_841;
assign x_32133 = x_842 & x_843;
assign x_32134 = x_32132 & x_32133;
assign x_32135 = x_844 & x_845;
assign x_32136 = x_846 & x_847;
assign x_32137 = x_32135 & x_32136;
assign x_32138 = x_32134 & x_32137;
assign x_32139 = x_848 & x_849;
assign x_32140 = x_850 & x_851;
assign x_32141 = x_32139 & x_32140;
assign x_32142 = x_852 & x_853;
assign x_32143 = x_854 & x_855;
assign x_32144 = x_32142 & x_32143;
assign x_32145 = x_32141 & x_32144;
assign x_32146 = x_32138 & x_32145;
assign x_32147 = x_32131 & x_32146;
assign x_32148 = x_32117 & x_32147;
assign x_32149 = x_32088 & x_32148;
assign x_32150 = x_857 & x_858;
assign x_32151 = x_856 & x_32150;
assign x_32152 = x_859 & x_860;
assign x_32153 = x_861 & x_862;
assign x_32154 = x_32152 & x_32153;
assign x_32155 = x_32151 & x_32154;
assign x_32156 = x_863 & x_864;
assign x_32157 = x_865 & x_866;
assign x_32158 = x_32156 & x_32157;
assign x_32159 = x_867 & x_868;
assign x_32160 = x_869 & x_870;
assign x_32161 = x_32159 & x_32160;
assign x_32162 = x_32158 & x_32161;
assign x_32163 = x_32155 & x_32162;
assign x_32164 = x_872 & x_873;
assign x_32165 = x_871 & x_32164;
assign x_32166 = x_874 & x_875;
assign x_32167 = x_876 & x_877;
assign x_32168 = x_32166 & x_32167;
assign x_32169 = x_32165 & x_32168;
assign x_32170 = x_878 & x_879;
assign x_32171 = x_880 & x_881;
assign x_32172 = x_32170 & x_32171;
assign x_32173 = x_882 & x_883;
assign x_32174 = x_884 & x_885;
assign x_32175 = x_32173 & x_32174;
assign x_32176 = x_32172 & x_32175;
assign x_32177 = x_32169 & x_32176;
assign x_32178 = x_32163 & x_32177;
assign x_32179 = x_887 & x_888;
assign x_32180 = x_886 & x_32179;
assign x_32181 = x_889 & x_890;
assign x_32182 = x_891 & x_892;
assign x_32183 = x_32181 & x_32182;
assign x_32184 = x_32180 & x_32183;
assign x_32185 = x_893 & x_894;
assign x_32186 = x_895 & x_896;
assign x_32187 = x_32185 & x_32186;
assign x_32188 = x_897 & x_898;
assign x_32189 = x_899 & x_900;
assign x_32190 = x_32188 & x_32189;
assign x_32191 = x_32187 & x_32190;
assign x_32192 = x_32184 & x_32191;
assign x_32193 = x_901 & x_902;
assign x_32194 = x_903 & x_904;
assign x_32195 = x_32193 & x_32194;
assign x_32196 = x_905 & x_906;
assign x_32197 = x_907 & x_908;
assign x_32198 = x_32196 & x_32197;
assign x_32199 = x_32195 & x_32198;
assign x_32200 = x_909 & x_910;
assign x_32201 = x_911 & x_912;
assign x_32202 = x_32200 & x_32201;
assign x_32203 = x_913 & x_914;
assign x_32204 = x_915 & x_916;
assign x_32205 = x_32203 & x_32204;
assign x_32206 = x_32202 & x_32205;
assign x_32207 = x_32199 & x_32206;
assign x_32208 = x_32192 & x_32207;
assign x_32209 = x_32178 & x_32208;
assign x_32210 = x_918 & x_919;
assign x_32211 = x_917 & x_32210;
assign x_32212 = x_920 & x_921;
assign x_32213 = x_922 & x_923;
assign x_32214 = x_32212 & x_32213;
assign x_32215 = x_32211 & x_32214;
assign x_32216 = x_924 & x_925;
assign x_32217 = x_926 & x_927;
assign x_32218 = x_32216 & x_32217;
assign x_32219 = x_928 & x_929;
assign x_32220 = x_930 & x_931;
assign x_32221 = x_32219 & x_32220;
assign x_32222 = x_32218 & x_32221;
assign x_32223 = x_32215 & x_32222;
assign x_32224 = x_932 & x_933;
assign x_32225 = x_934 & x_935;
assign x_32226 = x_32224 & x_32225;
assign x_32227 = x_936 & x_937;
assign x_32228 = x_938 & x_939;
assign x_32229 = x_32227 & x_32228;
assign x_32230 = x_32226 & x_32229;
assign x_32231 = x_940 & x_941;
assign x_32232 = x_942 & x_943;
assign x_32233 = x_32231 & x_32232;
assign x_32234 = x_944 & x_945;
assign x_32235 = x_946 & x_947;
assign x_32236 = x_32234 & x_32235;
assign x_32237 = x_32233 & x_32236;
assign x_32238 = x_32230 & x_32237;
assign x_32239 = x_32223 & x_32238;
assign x_32240 = x_949 & x_950;
assign x_32241 = x_948 & x_32240;
assign x_32242 = x_951 & x_952;
assign x_32243 = x_953 & x_954;
assign x_32244 = x_32242 & x_32243;
assign x_32245 = x_32241 & x_32244;
assign x_32246 = x_955 & x_956;
assign x_32247 = x_957 & x_958;
assign x_32248 = x_32246 & x_32247;
assign x_32249 = x_959 & x_960;
assign x_32250 = x_961 & x_962;
assign x_32251 = x_32249 & x_32250;
assign x_32252 = x_32248 & x_32251;
assign x_32253 = x_32245 & x_32252;
assign x_32254 = x_963 & x_964;
assign x_32255 = x_965 & x_966;
assign x_32256 = x_32254 & x_32255;
assign x_32257 = x_967 & x_968;
assign x_32258 = x_969 & x_970;
assign x_32259 = x_32257 & x_32258;
assign x_32260 = x_32256 & x_32259;
assign x_32261 = x_971 & x_972;
assign x_32262 = x_973 & x_974;
assign x_32263 = x_32261 & x_32262;
assign x_32264 = x_975 & x_976;
assign x_32265 = x_977 & x_978;
assign x_32266 = x_32264 & x_32265;
assign x_32267 = x_32263 & x_32266;
assign x_32268 = x_32260 & x_32267;
assign x_32269 = x_32253 & x_32268;
assign x_32270 = x_32239 & x_32269;
assign x_32271 = x_32209 & x_32270;
assign x_32272 = x_32149 & x_32271;
assign x_32273 = x_32028 & x_32272;
assign x_32274 = x_31785 & x_32273;
assign x_32275 = x_980 & x_981;
assign x_32276 = x_979 & x_32275;
assign x_32277 = x_982 & x_983;
assign x_32278 = x_984 & x_985;
assign x_32279 = x_32277 & x_32278;
assign x_32280 = x_32276 & x_32279;
assign x_32281 = x_986 & x_987;
assign x_32282 = x_988 & x_989;
assign x_32283 = x_32281 & x_32282;
assign x_32284 = x_990 & x_991;
assign x_32285 = x_992 & x_993;
assign x_32286 = x_32284 & x_32285;
assign x_32287 = x_32283 & x_32286;
assign x_32288 = x_32280 & x_32287;
assign x_32289 = x_995 & x_996;
assign x_32290 = x_994 & x_32289;
assign x_32291 = x_997 & x_998;
assign x_32292 = x_999 & x_1000;
assign x_32293 = x_32291 & x_32292;
assign x_32294 = x_32290 & x_32293;
assign x_32295 = x_1001 & x_1002;
assign x_32296 = x_1003 & x_1004;
assign x_32297 = x_32295 & x_32296;
assign x_32298 = x_1005 & x_1006;
assign x_32299 = x_1007 & x_1008;
assign x_32300 = x_32298 & x_32299;
assign x_32301 = x_32297 & x_32300;
assign x_32302 = x_32294 & x_32301;
assign x_32303 = x_32288 & x_32302;
assign x_32304 = x_1010 & x_1011;
assign x_32305 = x_1009 & x_32304;
assign x_32306 = x_1012 & x_1013;
assign x_32307 = x_1014 & x_1015;
assign x_32308 = x_32306 & x_32307;
assign x_32309 = x_32305 & x_32308;
assign x_32310 = x_1016 & x_1017;
assign x_32311 = x_1018 & x_1019;
assign x_32312 = x_32310 & x_32311;
assign x_32313 = x_1020 & x_1021;
assign x_32314 = x_1022 & x_1023;
assign x_32315 = x_32313 & x_32314;
assign x_32316 = x_32312 & x_32315;
assign x_32317 = x_32309 & x_32316;
assign x_32318 = x_1024 & x_1025;
assign x_32319 = x_1026 & x_1027;
assign x_32320 = x_32318 & x_32319;
assign x_32321 = x_1028 & x_1029;
assign x_32322 = x_1030 & x_1031;
assign x_32323 = x_32321 & x_32322;
assign x_32324 = x_32320 & x_32323;
assign x_32325 = x_1032 & x_1033;
assign x_32326 = x_1034 & x_1035;
assign x_32327 = x_32325 & x_32326;
assign x_32328 = x_1036 & x_1037;
assign x_32329 = x_1038 & x_1039;
assign x_32330 = x_32328 & x_32329;
assign x_32331 = x_32327 & x_32330;
assign x_32332 = x_32324 & x_32331;
assign x_32333 = x_32317 & x_32332;
assign x_32334 = x_32303 & x_32333;
assign x_32335 = x_1041 & x_1042;
assign x_32336 = x_1040 & x_32335;
assign x_32337 = x_1043 & x_1044;
assign x_32338 = x_1045 & x_1046;
assign x_32339 = x_32337 & x_32338;
assign x_32340 = x_32336 & x_32339;
assign x_32341 = x_1047 & x_1048;
assign x_32342 = x_1049 & x_1050;
assign x_32343 = x_32341 & x_32342;
assign x_32344 = x_1051 & x_1052;
assign x_32345 = x_1053 & x_1054;
assign x_32346 = x_32344 & x_32345;
assign x_32347 = x_32343 & x_32346;
assign x_32348 = x_32340 & x_32347;
assign x_32349 = x_1056 & x_1057;
assign x_32350 = x_1055 & x_32349;
assign x_32351 = x_1058 & x_1059;
assign x_32352 = x_1060 & x_1061;
assign x_32353 = x_32351 & x_32352;
assign x_32354 = x_32350 & x_32353;
assign x_32355 = x_1062 & x_1063;
assign x_32356 = x_1064 & x_1065;
assign x_32357 = x_32355 & x_32356;
assign x_32358 = x_1066 & x_1067;
assign x_32359 = x_1068 & x_1069;
assign x_32360 = x_32358 & x_32359;
assign x_32361 = x_32357 & x_32360;
assign x_32362 = x_32354 & x_32361;
assign x_32363 = x_32348 & x_32362;
assign x_32364 = x_1071 & x_1072;
assign x_32365 = x_1070 & x_32364;
assign x_32366 = x_1073 & x_1074;
assign x_32367 = x_1075 & x_1076;
assign x_32368 = x_32366 & x_32367;
assign x_32369 = x_32365 & x_32368;
assign x_32370 = x_1077 & x_1078;
assign x_32371 = x_1079 & x_1080;
assign x_32372 = x_32370 & x_32371;
assign x_32373 = x_1081 & x_1082;
assign x_32374 = x_1083 & x_1084;
assign x_32375 = x_32373 & x_32374;
assign x_32376 = x_32372 & x_32375;
assign x_32377 = x_32369 & x_32376;
assign x_32378 = x_1085 & x_1086;
assign x_32379 = x_1087 & x_1088;
assign x_32380 = x_32378 & x_32379;
assign x_32381 = x_1089 & x_1090;
assign x_32382 = x_1091 & x_1092;
assign x_32383 = x_32381 & x_32382;
assign x_32384 = x_32380 & x_32383;
assign x_32385 = x_1093 & x_1094;
assign x_32386 = x_1095 & x_1096;
assign x_32387 = x_32385 & x_32386;
assign x_32388 = x_1097 & x_1098;
assign x_32389 = x_1099 & x_1100;
assign x_32390 = x_32388 & x_32389;
assign x_32391 = x_32387 & x_32390;
assign x_32392 = x_32384 & x_32391;
assign x_32393 = x_32377 & x_32392;
assign x_32394 = x_32363 & x_32393;
assign x_32395 = x_32334 & x_32394;
assign x_32396 = x_1102 & x_1103;
assign x_32397 = x_1101 & x_32396;
assign x_32398 = x_1104 & x_1105;
assign x_32399 = x_1106 & x_1107;
assign x_32400 = x_32398 & x_32399;
assign x_32401 = x_32397 & x_32400;
assign x_32402 = x_1108 & x_1109;
assign x_32403 = x_1110 & x_1111;
assign x_32404 = x_32402 & x_32403;
assign x_32405 = x_1112 & x_1113;
assign x_32406 = x_1114 & x_1115;
assign x_32407 = x_32405 & x_32406;
assign x_32408 = x_32404 & x_32407;
assign x_32409 = x_32401 & x_32408;
assign x_32410 = x_1117 & x_1118;
assign x_32411 = x_1116 & x_32410;
assign x_32412 = x_1119 & x_1120;
assign x_32413 = x_1121 & x_1122;
assign x_32414 = x_32412 & x_32413;
assign x_32415 = x_32411 & x_32414;
assign x_32416 = x_1123 & x_1124;
assign x_32417 = x_1125 & x_1126;
assign x_32418 = x_32416 & x_32417;
assign x_32419 = x_1127 & x_1128;
assign x_32420 = x_1129 & x_1130;
assign x_32421 = x_32419 & x_32420;
assign x_32422 = x_32418 & x_32421;
assign x_32423 = x_32415 & x_32422;
assign x_32424 = x_32409 & x_32423;
assign x_32425 = x_1132 & x_1133;
assign x_32426 = x_1131 & x_32425;
assign x_32427 = x_1134 & x_1135;
assign x_32428 = x_1136 & x_1137;
assign x_32429 = x_32427 & x_32428;
assign x_32430 = x_32426 & x_32429;
assign x_32431 = x_1138 & x_1139;
assign x_32432 = x_1140 & x_1141;
assign x_32433 = x_32431 & x_32432;
assign x_32434 = x_1142 & x_1143;
assign x_32435 = x_1144 & x_1145;
assign x_32436 = x_32434 & x_32435;
assign x_32437 = x_32433 & x_32436;
assign x_32438 = x_32430 & x_32437;
assign x_32439 = x_1146 & x_1147;
assign x_32440 = x_1148 & x_1149;
assign x_32441 = x_32439 & x_32440;
assign x_32442 = x_1150 & x_1151;
assign x_32443 = x_1152 & x_1153;
assign x_32444 = x_32442 & x_32443;
assign x_32445 = x_32441 & x_32444;
assign x_32446 = x_1154 & x_1155;
assign x_32447 = x_1156 & x_1157;
assign x_32448 = x_32446 & x_32447;
assign x_32449 = x_1158 & x_1159;
assign x_32450 = x_1160 & x_1161;
assign x_32451 = x_32449 & x_32450;
assign x_32452 = x_32448 & x_32451;
assign x_32453 = x_32445 & x_32452;
assign x_32454 = x_32438 & x_32453;
assign x_32455 = x_32424 & x_32454;
assign x_32456 = x_1163 & x_1164;
assign x_32457 = x_1162 & x_32456;
assign x_32458 = x_1165 & x_1166;
assign x_32459 = x_1167 & x_1168;
assign x_32460 = x_32458 & x_32459;
assign x_32461 = x_32457 & x_32460;
assign x_32462 = x_1169 & x_1170;
assign x_32463 = x_1171 & x_1172;
assign x_32464 = x_32462 & x_32463;
assign x_32465 = x_1173 & x_1174;
assign x_32466 = x_1175 & x_1176;
assign x_32467 = x_32465 & x_32466;
assign x_32468 = x_32464 & x_32467;
assign x_32469 = x_32461 & x_32468;
assign x_32470 = x_1178 & x_1179;
assign x_32471 = x_1177 & x_32470;
assign x_32472 = x_1180 & x_1181;
assign x_32473 = x_1182 & x_1183;
assign x_32474 = x_32472 & x_32473;
assign x_32475 = x_32471 & x_32474;
assign x_32476 = x_1184 & x_1185;
assign x_32477 = x_1186 & x_1187;
assign x_32478 = x_32476 & x_32477;
assign x_32479 = x_1188 & x_1189;
assign x_32480 = x_1190 & x_1191;
assign x_32481 = x_32479 & x_32480;
assign x_32482 = x_32478 & x_32481;
assign x_32483 = x_32475 & x_32482;
assign x_32484 = x_32469 & x_32483;
assign x_32485 = x_1193 & x_1194;
assign x_32486 = x_1192 & x_32485;
assign x_32487 = x_1195 & x_1196;
assign x_32488 = x_1197 & x_1198;
assign x_32489 = x_32487 & x_32488;
assign x_32490 = x_32486 & x_32489;
assign x_32491 = x_1199 & x_1200;
assign x_32492 = x_1201 & x_1202;
assign x_32493 = x_32491 & x_32492;
assign x_32494 = x_1203 & x_1204;
assign x_32495 = x_1205 & x_1206;
assign x_32496 = x_32494 & x_32495;
assign x_32497 = x_32493 & x_32496;
assign x_32498 = x_32490 & x_32497;
assign x_32499 = x_1207 & x_1208;
assign x_32500 = x_1209 & x_1210;
assign x_32501 = x_32499 & x_32500;
assign x_32502 = x_1211 & x_1212;
assign x_32503 = x_1213 & x_1214;
assign x_32504 = x_32502 & x_32503;
assign x_32505 = x_32501 & x_32504;
assign x_32506 = x_1215 & x_1216;
assign x_32507 = x_1217 & x_1218;
assign x_32508 = x_32506 & x_32507;
assign x_32509 = x_1219 & x_1220;
assign x_32510 = x_1221 & x_1222;
assign x_32511 = x_32509 & x_32510;
assign x_32512 = x_32508 & x_32511;
assign x_32513 = x_32505 & x_32512;
assign x_32514 = x_32498 & x_32513;
assign x_32515 = x_32484 & x_32514;
assign x_32516 = x_32455 & x_32515;
assign x_32517 = x_32395 & x_32516;
assign x_32518 = x_1224 & x_1225;
assign x_32519 = x_1223 & x_32518;
assign x_32520 = x_1226 & x_1227;
assign x_32521 = x_1228 & x_1229;
assign x_32522 = x_32520 & x_32521;
assign x_32523 = x_32519 & x_32522;
assign x_32524 = x_1230 & x_1231;
assign x_32525 = x_1232 & x_1233;
assign x_32526 = x_32524 & x_32525;
assign x_32527 = x_1234 & x_1235;
assign x_32528 = x_1236 & x_1237;
assign x_32529 = x_32527 & x_32528;
assign x_32530 = x_32526 & x_32529;
assign x_32531 = x_32523 & x_32530;
assign x_32532 = x_1239 & x_1240;
assign x_32533 = x_1238 & x_32532;
assign x_32534 = x_1241 & x_1242;
assign x_32535 = x_1243 & x_1244;
assign x_32536 = x_32534 & x_32535;
assign x_32537 = x_32533 & x_32536;
assign x_32538 = x_1245 & x_1246;
assign x_32539 = x_1247 & x_1248;
assign x_32540 = x_32538 & x_32539;
assign x_32541 = x_1249 & x_1250;
assign x_32542 = x_1251 & x_1252;
assign x_32543 = x_32541 & x_32542;
assign x_32544 = x_32540 & x_32543;
assign x_32545 = x_32537 & x_32544;
assign x_32546 = x_32531 & x_32545;
assign x_32547 = x_1254 & x_1255;
assign x_32548 = x_1253 & x_32547;
assign x_32549 = x_1256 & x_1257;
assign x_32550 = x_1258 & x_1259;
assign x_32551 = x_32549 & x_32550;
assign x_32552 = x_32548 & x_32551;
assign x_32553 = x_1260 & x_1261;
assign x_32554 = x_1262 & x_1263;
assign x_32555 = x_32553 & x_32554;
assign x_32556 = x_1264 & x_1265;
assign x_32557 = x_1266 & x_1267;
assign x_32558 = x_32556 & x_32557;
assign x_32559 = x_32555 & x_32558;
assign x_32560 = x_32552 & x_32559;
assign x_32561 = x_1268 & x_1269;
assign x_32562 = x_1270 & x_1271;
assign x_32563 = x_32561 & x_32562;
assign x_32564 = x_1272 & x_1273;
assign x_32565 = x_1274 & x_1275;
assign x_32566 = x_32564 & x_32565;
assign x_32567 = x_32563 & x_32566;
assign x_32568 = x_1276 & x_1277;
assign x_32569 = x_1278 & x_1279;
assign x_32570 = x_32568 & x_32569;
assign x_32571 = x_1280 & x_1281;
assign x_32572 = x_1282 & x_1283;
assign x_32573 = x_32571 & x_32572;
assign x_32574 = x_32570 & x_32573;
assign x_32575 = x_32567 & x_32574;
assign x_32576 = x_32560 & x_32575;
assign x_32577 = x_32546 & x_32576;
assign x_32578 = x_1285 & x_1286;
assign x_32579 = x_1284 & x_32578;
assign x_32580 = x_1287 & x_1288;
assign x_32581 = x_1289 & x_1290;
assign x_32582 = x_32580 & x_32581;
assign x_32583 = x_32579 & x_32582;
assign x_32584 = x_1291 & x_1292;
assign x_32585 = x_1293 & x_1294;
assign x_32586 = x_32584 & x_32585;
assign x_32587 = x_1295 & x_1296;
assign x_32588 = x_1297 & x_1298;
assign x_32589 = x_32587 & x_32588;
assign x_32590 = x_32586 & x_32589;
assign x_32591 = x_32583 & x_32590;
assign x_32592 = x_1300 & x_1301;
assign x_32593 = x_1299 & x_32592;
assign x_32594 = x_1302 & x_1303;
assign x_32595 = x_1304 & x_1305;
assign x_32596 = x_32594 & x_32595;
assign x_32597 = x_32593 & x_32596;
assign x_32598 = x_1306 & x_1307;
assign x_32599 = x_1308 & x_1309;
assign x_32600 = x_32598 & x_32599;
assign x_32601 = x_1310 & x_1311;
assign x_32602 = x_1312 & x_1313;
assign x_32603 = x_32601 & x_32602;
assign x_32604 = x_32600 & x_32603;
assign x_32605 = x_32597 & x_32604;
assign x_32606 = x_32591 & x_32605;
assign x_32607 = x_1315 & x_1316;
assign x_32608 = x_1314 & x_32607;
assign x_32609 = x_1317 & x_1318;
assign x_32610 = x_1319 & x_1320;
assign x_32611 = x_32609 & x_32610;
assign x_32612 = x_32608 & x_32611;
assign x_32613 = x_1321 & x_1322;
assign x_32614 = x_1323 & x_1324;
assign x_32615 = x_32613 & x_32614;
assign x_32616 = x_1325 & x_1326;
assign x_32617 = x_1327 & x_1328;
assign x_32618 = x_32616 & x_32617;
assign x_32619 = x_32615 & x_32618;
assign x_32620 = x_32612 & x_32619;
assign x_32621 = x_1329 & x_1330;
assign x_32622 = x_1331 & x_1332;
assign x_32623 = x_32621 & x_32622;
assign x_32624 = x_1333 & x_1334;
assign x_32625 = x_1335 & x_1336;
assign x_32626 = x_32624 & x_32625;
assign x_32627 = x_32623 & x_32626;
assign x_32628 = x_1337 & x_1338;
assign x_32629 = x_1339 & x_1340;
assign x_32630 = x_32628 & x_32629;
assign x_32631 = x_1341 & x_1342;
assign x_32632 = x_1343 & x_1344;
assign x_32633 = x_32631 & x_32632;
assign x_32634 = x_32630 & x_32633;
assign x_32635 = x_32627 & x_32634;
assign x_32636 = x_32620 & x_32635;
assign x_32637 = x_32606 & x_32636;
assign x_32638 = x_32577 & x_32637;
assign x_32639 = x_1346 & x_1347;
assign x_32640 = x_1345 & x_32639;
assign x_32641 = x_1348 & x_1349;
assign x_32642 = x_1350 & x_1351;
assign x_32643 = x_32641 & x_32642;
assign x_32644 = x_32640 & x_32643;
assign x_32645 = x_1352 & x_1353;
assign x_32646 = x_1354 & x_1355;
assign x_32647 = x_32645 & x_32646;
assign x_32648 = x_1356 & x_1357;
assign x_32649 = x_1358 & x_1359;
assign x_32650 = x_32648 & x_32649;
assign x_32651 = x_32647 & x_32650;
assign x_32652 = x_32644 & x_32651;
assign x_32653 = x_1361 & x_1362;
assign x_32654 = x_1360 & x_32653;
assign x_32655 = x_1363 & x_1364;
assign x_32656 = x_1365 & x_1366;
assign x_32657 = x_32655 & x_32656;
assign x_32658 = x_32654 & x_32657;
assign x_32659 = x_1367 & x_1368;
assign x_32660 = x_1369 & x_1370;
assign x_32661 = x_32659 & x_32660;
assign x_32662 = x_1371 & x_1372;
assign x_32663 = x_1373 & x_1374;
assign x_32664 = x_32662 & x_32663;
assign x_32665 = x_32661 & x_32664;
assign x_32666 = x_32658 & x_32665;
assign x_32667 = x_32652 & x_32666;
assign x_32668 = x_1376 & x_1377;
assign x_32669 = x_1375 & x_32668;
assign x_32670 = x_1378 & x_1379;
assign x_32671 = x_1380 & x_1381;
assign x_32672 = x_32670 & x_32671;
assign x_32673 = x_32669 & x_32672;
assign x_32674 = x_1382 & x_1383;
assign x_32675 = x_1384 & x_1385;
assign x_32676 = x_32674 & x_32675;
assign x_32677 = x_1386 & x_1387;
assign x_32678 = x_1388 & x_1389;
assign x_32679 = x_32677 & x_32678;
assign x_32680 = x_32676 & x_32679;
assign x_32681 = x_32673 & x_32680;
assign x_32682 = x_1390 & x_1391;
assign x_32683 = x_1392 & x_1393;
assign x_32684 = x_32682 & x_32683;
assign x_32685 = x_1394 & x_1395;
assign x_32686 = x_1396 & x_1397;
assign x_32687 = x_32685 & x_32686;
assign x_32688 = x_32684 & x_32687;
assign x_32689 = x_1398 & x_1399;
assign x_32690 = x_1400 & x_1401;
assign x_32691 = x_32689 & x_32690;
assign x_32692 = x_1402 & x_1403;
assign x_32693 = x_1404 & x_1405;
assign x_32694 = x_32692 & x_32693;
assign x_32695 = x_32691 & x_32694;
assign x_32696 = x_32688 & x_32695;
assign x_32697 = x_32681 & x_32696;
assign x_32698 = x_32667 & x_32697;
assign x_32699 = x_1407 & x_1408;
assign x_32700 = x_1406 & x_32699;
assign x_32701 = x_1409 & x_1410;
assign x_32702 = x_1411 & x_1412;
assign x_32703 = x_32701 & x_32702;
assign x_32704 = x_32700 & x_32703;
assign x_32705 = x_1413 & x_1414;
assign x_32706 = x_1415 & x_1416;
assign x_32707 = x_32705 & x_32706;
assign x_32708 = x_1417 & x_1418;
assign x_32709 = x_1419 & x_1420;
assign x_32710 = x_32708 & x_32709;
assign x_32711 = x_32707 & x_32710;
assign x_32712 = x_32704 & x_32711;
assign x_32713 = x_1421 & x_1422;
assign x_32714 = x_1423 & x_1424;
assign x_32715 = x_32713 & x_32714;
assign x_32716 = x_1425 & x_1426;
assign x_32717 = x_1427 & x_1428;
assign x_32718 = x_32716 & x_32717;
assign x_32719 = x_32715 & x_32718;
assign x_32720 = x_1429 & x_1430;
assign x_32721 = x_1431 & x_1432;
assign x_32722 = x_32720 & x_32721;
assign x_32723 = x_1433 & x_1434;
assign x_32724 = x_1435 & x_1436;
assign x_32725 = x_32723 & x_32724;
assign x_32726 = x_32722 & x_32725;
assign x_32727 = x_32719 & x_32726;
assign x_32728 = x_32712 & x_32727;
assign x_32729 = x_1438 & x_1439;
assign x_32730 = x_1437 & x_32729;
assign x_32731 = x_1440 & x_1441;
assign x_32732 = x_1442 & x_1443;
assign x_32733 = x_32731 & x_32732;
assign x_32734 = x_32730 & x_32733;
assign x_32735 = x_1444 & x_1445;
assign x_32736 = x_1446 & x_1447;
assign x_32737 = x_32735 & x_32736;
assign x_32738 = x_1448 & x_1449;
assign x_32739 = x_1450 & x_1451;
assign x_32740 = x_32738 & x_32739;
assign x_32741 = x_32737 & x_32740;
assign x_32742 = x_32734 & x_32741;
assign x_32743 = x_1452 & x_1453;
assign x_32744 = x_1454 & x_1455;
assign x_32745 = x_32743 & x_32744;
assign x_32746 = x_1456 & x_1457;
assign x_32747 = x_1458 & x_1459;
assign x_32748 = x_32746 & x_32747;
assign x_32749 = x_32745 & x_32748;
assign x_32750 = x_1460 & x_1461;
assign x_32751 = x_1462 & x_1463;
assign x_32752 = x_32750 & x_32751;
assign x_32753 = x_1464 & x_1465;
assign x_32754 = x_1466 & x_1467;
assign x_32755 = x_32753 & x_32754;
assign x_32756 = x_32752 & x_32755;
assign x_32757 = x_32749 & x_32756;
assign x_32758 = x_32742 & x_32757;
assign x_32759 = x_32728 & x_32758;
assign x_32760 = x_32698 & x_32759;
assign x_32761 = x_32638 & x_32760;
assign x_32762 = x_32517 & x_32761;
assign x_32763 = x_1469 & x_1470;
assign x_32764 = x_1468 & x_32763;
assign x_32765 = x_1471 & x_1472;
assign x_32766 = x_1473 & x_1474;
assign x_32767 = x_32765 & x_32766;
assign x_32768 = x_32764 & x_32767;
assign x_32769 = x_1475 & x_1476;
assign x_32770 = x_1477 & x_1478;
assign x_32771 = x_32769 & x_32770;
assign x_32772 = x_1479 & x_1480;
assign x_32773 = x_1481 & x_1482;
assign x_32774 = x_32772 & x_32773;
assign x_32775 = x_32771 & x_32774;
assign x_32776 = x_32768 & x_32775;
assign x_32777 = x_1484 & x_1485;
assign x_32778 = x_1483 & x_32777;
assign x_32779 = x_1486 & x_1487;
assign x_32780 = x_1488 & x_1489;
assign x_32781 = x_32779 & x_32780;
assign x_32782 = x_32778 & x_32781;
assign x_32783 = x_1490 & x_1491;
assign x_32784 = x_1492 & x_1493;
assign x_32785 = x_32783 & x_32784;
assign x_32786 = x_1494 & x_1495;
assign x_32787 = x_1496 & x_1497;
assign x_32788 = x_32786 & x_32787;
assign x_32789 = x_32785 & x_32788;
assign x_32790 = x_32782 & x_32789;
assign x_32791 = x_32776 & x_32790;
assign x_32792 = x_1499 & x_1500;
assign x_32793 = x_1498 & x_32792;
assign x_32794 = x_1501 & x_1502;
assign x_32795 = x_1503 & x_1504;
assign x_32796 = x_32794 & x_32795;
assign x_32797 = x_32793 & x_32796;
assign x_32798 = x_1505 & x_1506;
assign x_32799 = x_1507 & x_1508;
assign x_32800 = x_32798 & x_32799;
assign x_32801 = x_1509 & x_1510;
assign x_32802 = x_1511 & x_1512;
assign x_32803 = x_32801 & x_32802;
assign x_32804 = x_32800 & x_32803;
assign x_32805 = x_32797 & x_32804;
assign x_32806 = x_1513 & x_1514;
assign x_32807 = x_1515 & x_1516;
assign x_32808 = x_32806 & x_32807;
assign x_32809 = x_1517 & x_1518;
assign x_32810 = x_1519 & x_1520;
assign x_32811 = x_32809 & x_32810;
assign x_32812 = x_32808 & x_32811;
assign x_32813 = x_1521 & x_1522;
assign x_32814 = x_1523 & x_1524;
assign x_32815 = x_32813 & x_32814;
assign x_32816 = x_1525 & x_1526;
assign x_32817 = x_1527 & x_1528;
assign x_32818 = x_32816 & x_32817;
assign x_32819 = x_32815 & x_32818;
assign x_32820 = x_32812 & x_32819;
assign x_32821 = x_32805 & x_32820;
assign x_32822 = x_32791 & x_32821;
assign x_32823 = x_1530 & x_1531;
assign x_32824 = x_1529 & x_32823;
assign x_32825 = x_1532 & x_1533;
assign x_32826 = x_1534 & x_1535;
assign x_32827 = x_32825 & x_32826;
assign x_32828 = x_32824 & x_32827;
assign x_32829 = x_1536 & x_1537;
assign x_32830 = x_1538 & x_1539;
assign x_32831 = x_32829 & x_32830;
assign x_32832 = x_1540 & x_1541;
assign x_32833 = x_1542 & x_1543;
assign x_32834 = x_32832 & x_32833;
assign x_32835 = x_32831 & x_32834;
assign x_32836 = x_32828 & x_32835;
assign x_32837 = x_1545 & x_1546;
assign x_32838 = x_1544 & x_32837;
assign x_32839 = x_1547 & x_1548;
assign x_32840 = x_1549 & x_1550;
assign x_32841 = x_32839 & x_32840;
assign x_32842 = x_32838 & x_32841;
assign x_32843 = x_1551 & x_1552;
assign x_32844 = x_1553 & x_1554;
assign x_32845 = x_32843 & x_32844;
assign x_32846 = x_1555 & x_1556;
assign x_32847 = x_1557 & x_1558;
assign x_32848 = x_32846 & x_32847;
assign x_32849 = x_32845 & x_32848;
assign x_32850 = x_32842 & x_32849;
assign x_32851 = x_32836 & x_32850;
assign x_32852 = x_1560 & x_1561;
assign x_32853 = x_1559 & x_32852;
assign x_32854 = x_1562 & x_1563;
assign x_32855 = x_1564 & x_1565;
assign x_32856 = x_32854 & x_32855;
assign x_32857 = x_32853 & x_32856;
assign x_32858 = x_1566 & x_1567;
assign x_32859 = x_1568 & x_1569;
assign x_32860 = x_32858 & x_32859;
assign x_32861 = x_1570 & x_1571;
assign x_32862 = x_1572 & x_1573;
assign x_32863 = x_32861 & x_32862;
assign x_32864 = x_32860 & x_32863;
assign x_32865 = x_32857 & x_32864;
assign x_32866 = x_1574 & x_1575;
assign x_32867 = x_1576 & x_1577;
assign x_32868 = x_32866 & x_32867;
assign x_32869 = x_1578 & x_1579;
assign x_32870 = x_1580 & x_1581;
assign x_32871 = x_32869 & x_32870;
assign x_32872 = x_32868 & x_32871;
assign x_32873 = x_1582 & x_1583;
assign x_32874 = x_1584 & x_1585;
assign x_32875 = x_32873 & x_32874;
assign x_32876 = x_1586 & x_1587;
assign x_32877 = x_1588 & x_1589;
assign x_32878 = x_32876 & x_32877;
assign x_32879 = x_32875 & x_32878;
assign x_32880 = x_32872 & x_32879;
assign x_32881 = x_32865 & x_32880;
assign x_32882 = x_32851 & x_32881;
assign x_32883 = x_32822 & x_32882;
assign x_32884 = x_1591 & x_1592;
assign x_32885 = x_1590 & x_32884;
assign x_32886 = x_1593 & x_1594;
assign x_32887 = x_1595 & x_1596;
assign x_32888 = x_32886 & x_32887;
assign x_32889 = x_32885 & x_32888;
assign x_32890 = x_1597 & x_1598;
assign x_32891 = x_1599 & x_1600;
assign x_32892 = x_32890 & x_32891;
assign x_32893 = x_1601 & x_1602;
assign x_32894 = x_1603 & x_1604;
assign x_32895 = x_32893 & x_32894;
assign x_32896 = x_32892 & x_32895;
assign x_32897 = x_32889 & x_32896;
assign x_32898 = x_1606 & x_1607;
assign x_32899 = x_1605 & x_32898;
assign x_32900 = x_1608 & x_1609;
assign x_32901 = x_1610 & x_1611;
assign x_32902 = x_32900 & x_32901;
assign x_32903 = x_32899 & x_32902;
assign x_32904 = x_1612 & x_1613;
assign x_32905 = x_1614 & x_1615;
assign x_32906 = x_32904 & x_32905;
assign x_32907 = x_1616 & x_1617;
assign x_32908 = x_1618 & x_1619;
assign x_32909 = x_32907 & x_32908;
assign x_32910 = x_32906 & x_32909;
assign x_32911 = x_32903 & x_32910;
assign x_32912 = x_32897 & x_32911;
assign x_32913 = x_1621 & x_1622;
assign x_32914 = x_1620 & x_32913;
assign x_32915 = x_1623 & x_1624;
assign x_32916 = x_1625 & x_1626;
assign x_32917 = x_32915 & x_32916;
assign x_32918 = x_32914 & x_32917;
assign x_32919 = x_1627 & x_1628;
assign x_32920 = x_1629 & x_1630;
assign x_32921 = x_32919 & x_32920;
assign x_32922 = x_1631 & x_1632;
assign x_32923 = x_1633 & x_1634;
assign x_32924 = x_32922 & x_32923;
assign x_32925 = x_32921 & x_32924;
assign x_32926 = x_32918 & x_32925;
assign x_32927 = x_1635 & x_1636;
assign x_32928 = x_1637 & x_1638;
assign x_32929 = x_32927 & x_32928;
assign x_32930 = x_1639 & x_1640;
assign x_32931 = x_1641 & x_1642;
assign x_32932 = x_32930 & x_32931;
assign x_32933 = x_32929 & x_32932;
assign x_32934 = x_1643 & x_1644;
assign x_32935 = x_1645 & x_1646;
assign x_32936 = x_32934 & x_32935;
assign x_32937 = x_1647 & x_1648;
assign x_32938 = x_1649 & x_1650;
assign x_32939 = x_32937 & x_32938;
assign x_32940 = x_32936 & x_32939;
assign x_32941 = x_32933 & x_32940;
assign x_32942 = x_32926 & x_32941;
assign x_32943 = x_32912 & x_32942;
assign x_32944 = x_1652 & x_1653;
assign x_32945 = x_1651 & x_32944;
assign x_32946 = x_1654 & x_1655;
assign x_32947 = x_1656 & x_1657;
assign x_32948 = x_32946 & x_32947;
assign x_32949 = x_32945 & x_32948;
assign x_32950 = x_1658 & x_1659;
assign x_32951 = x_1660 & x_1661;
assign x_32952 = x_32950 & x_32951;
assign x_32953 = x_1662 & x_1663;
assign x_32954 = x_1664 & x_1665;
assign x_32955 = x_32953 & x_32954;
assign x_32956 = x_32952 & x_32955;
assign x_32957 = x_32949 & x_32956;
assign x_32958 = x_1667 & x_1668;
assign x_32959 = x_1666 & x_32958;
assign x_32960 = x_1669 & x_1670;
assign x_32961 = x_1671 & x_1672;
assign x_32962 = x_32960 & x_32961;
assign x_32963 = x_32959 & x_32962;
assign x_32964 = x_1673 & x_1674;
assign x_32965 = x_1675 & x_1676;
assign x_32966 = x_32964 & x_32965;
assign x_32967 = x_1677 & x_1678;
assign x_32968 = x_1679 & x_1680;
assign x_32969 = x_32967 & x_32968;
assign x_32970 = x_32966 & x_32969;
assign x_32971 = x_32963 & x_32970;
assign x_32972 = x_32957 & x_32971;
assign x_32973 = x_1682 & x_1683;
assign x_32974 = x_1681 & x_32973;
assign x_32975 = x_1684 & x_1685;
assign x_32976 = x_1686 & x_1687;
assign x_32977 = x_32975 & x_32976;
assign x_32978 = x_32974 & x_32977;
assign x_32979 = x_1688 & x_1689;
assign x_32980 = x_1690 & x_1691;
assign x_32981 = x_32979 & x_32980;
assign x_32982 = x_1692 & x_1693;
assign x_32983 = x_1694 & x_1695;
assign x_32984 = x_32982 & x_32983;
assign x_32985 = x_32981 & x_32984;
assign x_32986 = x_32978 & x_32985;
assign x_32987 = x_1696 & x_1697;
assign x_32988 = x_1698 & x_1699;
assign x_32989 = x_32987 & x_32988;
assign x_32990 = x_1700 & x_1701;
assign x_32991 = x_1702 & x_1703;
assign x_32992 = x_32990 & x_32991;
assign x_32993 = x_32989 & x_32992;
assign x_32994 = x_1704 & x_1705;
assign x_32995 = x_1706 & x_1707;
assign x_32996 = x_32994 & x_32995;
assign x_32997 = x_1708 & x_1709;
assign x_32998 = x_1710 & x_1711;
assign x_32999 = x_32997 & x_32998;
assign x_33000 = x_32996 & x_32999;
assign x_33001 = x_32993 & x_33000;
assign x_33002 = x_32986 & x_33001;
assign x_33003 = x_32972 & x_33002;
assign x_33004 = x_32943 & x_33003;
assign x_33005 = x_32883 & x_33004;
assign x_33006 = x_1713 & x_1714;
assign x_33007 = x_1712 & x_33006;
assign x_33008 = x_1715 & x_1716;
assign x_33009 = x_1717 & x_1718;
assign x_33010 = x_33008 & x_33009;
assign x_33011 = x_33007 & x_33010;
assign x_33012 = x_1719 & x_1720;
assign x_33013 = x_1721 & x_1722;
assign x_33014 = x_33012 & x_33013;
assign x_33015 = x_1723 & x_1724;
assign x_33016 = x_1725 & x_1726;
assign x_33017 = x_33015 & x_33016;
assign x_33018 = x_33014 & x_33017;
assign x_33019 = x_33011 & x_33018;
assign x_33020 = x_1728 & x_1729;
assign x_33021 = x_1727 & x_33020;
assign x_33022 = x_1730 & x_1731;
assign x_33023 = x_1732 & x_1733;
assign x_33024 = x_33022 & x_33023;
assign x_33025 = x_33021 & x_33024;
assign x_33026 = x_1734 & x_1735;
assign x_33027 = x_1736 & x_1737;
assign x_33028 = x_33026 & x_33027;
assign x_33029 = x_1738 & x_1739;
assign x_33030 = x_1740 & x_1741;
assign x_33031 = x_33029 & x_33030;
assign x_33032 = x_33028 & x_33031;
assign x_33033 = x_33025 & x_33032;
assign x_33034 = x_33019 & x_33033;
assign x_33035 = x_1743 & x_1744;
assign x_33036 = x_1742 & x_33035;
assign x_33037 = x_1745 & x_1746;
assign x_33038 = x_1747 & x_1748;
assign x_33039 = x_33037 & x_33038;
assign x_33040 = x_33036 & x_33039;
assign x_33041 = x_1749 & x_1750;
assign x_33042 = x_1751 & x_1752;
assign x_33043 = x_33041 & x_33042;
assign x_33044 = x_1753 & x_1754;
assign x_33045 = x_1755 & x_1756;
assign x_33046 = x_33044 & x_33045;
assign x_33047 = x_33043 & x_33046;
assign x_33048 = x_33040 & x_33047;
assign x_33049 = x_1757 & x_1758;
assign x_33050 = x_1759 & x_1760;
assign x_33051 = x_33049 & x_33050;
assign x_33052 = x_1761 & x_1762;
assign x_33053 = x_1763 & x_1764;
assign x_33054 = x_33052 & x_33053;
assign x_33055 = x_33051 & x_33054;
assign x_33056 = x_1765 & x_1766;
assign x_33057 = x_1767 & x_1768;
assign x_33058 = x_33056 & x_33057;
assign x_33059 = x_1769 & x_1770;
assign x_33060 = x_1771 & x_1772;
assign x_33061 = x_33059 & x_33060;
assign x_33062 = x_33058 & x_33061;
assign x_33063 = x_33055 & x_33062;
assign x_33064 = x_33048 & x_33063;
assign x_33065 = x_33034 & x_33064;
assign x_33066 = x_1774 & x_1775;
assign x_33067 = x_1773 & x_33066;
assign x_33068 = x_1776 & x_1777;
assign x_33069 = x_1778 & x_1779;
assign x_33070 = x_33068 & x_33069;
assign x_33071 = x_33067 & x_33070;
assign x_33072 = x_1780 & x_1781;
assign x_33073 = x_1782 & x_1783;
assign x_33074 = x_33072 & x_33073;
assign x_33075 = x_1784 & x_1785;
assign x_33076 = x_1786 & x_1787;
assign x_33077 = x_33075 & x_33076;
assign x_33078 = x_33074 & x_33077;
assign x_33079 = x_33071 & x_33078;
assign x_33080 = x_1789 & x_1790;
assign x_33081 = x_1788 & x_33080;
assign x_33082 = x_1791 & x_1792;
assign x_33083 = x_1793 & x_1794;
assign x_33084 = x_33082 & x_33083;
assign x_33085 = x_33081 & x_33084;
assign x_33086 = x_1795 & x_1796;
assign x_33087 = x_1797 & x_1798;
assign x_33088 = x_33086 & x_33087;
assign x_33089 = x_1799 & x_1800;
assign x_33090 = x_1801 & x_1802;
assign x_33091 = x_33089 & x_33090;
assign x_33092 = x_33088 & x_33091;
assign x_33093 = x_33085 & x_33092;
assign x_33094 = x_33079 & x_33093;
assign x_33095 = x_1804 & x_1805;
assign x_33096 = x_1803 & x_33095;
assign x_33097 = x_1806 & x_1807;
assign x_33098 = x_1808 & x_1809;
assign x_33099 = x_33097 & x_33098;
assign x_33100 = x_33096 & x_33099;
assign x_33101 = x_1810 & x_1811;
assign x_33102 = x_1812 & x_1813;
assign x_33103 = x_33101 & x_33102;
assign x_33104 = x_1814 & x_1815;
assign x_33105 = x_1816 & x_1817;
assign x_33106 = x_33104 & x_33105;
assign x_33107 = x_33103 & x_33106;
assign x_33108 = x_33100 & x_33107;
assign x_33109 = x_1818 & x_1819;
assign x_33110 = x_1820 & x_1821;
assign x_33111 = x_33109 & x_33110;
assign x_33112 = x_1822 & x_1823;
assign x_33113 = x_1824 & x_1825;
assign x_33114 = x_33112 & x_33113;
assign x_33115 = x_33111 & x_33114;
assign x_33116 = x_1826 & x_1827;
assign x_33117 = x_1828 & x_1829;
assign x_33118 = x_33116 & x_33117;
assign x_33119 = x_1830 & x_1831;
assign x_33120 = x_1832 & x_1833;
assign x_33121 = x_33119 & x_33120;
assign x_33122 = x_33118 & x_33121;
assign x_33123 = x_33115 & x_33122;
assign x_33124 = x_33108 & x_33123;
assign x_33125 = x_33094 & x_33124;
assign x_33126 = x_33065 & x_33125;
assign x_33127 = x_1835 & x_1836;
assign x_33128 = x_1834 & x_33127;
assign x_33129 = x_1837 & x_1838;
assign x_33130 = x_1839 & x_1840;
assign x_33131 = x_33129 & x_33130;
assign x_33132 = x_33128 & x_33131;
assign x_33133 = x_1841 & x_1842;
assign x_33134 = x_1843 & x_1844;
assign x_33135 = x_33133 & x_33134;
assign x_33136 = x_1845 & x_1846;
assign x_33137 = x_1847 & x_1848;
assign x_33138 = x_33136 & x_33137;
assign x_33139 = x_33135 & x_33138;
assign x_33140 = x_33132 & x_33139;
assign x_33141 = x_1850 & x_1851;
assign x_33142 = x_1849 & x_33141;
assign x_33143 = x_1852 & x_1853;
assign x_33144 = x_1854 & x_1855;
assign x_33145 = x_33143 & x_33144;
assign x_33146 = x_33142 & x_33145;
assign x_33147 = x_1856 & x_1857;
assign x_33148 = x_1858 & x_1859;
assign x_33149 = x_33147 & x_33148;
assign x_33150 = x_1860 & x_1861;
assign x_33151 = x_1862 & x_1863;
assign x_33152 = x_33150 & x_33151;
assign x_33153 = x_33149 & x_33152;
assign x_33154 = x_33146 & x_33153;
assign x_33155 = x_33140 & x_33154;
assign x_33156 = x_1865 & x_1866;
assign x_33157 = x_1864 & x_33156;
assign x_33158 = x_1867 & x_1868;
assign x_33159 = x_1869 & x_1870;
assign x_33160 = x_33158 & x_33159;
assign x_33161 = x_33157 & x_33160;
assign x_33162 = x_1871 & x_1872;
assign x_33163 = x_1873 & x_1874;
assign x_33164 = x_33162 & x_33163;
assign x_33165 = x_1875 & x_1876;
assign x_33166 = x_1877 & x_1878;
assign x_33167 = x_33165 & x_33166;
assign x_33168 = x_33164 & x_33167;
assign x_33169 = x_33161 & x_33168;
assign x_33170 = x_1879 & x_1880;
assign x_33171 = x_1881 & x_1882;
assign x_33172 = x_33170 & x_33171;
assign x_33173 = x_1883 & x_1884;
assign x_33174 = x_1885 & x_1886;
assign x_33175 = x_33173 & x_33174;
assign x_33176 = x_33172 & x_33175;
assign x_33177 = x_1887 & x_1888;
assign x_33178 = x_1889 & x_1890;
assign x_33179 = x_33177 & x_33178;
assign x_33180 = x_1891 & x_1892;
assign x_33181 = x_1893 & x_1894;
assign x_33182 = x_33180 & x_33181;
assign x_33183 = x_33179 & x_33182;
assign x_33184 = x_33176 & x_33183;
assign x_33185 = x_33169 & x_33184;
assign x_33186 = x_33155 & x_33185;
assign x_33187 = x_1896 & x_1897;
assign x_33188 = x_1895 & x_33187;
assign x_33189 = x_1898 & x_1899;
assign x_33190 = x_1900 & x_1901;
assign x_33191 = x_33189 & x_33190;
assign x_33192 = x_33188 & x_33191;
assign x_33193 = x_1902 & x_1903;
assign x_33194 = x_1904 & x_1905;
assign x_33195 = x_33193 & x_33194;
assign x_33196 = x_1906 & x_1907;
assign x_33197 = x_1908 & x_1909;
assign x_33198 = x_33196 & x_33197;
assign x_33199 = x_33195 & x_33198;
assign x_33200 = x_33192 & x_33199;
assign x_33201 = x_1910 & x_1911;
assign x_33202 = x_1912 & x_1913;
assign x_33203 = x_33201 & x_33202;
assign x_33204 = x_1914 & x_1915;
assign x_33205 = x_1916 & x_1917;
assign x_33206 = x_33204 & x_33205;
assign x_33207 = x_33203 & x_33206;
assign x_33208 = x_1918 & x_1919;
assign x_33209 = x_1920 & x_1921;
assign x_33210 = x_33208 & x_33209;
assign x_33211 = x_1922 & x_1923;
assign x_33212 = x_1924 & x_1925;
assign x_33213 = x_33211 & x_33212;
assign x_33214 = x_33210 & x_33213;
assign x_33215 = x_33207 & x_33214;
assign x_33216 = x_33200 & x_33215;
assign x_33217 = x_1927 & x_1928;
assign x_33218 = x_1926 & x_33217;
assign x_33219 = x_1929 & x_1930;
assign x_33220 = x_1931 & x_1932;
assign x_33221 = x_33219 & x_33220;
assign x_33222 = x_33218 & x_33221;
assign x_33223 = x_1933 & x_1934;
assign x_33224 = x_1935 & x_1936;
assign x_33225 = x_33223 & x_33224;
assign x_33226 = x_1937 & x_1938;
assign x_33227 = x_1939 & x_1940;
assign x_33228 = x_33226 & x_33227;
assign x_33229 = x_33225 & x_33228;
assign x_33230 = x_33222 & x_33229;
assign x_33231 = x_1941 & x_1942;
assign x_33232 = x_1943 & x_1944;
assign x_33233 = x_33231 & x_33232;
assign x_33234 = x_1945 & x_1946;
assign x_33235 = x_1947 & x_1948;
assign x_33236 = x_33234 & x_33235;
assign x_33237 = x_33233 & x_33236;
assign x_33238 = x_1949 & x_1950;
assign x_33239 = x_1951 & x_1952;
assign x_33240 = x_33238 & x_33239;
assign x_33241 = x_1953 & x_1954;
assign x_33242 = x_1955 & x_1956;
assign x_33243 = x_33241 & x_33242;
assign x_33244 = x_33240 & x_33243;
assign x_33245 = x_33237 & x_33244;
assign x_33246 = x_33230 & x_33245;
assign x_33247 = x_33216 & x_33246;
assign x_33248 = x_33186 & x_33247;
assign x_33249 = x_33126 & x_33248;
assign x_33250 = x_33005 & x_33249;
assign x_33251 = x_32762 & x_33250;
assign x_33252 = x_32274 & x_33251;
assign x_33253 = x_1958 & x_1959;
assign x_33254 = x_1957 & x_33253;
assign x_33255 = x_1960 & x_1961;
assign x_33256 = x_1962 & x_1963;
assign x_33257 = x_33255 & x_33256;
assign x_33258 = x_33254 & x_33257;
assign x_33259 = x_1964 & x_1965;
assign x_33260 = x_1966 & x_1967;
assign x_33261 = x_33259 & x_33260;
assign x_33262 = x_1968 & x_1969;
assign x_33263 = x_1970 & x_1971;
assign x_33264 = x_33262 & x_33263;
assign x_33265 = x_33261 & x_33264;
assign x_33266 = x_33258 & x_33265;
assign x_33267 = x_1973 & x_1974;
assign x_33268 = x_1972 & x_33267;
assign x_33269 = x_1975 & x_1976;
assign x_33270 = x_1977 & x_1978;
assign x_33271 = x_33269 & x_33270;
assign x_33272 = x_33268 & x_33271;
assign x_33273 = x_1979 & x_1980;
assign x_33274 = x_1981 & x_1982;
assign x_33275 = x_33273 & x_33274;
assign x_33276 = x_1983 & x_1984;
assign x_33277 = x_1985 & x_1986;
assign x_33278 = x_33276 & x_33277;
assign x_33279 = x_33275 & x_33278;
assign x_33280 = x_33272 & x_33279;
assign x_33281 = x_33266 & x_33280;
assign x_33282 = x_1988 & x_1989;
assign x_33283 = x_1987 & x_33282;
assign x_33284 = x_1990 & x_1991;
assign x_33285 = x_1992 & x_1993;
assign x_33286 = x_33284 & x_33285;
assign x_33287 = x_33283 & x_33286;
assign x_33288 = x_1994 & x_1995;
assign x_33289 = x_1996 & x_1997;
assign x_33290 = x_33288 & x_33289;
assign x_33291 = x_1998 & x_1999;
assign x_33292 = x_2000 & x_2001;
assign x_33293 = x_33291 & x_33292;
assign x_33294 = x_33290 & x_33293;
assign x_33295 = x_33287 & x_33294;
assign x_33296 = x_2002 & x_2003;
assign x_33297 = x_2004 & x_2005;
assign x_33298 = x_33296 & x_33297;
assign x_33299 = x_2006 & x_2007;
assign x_33300 = x_2008 & x_2009;
assign x_33301 = x_33299 & x_33300;
assign x_33302 = x_33298 & x_33301;
assign x_33303 = x_2010 & x_2011;
assign x_33304 = x_2012 & x_2013;
assign x_33305 = x_33303 & x_33304;
assign x_33306 = x_2014 & x_2015;
assign x_33307 = x_2016 & x_2017;
assign x_33308 = x_33306 & x_33307;
assign x_33309 = x_33305 & x_33308;
assign x_33310 = x_33302 & x_33309;
assign x_33311 = x_33295 & x_33310;
assign x_33312 = x_33281 & x_33311;
assign x_33313 = x_2019 & x_2020;
assign x_33314 = x_2018 & x_33313;
assign x_33315 = x_2021 & x_2022;
assign x_33316 = x_2023 & x_2024;
assign x_33317 = x_33315 & x_33316;
assign x_33318 = x_33314 & x_33317;
assign x_33319 = x_2025 & x_2026;
assign x_33320 = x_2027 & x_2028;
assign x_33321 = x_33319 & x_33320;
assign x_33322 = x_2029 & x_2030;
assign x_33323 = x_2031 & x_2032;
assign x_33324 = x_33322 & x_33323;
assign x_33325 = x_33321 & x_33324;
assign x_33326 = x_33318 & x_33325;
assign x_33327 = x_2034 & x_2035;
assign x_33328 = x_2033 & x_33327;
assign x_33329 = x_2036 & x_2037;
assign x_33330 = x_2038 & x_2039;
assign x_33331 = x_33329 & x_33330;
assign x_33332 = x_33328 & x_33331;
assign x_33333 = x_2040 & x_2041;
assign x_33334 = x_2042 & x_2043;
assign x_33335 = x_33333 & x_33334;
assign x_33336 = x_2044 & x_2045;
assign x_33337 = x_2046 & x_2047;
assign x_33338 = x_33336 & x_33337;
assign x_33339 = x_33335 & x_33338;
assign x_33340 = x_33332 & x_33339;
assign x_33341 = x_33326 & x_33340;
assign x_33342 = x_2049 & x_2050;
assign x_33343 = x_2048 & x_33342;
assign x_33344 = x_2051 & x_2052;
assign x_33345 = x_2053 & x_2054;
assign x_33346 = x_33344 & x_33345;
assign x_33347 = x_33343 & x_33346;
assign x_33348 = x_2055 & x_2056;
assign x_33349 = x_2057 & x_2058;
assign x_33350 = x_33348 & x_33349;
assign x_33351 = x_2059 & x_2060;
assign x_33352 = x_2061 & x_2062;
assign x_33353 = x_33351 & x_33352;
assign x_33354 = x_33350 & x_33353;
assign x_33355 = x_33347 & x_33354;
assign x_33356 = x_2063 & x_2064;
assign x_33357 = x_2065 & x_2066;
assign x_33358 = x_33356 & x_33357;
assign x_33359 = x_2067 & x_2068;
assign x_33360 = x_2069 & x_2070;
assign x_33361 = x_33359 & x_33360;
assign x_33362 = x_33358 & x_33361;
assign x_33363 = x_2071 & x_2072;
assign x_33364 = x_2073 & x_2074;
assign x_33365 = x_33363 & x_33364;
assign x_33366 = x_2075 & x_2076;
assign x_33367 = x_2077 & x_2078;
assign x_33368 = x_33366 & x_33367;
assign x_33369 = x_33365 & x_33368;
assign x_33370 = x_33362 & x_33369;
assign x_33371 = x_33355 & x_33370;
assign x_33372 = x_33341 & x_33371;
assign x_33373 = x_33312 & x_33372;
assign x_33374 = x_2080 & x_2081;
assign x_33375 = x_2079 & x_33374;
assign x_33376 = x_2082 & x_2083;
assign x_33377 = x_2084 & x_2085;
assign x_33378 = x_33376 & x_33377;
assign x_33379 = x_33375 & x_33378;
assign x_33380 = x_2086 & x_2087;
assign x_33381 = x_2088 & x_2089;
assign x_33382 = x_33380 & x_33381;
assign x_33383 = x_2090 & x_2091;
assign x_33384 = x_2092 & x_2093;
assign x_33385 = x_33383 & x_33384;
assign x_33386 = x_33382 & x_33385;
assign x_33387 = x_33379 & x_33386;
assign x_33388 = x_2095 & x_2096;
assign x_33389 = x_2094 & x_33388;
assign x_33390 = x_2097 & x_2098;
assign x_33391 = x_2099 & x_2100;
assign x_33392 = x_33390 & x_33391;
assign x_33393 = x_33389 & x_33392;
assign x_33394 = x_2101 & x_2102;
assign x_33395 = x_2103 & x_2104;
assign x_33396 = x_33394 & x_33395;
assign x_33397 = x_2105 & x_2106;
assign x_33398 = x_2107 & x_2108;
assign x_33399 = x_33397 & x_33398;
assign x_33400 = x_33396 & x_33399;
assign x_33401 = x_33393 & x_33400;
assign x_33402 = x_33387 & x_33401;
assign x_33403 = x_2110 & x_2111;
assign x_33404 = x_2109 & x_33403;
assign x_33405 = x_2112 & x_2113;
assign x_33406 = x_2114 & x_2115;
assign x_33407 = x_33405 & x_33406;
assign x_33408 = x_33404 & x_33407;
assign x_33409 = x_2116 & x_2117;
assign x_33410 = x_2118 & x_2119;
assign x_33411 = x_33409 & x_33410;
assign x_33412 = x_2120 & x_2121;
assign x_33413 = x_2122 & x_2123;
assign x_33414 = x_33412 & x_33413;
assign x_33415 = x_33411 & x_33414;
assign x_33416 = x_33408 & x_33415;
assign x_33417 = x_2124 & x_2125;
assign x_33418 = x_2126 & x_2127;
assign x_33419 = x_33417 & x_33418;
assign x_33420 = x_2128 & x_2129;
assign x_33421 = x_2130 & x_2131;
assign x_33422 = x_33420 & x_33421;
assign x_33423 = x_33419 & x_33422;
assign x_33424 = x_2132 & x_2133;
assign x_33425 = x_2134 & x_2135;
assign x_33426 = x_33424 & x_33425;
assign x_33427 = x_2136 & x_2137;
assign x_33428 = x_2138 & x_2139;
assign x_33429 = x_33427 & x_33428;
assign x_33430 = x_33426 & x_33429;
assign x_33431 = x_33423 & x_33430;
assign x_33432 = x_33416 & x_33431;
assign x_33433 = x_33402 & x_33432;
assign x_33434 = x_2141 & x_2142;
assign x_33435 = x_2140 & x_33434;
assign x_33436 = x_2143 & x_2144;
assign x_33437 = x_2145 & x_2146;
assign x_33438 = x_33436 & x_33437;
assign x_33439 = x_33435 & x_33438;
assign x_33440 = x_2147 & x_2148;
assign x_33441 = x_2149 & x_2150;
assign x_33442 = x_33440 & x_33441;
assign x_33443 = x_2151 & x_2152;
assign x_33444 = x_2153 & x_2154;
assign x_33445 = x_33443 & x_33444;
assign x_33446 = x_33442 & x_33445;
assign x_33447 = x_33439 & x_33446;
assign x_33448 = x_2156 & x_2157;
assign x_33449 = x_2155 & x_33448;
assign x_33450 = x_2158 & x_2159;
assign x_33451 = x_2160 & x_2161;
assign x_33452 = x_33450 & x_33451;
assign x_33453 = x_33449 & x_33452;
assign x_33454 = x_2162 & x_2163;
assign x_33455 = x_2164 & x_2165;
assign x_33456 = x_33454 & x_33455;
assign x_33457 = x_2166 & x_2167;
assign x_33458 = x_2168 & x_2169;
assign x_33459 = x_33457 & x_33458;
assign x_33460 = x_33456 & x_33459;
assign x_33461 = x_33453 & x_33460;
assign x_33462 = x_33447 & x_33461;
assign x_33463 = x_2171 & x_2172;
assign x_33464 = x_2170 & x_33463;
assign x_33465 = x_2173 & x_2174;
assign x_33466 = x_2175 & x_2176;
assign x_33467 = x_33465 & x_33466;
assign x_33468 = x_33464 & x_33467;
assign x_33469 = x_2177 & x_2178;
assign x_33470 = x_2179 & x_2180;
assign x_33471 = x_33469 & x_33470;
assign x_33472 = x_2181 & x_2182;
assign x_33473 = x_2183 & x_2184;
assign x_33474 = x_33472 & x_33473;
assign x_33475 = x_33471 & x_33474;
assign x_33476 = x_33468 & x_33475;
assign x_33477 = x_2185 & x_2186;
assign x_33478 = x_2187 & x_2188;
assign x_33479 = x_33477 & x_33478;
assign x_33480 = x_2189 & x_2190;
assign x_33481 = x_2191 & x_2192;
assign x_33482 = x_33480 & x_33481;
assign x_33483 = x_33479 & x_33482;
assign x_33484 = x_2193 & x_2194;
assign x_33485 = x_2195 & x_2196;
assign x_33486 = x_33484 & x_33485;
assign x_33487 = x_2197 & x_2198;
assign x_33488 = x_2199 & x_2200;
assign x_33489 = x_33487 & x_33488;
assign x_33490 = x_33486 & x_33489;
assign x_33491 = x_33483 & x_33490;
assign x_33492 = x_33476 & x_33491;
assign x_33493 = x_33462 & x_33492;
assign x_33494 = x_33433 & x_33493;
assign x_33495 = x_33373 & x_33494;
assign x_33496 = x_2202 & x_2203;
assign x_33497 = x_2201 & x_33496;
assign x_33498 = x_2204 & x_2205;
assign x_33499 = x_2206 & x_2207;
assign x_33500 = x_33498 & x_33499;
assign x_33501 = x_33497 & x_33500;
assign x_33502 = x_2208 & x_2209;
assign x_33503 = x_2210 & x_2211;
assign x_33504 = x_33502 & x_33503;
assign x_33505 = x_2212 & x_2213;
assign x_33506 = x_2214 & x_2215;
assign x_33507 = x_33505 & x_33506;
assign x_33508 = x_33504 & x_33507;
assign x_33509 = x_33501 & x_33508;
assign x_33510 = x_2217 & x_2218;
assign x_33511 = x_2216 & x_33510;
assign x_33512 = x_2219 & x_2220;
assign x_33513 = x_2221 & x_2222;
assign x_33514 = x_33512 & x_33513;
assign x_33515 = x_33511 & x_33514;
assign x_33516 = x_2223 & x_2224;
assign x_33517 = x_2225 & x_2226;
assign x_33518 = x_33516 & x_33517;
assign x_33519 = x_2227 & x_2228;
assign x_33520 = x_2229 & x_2230;
assign x_33521 = x_33519 & x_33520;
assign x_33522 = x_33518 & x_33521;
assign x_33523 = x_33515 & x_33522;
assign x_33524 = x_33509 & x_33523;
assign x_33525 = x_2232 & x_2233;
assign x_33526 = x_2231 & x_33525;
assign x_33527 = x_2234 & x_2235;
assign x_33528 = x_2236 & x_2237;
assign x_33529 = x_33527 & x_33528;
assign x_33530 = x_33526 & x_33529;
assign x_33531 = x_2238 & x_2239;
assign x_33532 = x_2240 & x_2241;
assign x_33533 = x_33531 & x_33532;
assign x_33534 = x_2242 & x_2243;
assign x_33535 = x_2244 & x_2245;
assign x_33536 = x_33534 & x_33535;
assign x_33537 = x_33533 & x_33536;
assign x_33538 = x_33530 & x_33537;
assign x_33539 = x_2246 & x_2247;
assign x_33540 = x_2248 & x_2249;
assign x_33541 = x_33539 & x_33540;
assign x_33542 = x_2250 & x_2251;
assign x_33543 = x_2252 & x_2253;
assign x_33544 = x_33542 & x_33543;
assign x_33545 = x_33541 & x_33544;
assign x_33546 = x_2254 & x_2255;
assign x_33547 = x_2256 & x_2257;
assign x_33548 = x_33546 & x_33547;
assign x_33549 = x_2258 & x_2259;
assign x_33550 = x_2260 & x_2261;
assign x_33551 = x_33549 & x_33550;
assign x_33552 = x_33548 & x_33551;
assign x_33553 = x_33545 & x_33552;
assign x_33554 = x_33538 & x_33553;
assign x_33555 = x_33524 & x_33554;
assign x_33556 = x_2263 & x_2264;
assign x_33557 = x_2262 & x_33556;
assign x_33558 = x_2265 & x_2266;
assign x_33559 = x_2267 & x_2268;
assign x_33560 = x_33558 & x_33559;
assign x_33561 = x_33557 & x_33560;
assign x_33562 = x_2269 & x_2270;
assign x_33563 = x_2271 & x_2272;
assign x_33564 = x_33562 & x_33563;
assign x_33565 = x_2273 & x_2274;
assign x_33566 = x_2275 & x_2276;
assign x_33567 = x_33565 & x_33566;
assign x_33568 = x_33564 & x_33567;
assign x_33569 = x_33561 & x_33568;
assign x_33570 = x_2278 & x_2279;
assign x_33571 = x_2277 & x_33570;
assign x_33572 = x_2280 & x_2281;
assign x_33573 = x_2282 & x_2283;
assign x_33574 = x_33572 & x_33573;
assign x_33575 = x_33571 & x_33574;
assign x_33576 = x_2284 & x_2285;
assign x_33577 = x_2286 & x_2287;
assign x_33578 = x_33576 & x_33577;
assign x_33579 = x_2288 & x_2289;
assign x_33580 = x_2290 & x_2291;
assign x_33581 = x_33579 & x_33580;
assign x_33582 = x_33578 & x_33581;
assign x_33583 = x_33575 & x_33582;
assign x_33584 = x_33569 & x_33583;
assign x_33585 = x_2293 & x_2294;
assign x_33586 = x_2292 & x_33585;
assign x_33587 = x_2295 & x_2296;
assign x_33588 = x_2297 & x_2298;
assign x_33589 = x_33587 & x_33588;
assign x_33590 = x_33586 & x_33589;
assign x_33591 = x_2299 & x_2300;
assign x_33592 = x_2301 & x_2302;
assign x_33593 = x_33591 & x_33592;
assign x_33594 = x_2303 & x_2304;
assign x_33595 = x_2305 & x_2306;
assign x_33596 = x_33594 & x_33595;
assign x_33597 = x_33593 & x_33596;
assign x_33598 = x_33590 & x_33597;
assign x_33599 = x_2307 & x_2308;
assign x_33600 = x_2309 & x_2310;
assign x_33601 = x_33599 & x_33600;
assign x_33602 = x_2311 & x_2312;
assign x_33603 = x_2313 & x_2314;
assign x_33604 = x_33602 & x_33603;
assign x_33605 = x_33601 & x_33604;
assign x_33606 = x_2315 & x_2316;
assign x_33607 = x_2317 & x_2318;
assign x_33608 = x_33606 & x_33607;
assign x_33609 = x_2319 & x_2320;
assign x_33610 = x_2321 & x_2322;
assign x_33611 = x_33609 & x_33610;
assign x_33612 = x_33608 & x_33611;
assign x_33613 = x_33605 & x_33612;
assign x_33614 = x_33598 & x_33613;
assign x_33615 = x_33584 & x_33614;
assign x_33616 = x_33555 & x_33615;
assign x_33617 = x_2324 & x_2325;
assign x_33618 = x_2323 & x_33617;
assign x_33619 = x_2326 & x_2327;
assign x_33620 = x_2328 & x_2329;
assign x_33621 = x_33619 & x_33620;
assign x_33622 = x_33618 & x_33621;
assign x_33623 = x_2330 & x_2331;
assign x_33624 = x_2332 & x_2333;
assign x_33625 = x_33623 & x_33624;
assign x_33626 = x_2334 & x_2335;
assign x_33627 = x_2336 & x_2337;
assign x_33628 = x_33626 & x_33627;
assign x_33629 = x_33625 & x_33628;
assign x_33630 = x_33622 & x_33629;
assign x_33631 = x_2339 & x_2340;
assign x_33632 = x_2338 & x_33631;
assign x_33633 = x_2341 & x_2342;
assign x_33634 = x_2343 & x_2344;
assign x_33635 = x_33633 & x_33634;
assign x_33636 = x_33632 & x_33635;
assign x_33637 = x_2345 & x_2346;
assign x_33638 = x_2347 & x_2348;
assign x_33639 = x_33637 & x_33638;
assign x_33640 = x_2349 & x_2350;
assign x_33641 = x_2351 & x_2352;
assign x_33642 = x_33640 & x_33641;
assign x_33643 = x_33639 & x_33642;
assign x_33644 = x_33636 & x_33643;
assign x_33645 = x_33630 & x_33644;
assign x_33646 = x_2354 & x_2355;
assign x_33647 = x_2353 & x_33646;
assign x_33648 = x_2356 & x_2357;
assign x_33649 = x_2358 & x_2359;
assign x_33650 = x_33648 & x_33649;
assign x_33651 = x_33647 & x_33650;
assign x_33652 = x_2360 & x_2361;
assign x_33653 = x_2362 & x_2363;
assign x_33654 = x_33652 & x_33653;
assign x_33655 = x_2364 & x_2365;
assign x_33656 = x_2366 & x_2367;
assign x_33657 = x_33655 & x_33656;
assign x_33658 = x_33654 & x_33657;
assign x_33659 = x_33651 & x_33658;
assign x_33660 = x_2368 & x_2369;
assign x_33661 = x_2370 & x_2371;
assign x_33662 = x_33660 & x_33661;
assign x_33663 = x_2372 & x_2373;
assign x_33664 = x_2374 & x_2375;
assign x_33665 = x_33663 & x_33664;
assign x_33666 = x_33662 & x_33665;
assign x_33667 = x_2376 & x_2377;
assign x_33668 = x_2378 & x_2379;
assign x_33669 = x_33667 & x_33668;
assign x_33670 = x_2380 & x_2381;
assign x_33671 = x_2382 & x_2383;
assign x_33672 = x_33670 & x_33671;
assign x_33673 = x_33669 & x_33672;
assign x_33674 = x_33666 & x_33673;
assign x_33675 = x_33659 & x_33674;
assign x_33676 = x_33645 & x_33675;
assign x_33677 = x_2385 & x_2386;
assign x_33678 = x_2384 & x_33677;
assign x_33679 = x_2387 & x_2388;
assign x_33680 = x_2389 & x_2390;
assign x_33681 = x_33679 & x_33680;
assign x_33682 = x_33678 & x_33681;
assign x_33683 = x_2391 & x_2392;
assign x_33684 = x_2393 & x_2394;
assign x_33685 = x_33683 & x_33684;
assign x_33686 = x_2395 & x_2396;
assign x_33687 = x_2397 & x_2398;
assign x_33688 = x_33686 & x_33687;
assign x_33689 = x_33685 & x_33688;
assign x_33690 = x_33682 & x_33689;
assign x_33691 = x_2399 & x_2400;
assign x_33692 = x_2401 & x_2402;
assign x_33693 = x_33691 & x_33692;
assign x_33694 = x_2403 & x_2404;
assign x_33695 = x_2405 & x_2406;
assign x_33696 = x_33694 & x_33695;
assign x_33697 = x_33693 & x_33696;
assign x_33698 = x_2407 & x_2408;
assign x_33699 = x_2409 & x_2410;
assign x_33700 = x_33698 & x_33699;
assign x_33701 = x_2411 & x_2412;
assign x_33702 = x_2413 & x_2414;
assign x_33703 = x_33701 & x_33702;
assign x_33704 = x_33700 & x_33703;
assign x_33705 = x_33697 & x_33704;
assign x_33706 = x_33690 & x_33705;
assign x_33707 = x_2416 & x_2417;
assign x_33708 = x_2415 & x_33707;
assign x_33709 = x_2418 & x_2419;
assign x_33710 = x_2420 & x_2421;
assign x_33711 = x_33709 & x_33710;
assign x_33712 = x_33708 & x_33711;
assign x_33713 = x_2422 & x_2423;
assign x_33714 = x_2424 & x_2425;
assign x_33715 = x_33713 & x_33714;
assign x_33716 = x_2426 & x_2427;
assign x_33717 = x_2428 & x_2429;
assign x_33718 = x_33716 & x_33717;
assign x_33719 = x_33715 & x_33718;
assign x_33720 = x_33712 & x_33719;
assign x_33721 = x_2430 & x_2431;
assign x_33722 = x_2432 & x_2433;
assign x_33723 = x_33721 & x_33722;
assign x_33724 = x_2434 & x_2435;
assign x_33725 = x_2436 & x_2437;
assign x_33726 = x_33724 & x_33725;
assign x_33727 = x_33723 & x_33726;
assign x_33728 = x_2438 & x_2439;
assign x_33729 = x_2440 & x_2441;
assign x_33730 = x_33728 & x_33729;
assign x_33731 = x_2442 & x_2443;
assign x_33732 = x_2444 & x_2445;
assign x_33733 = x_33731 & x_33732;
assign x_33734 = x_33730 & x_33733;
assign x_33735 = x_33727 & x_33734;
assign x_33736 = x_33720 & x_33735;
assign x_33737 = x_33706 & x_33736;
assign x_33738 = x_33676 & x_33737;
assign x_33739 = x_33616 & x_33738;
assign x_33740 = x_33495 & x_33739;
assign x_33741 = x_2447 & x_2448;
assign x_33742 = x_2446 & x_33741;
assign x_33743 = x_2449 & x_2450;
assign x_33744 = x_2451 & x_2452;
assign x_33745 = x_33743 & x_33744;
assign x_33746 = x_33742 & x_33745;
assign x_33747 = x_2453 & x_2454;
assign x_33748 = x_2455 & x_2456;
assign x_33749 = x_33747 & x_33748;
assign x_33750 = x_2457 & x_2458;
assign x_33751 = x_2459 & x_2460;
assign x_33752 = x_33750 & x_33751;
assign x_33753 = x_33749 & x_33752;
assign x_33754 = x_33746 & x_33753;
assign x_33755 = x_2462 & x_2463;
assign x_33756 = x_2461 & x_33755;
assign x_33757 = x_2464 & x_2465;
assign x_33758 = x_2466 & x_2467;
assign x_33759 = x_33757 & x_33758;
assign x_33760 = x_33756 & x_33759;
assign x_33761 = x_2468 & x_2469;
assign x_33762 = x_2470 & x_2471;
assign x_33763 = x_33761 & x_33762;
assign x_33764 = x_2472 & x_2473;
assign x_33765 = x_2474 & x_2475;
assign x_33766 = x_33764 & x_33765;
assign x_33767 = x_33763 & x_33766;
assign x_33768 = x_33760 & x_33767;
assign x_33769 = x_33754 & x_33768;
assign x_33770 = x_2477 & x_2478;
assign x_33771 = x_2476 & x_33770;
assign x_33772 = x_2479 & x_2480;
assign x_33773 = x_2481 & x_2482;
assign x_33774 = x_33772 & x_33773;
assign x_33775 = x_33771 & x_33774;
assign x_33776 = x_2483 & x_2484;
assign x_33777 = x_2485 & x_2486;
assign x_33778 = x_33776 & x_33777;
assign x_33779 = x_2487 & x_2488;
assign x_33780 = x_2489 & x_2490;
assign x_33781 = x_33779 & x_33780;
assign x_33782 = x_33778 & x_33781;
assign x_33783 = x_33775 & x_33782;
assign x_33784 = x_2491 & x_2492;
assign x_33785 = x_2493 & x_2494;
assign x_33786 = x_33784 & x_33785;
assign x_33787 = x_2495 & x_2496;
assign x_33788 = x_2497 & x_2498;
assign x_33789 = x_33787 & x_33788;
assign x_33790 = x_33786 & x_33789;
assign x_33791 = x_2499 & x_2500;
assign x_33792 = x_2501 & x_2502;
assign x_33793 = x_33791 & x_33792;
assign x_33794 = x_2503 & x_2504;
assign x_33795 = x_2505 & x_2506;
assign x_33796 = x_33794 & x_33795;
assign x_33797 = x_33793 & x_33796;
assign x_33798 = x_33790 & x_33797;
assign x_33799 = x_33783 & x_33798;
assign x_33800 = x_33769 & x_33799;
assign x_33801 = x_2508 & x_2509;
assign x_33802 = x_2507 & x_33801;
assign x_33803 = x_2510 & x_2511;
assign x_33804 = x_2512 & x_2513;
assign x_33805 = x_33803 & x_33804;
assign x_33806 = x_33802 & x_33805;
assign x_33807 = x_2514 & x_2515;
assign x_33808 = x_2516 & x_2517;
assign x_33809 = x_33807 & x_33808;
assign x_33810 = x_2518 & x_2519;
assign x_33811 = x_2520 & x_2521;
assign x_33812 = x_33810 & x_33811;
assign x_33813 = x_33809 & x_33812;
assign x_33814 = x_33806 & x_33813;
assign x_33815 = x_2523 & x_2524;
assign x_33816 = x_2522 & x_33815;
assign x_33817 = x_2525 & x_2526;
assign x_33818 = x_2527 & x_2528;
assign x_33819 = x_33817 & x_33818;
assign x_33820 = x_33816 & x_33819;
assign x_33821 = x_2529 & x_2530;
assign x_33822 = x_2531 & x_2532;
assign x_33823 = x_33821 & x_33822;
assign x_33824 = x_2533 & x_2534;
assign x_33825 = x_2535 & x_2536;
assign x_33826 = x_33824 & x_33825;
assign x_33827 = x_33823 & x_33826;
assign x_33828 = x_33820 & x_33827;
assign x_33829 = x_33814 & x_33828;
assign x_33830 = x_2538 & x_2539;
assign x_33831 = x_2537 & x_33830;
assign x_33832 = x_2540 & x_2541;
assign x_33833 = x_2542 & x_2543;
assign x_33834 = x_33832 & x_33833;
assign x_33835 = x_33831 & x_33834;
assign x_33836 = x_2544 & x_2545;
assign x_33837 = x_2546 & x_2547;
assign x_33838 = x_33836 & x_33837;
assign x_33839 = x_2548 & x_2549;
assign x_33840 = x_2550 & x_2551;
assign x_33841 = x_33839 & x_33840;
assign x_33842 = x_33838 & x_33841;
assign x_33843 = x_33835 & x_33842;
assign x_33844 = x_2552 & x_2553;
assign x_33845 = x_2554 & x_2555;
assign x_33846 = x_33844 & x_33845;
assign x_33847 = x_2556 & x_2557;
assign x_33848 = x_2558 & x_2559;
assign x_33849 = x_33847 & x_33848;
assign x_33850 = x_33846 & x_33849;
assign x_33851 = x_2560 & x_2561;
assign x_33852 = x_2562 & x_2563;
assign x_33853 = x_33851 & x_33852;
assign x_33854 = x_2564 & x_2565;
assign x_33855 = x_2566 & x_2567;
assign x_33856 = x_33854 & x_33855;
assign x_33857 = x_33853 & x_33856;
assign x_33858 = x_33850 & x_33857;
assign x_33859 = x_33843 & x_33858;
assign x_33860 = x_33829 & x_33859;
assign x_33861 = x_33800 & x_33860;
assign x_33862 = x_2569 & x_2570;
assign x_33863 = x_2568 & x_33862;
assign x_33864 = x_2571 & x_2572;
assign x_33865 = x_2573 & x_2574;
assign x_33866 = x_33864 & x_33865;
assign x_33867 = x_33863 & x_33866;
assign x_33868 = x_2575 & x_2576;
assign x_33869 = x_2577 & x_2578;
assign x_33870 = x_33868 & x_33869;
assign x_33871 = x_2579 & x_2580;
assign x_33872 = x_2581 & x_2582;
assign x_33873 = x_33871 & x_33872;
assign x_33874 = x_33870 & x_33873;
assign x_33875 = x_33867 & x_33874;
assign x_33876 = x_2584 & x_2585;
assign x_33877 = x_2583 & x_33876;
assign x_33878 = x_2586 & x_2587;
assign x_33879 = x_2588 & x_2589;
assign x_33880 = x_33878 & x_33879;
assign x_33881 = x_33877 & x_33880;
assign x_33882 = x_2590 & x_2591;
assign x_33883 = x_2592 & x_2593;
assign x_33884 = x_33882 & x_33883;
assign x_33885 = x_2594 & x_2595;
assign x_33886 = x_2596 & x_2597;
assign x_33887 = x_33885 & x_33886;
assign x_33888 = x_33884 & x_33887;
assign x_33889 = x_33881 & x_33888;
assign x_33890 = x_33875 & x_33889;
assign x_33891 = x_2599 & x_2600;
assign x_33892 = x_2598 & x_33891;
assign x_33893 = x_2601 & x_2602;
assign x_33894 = x_2603 & x_2604;
assign x_33895 = x_33893 & x_33894;
assign x_33896 = x_33892 & x_33895;
assign x_33897 = x_2605 & x_2606;
assign x_33898 = x_2607 & x_2608;
assign x_33899 = x_33897 & x_33898;
assign x_33900 = x_2609 & x_2610;
assign x_33901 = x_2611 & x_2612;
assign x_33902 = x_33900 & x_33901;
assign x_33903 = x_33899 & x_33902;
assign x_33904 = x_33896 & x_33903;
assign x_33905 = x_2613 & x_2614;
assign x_33906 = x_2615 & x_2616;
assign x_33907 = x_33905 & x_33906;
assign x_33908 = x_2617 & x_2618;
assign x_33909 = x_2619 & x_2620;
assign x_33910 = x_33908 & x_33909;
assign x_33911 = x_33907 & x_33910;
assign x_33912 = x_2621 & x_2622;
assign x_33913 = x_2623 & x_2624;
assign x_33914 = x_33912 & x_33913;
assign x_33915 = x_2625 & x_2626;
assign x_33916 = x_2627 & x_2628;
assign x_33917 = x_33915 & x_33916;
assign x_33918 = x_33914 & x_33917;
assign x_33919 = x_33911 & x_33918;
assign x_33920 = x_33904 & x_33919;
assign x_33921 = x_33890 & x_33920;
assign x_33922 = x_2630 & x_2631;
assign x_33923 = x_2629 & x_33922;
assign x_33924 = x_2632 & x_2633;
assign x_33925 = x_2634 & x_2635;
assign x_33926 = x_33924 & x_33925;
assign x_33927 = x_33923 & x_33926;
assign x_33928 = x_2636 & x_2637;
assign x_33929 = x_2638 & x_2639;
assign x_33930 = x_33928 & x_33929;
assign x_33931 = x_2640 & x_2641;
assign x_33932 = x_2642 & x_2643;
assign x_33933 = x_33931 & x_33932;
assign x_33934 = x_33930 & x_33933;
assign x_33935 = x_33927 & x_33934;
assign x_33936 = x_2645 & x_2646;
assign x_33937 = x_2644 & x_33936;
assign x_33938 = x_2647 & x_2648;
assign x_33939 = x_2649 & x_2650;
assign x_33940 = x_33938 & x_33939;
assign x_33941 = x_33937 & x_33940;
assign x_33942 = x_2651 & x_2652;
assign x_33943 = x_2653 & x_2654;
assign x_33944 = x_33942 & x_33943;
assign x_33945 = x_2655 & x_2656;
assign x_33946 = x_2657 & x_2658;
assign x_33947 = x_33945 & x_33946;
assign x_33948 = x_33944 & x_33947;
assign x_33949 = x_33941 & x_33948;
assign x_33950 = x_33935 & x_33949;
assign x_33951 = x_2660 & x_2661;
assign x_33952 = x_2659 & x_33951;
assign x_33953 = x_2662 & x_2663;
assign x_33954 = x_2664 & x_2665;
assign x_33955 = x_33953 & x_33954;
assign x_33956 = x_33952 & x_33955;
assign x_33957 = x_2666 & x_2667;
assign x_33958 = x_2668 & x_2669;
assign x_33959 = x_33957 & x_33958;
assign x_33960 = x_2670 & x_2671;
assign x_33961 = x_2672 & x_2673;
assign x_33962 = x_33960 & x_33961;
assign x_33963 = x_33959 & x_33962;
assign x_33964 = x_33956 & x_33963;
assign x_33965 = x_2674 & x_2675;
assign x_33966 = x_2676 & x_2677;
assign x_33967 = x_33965 & x_33966;
assign x_33968 = x_2678 & x_2679;
assign x_33969 = x_2680 & x_2681;
assign x_33970 = x_33968 & x_33969;
assign x_33971 = x_33967 & x_33970;
assign x_33972 = x_2682 & x_2683;
assign x_33973 = x_2684 & x_2685;
assign x_33974 = x_33972 & x_33973;
assign x_33975 = x_2686 & x_2687;
assign x_33976 = x_2688 & x_2689;
assign x_33977 = x_33975 & x_33976;
assign x_33978 = x_33974 & x_33977;
assign x_33979 = x_33971 & x_33978;
assign x_33980 = x_33964 & x_33979;
assign x_33981 = x_33950 & x_33980;
assign x_33982 = x_33921 & x_33981;
assign x_33983 = x_33861 & x_33982;
assign x_33984 = x_2691 & x_2692;
assign x_33985 = x_2690 & x_33984;
assign x_33986 = x_2693 & x_2694;
assign x_33987 = x_2695 & x_2696;
assign x_33988 = x_33986 & x_33987;
assign x_33989 = x_33985 & x_33988;
assign x_33990 = x_2697 & x_2698;
assign x_33991 = x_2699 & x_2700;
assign x_33992 = x_33990 & x_33991;
assign x_33993 = x_2701 & x_2702;
assign x_33994 = x_2703 & x_2704;
assign x_33995 = x_33993 & x_33994;
assign x_33996 = x_33992 & x_33995;
assign x_33997 = x_33989 & x_33996;
assign x_33998 = x_2706 & x_2707;
assign x_33999 = x_2705 & x_33998;
assign x_34000 = x_2708 & x_2709;
assign x_34001 = x_2710 & x_2711;
assign x_34002 = x_34000 & x_34001;
assign x_34003 = x_33999 & x_34002;
assign x_34004 = x_2712 & x_2713;
assign x_34005 = x_2714 & x_2715;
assign x_34006 = x_34004 & x_34005;
assign x_34007 = x_2716 & x_2717;
assign x_34008 = x_2718 & x_2719;
assign x_34009 = x_34007 & x_34008;
assign x_34010 = x_34006 & x_34009;
assign x_34011 = x_34003 & x_34010;
assign x_34012 = x_33997 & x_34011;
assign x_34013 = x_2721 & x_2722;
assign x_34014 = x_2720 & x_34013;
assign x_34015 = x_2723 & x_2724;
assign x_34016 = x_2725 & x_2726;
assign x_34017 = x_34015 & x_34016;
assign x_34018 = x_34014 & x_34017;
assign x_34019 = x_2727 & x_2728;
assign x_34020 = x_2729 & x_2730;
assign x_34021 = x_34019 & x_34020;
assign x_34022 = x_2731 & x_2732;
assign x_34023 = x_2733 & x_2734;
assign x_34024 = x_34022 & x_34023;
assign x_34025 = x_34021 & x_34024;
assign x_34026 = x_34018 & x_34025;
assign x_34027 = x_2735 & x_2736;
assign x_34028 = x_2737 & x_2738;
assign x_34029 = x_34027 & x_34028;
assign x_34030 = x_2739 & x_2740;
assign x_34031 = x_2741 & x_2742;
assign x_34032 = x_34030 & x_34031;
assign x_34033 = x_34029 & x_34032;
assign x_34034 = x_2743 & x_2744;
assign x_34035 = x_2745 & x_2746;
assign x_34036 = x_34034 & x_34035;
assign x_34037 = x_2747 & x_2748;
assign x_34038 = x_2749 & x_2750;
assign x_34039 = x_34037 & x_34038;
assign x_34040 = x_34036 & x_34039;
assign x_34041 = x_34033 & x_34040;
assign x_34042 = x_34026 & x_34041;
assign x_34043 = x_34012 & x_34042;
assign x_34044 = x_2752 & x_2753;
assign x_34045 = x_2751 & x_34044;
assign x_34046 = x_2754 & x_2755;
assign x_34047 = x_2756 & x_2757;
assign x_34048 = x_34046 & x_34047;
assign x_34049 = x_34045 & x_34048;
assign x_34050 = x_2758 & x_2759;
assign x_34051 = x_2760 & x_2761;
assign x_34052 = x_34050 & x_34051;
assign x_34053 = x_2762 & x_2763;
assign x_34054 = x_2764 & x_2765;
assign x_34055 = x_34053 & x_34054;
assign x_34056 = x_34052 & x_34055;
assign x_34057 = x_34049 & x_34056;
assign x_34058 = x_2767 & x_2768;
assign x_34059 = x_2766 & x_34058;
assign x_34060 = x_2769 & x_2770;
assign x_34061 = x_2771 & x_2772;
assign x_34062 = x_34060 & x_34061;
assign x_34063 = x_34059 & x_34062;
assign x_34064 = x_2773 & x_2774;
assign x_34065 = x_2775 & x_2776;
assign x_34066 = x_34064 & x_34065;
assign x_34067 = x_2777 & x_2778;
assign x_34068 = x_2779 & x_2780;
assign x_34069 = x_34067 & x_34068;
assign x_34070 = x_34066 & x_34069;
assign x_34071 = x_34063 & x_34070;
assign x_34072 = x_34057 & x_34071;
assign x_34073 = x_2782 & x_2783;
assign x_34074 = x_2781 & x_34073;
assign x_34075 = x_2784 & x_2785;
assign x_34076 = x_2786 & x_2787;
assign x_34077 = x_34075 & x_34076;
assign x_34078 = x_34074 & x_34077;
assign x_34079 = x_2788 & x_2789;
assign x_34080 = x_2790 & x_2791;
assign x_34081 = x_34079 & x_34080;
assign x_34082 = x_2792 & x_2793;
assign x_34083 = x_2794 & x_2795;
assign x_34084 = x_34082 & x_34083;
assign x_34085 = x_34081 & x_34084;
assign x_34086 = x_34078 & x_34085;
assign x_34087 = x_2796 & x_2797;
assign x_34088 = x_2798 & x_2799;
assign x_34089 = x_34087 & x_34088;
assign x_34090 = x_2800 & x_2801;
assign x_34091 = x_2802 & x_2803;
assign x_34092 = x_34090 & x_34091;
assign x_34093 = x_34089 & x_34092;
assign x_34094 = x_2804 & x_2805;
assign x_34095 = x_2806 & x_2807;
assign x_34096 = x_34094 & x_34095;
assign x_34097 = x_2808 & x_2809;
assign x_34098 = x_2810 & x_2811;
assign x_34099 = x_34097 & x_34098;
assign x_34100 = x_34096 & x_34099;
assign x_34101 = x_34093 & x_34100;
assign x_34102 = x_34086 & x_34101;
assign x_34103 = x_34072 & x_34102;
assign x_34104 = x_34043 & x_34103;
assign x_34105 = x_2813 & x_2814;
assign x_34106 = x_2812 & x_34105;
assign x_34107 = x_2815 & x_2816;
assign x_34108 = x_2817 & x_2818;
assign x_34109 = x_34107 & x_34108;
assign x_34110 = x_34106 & x_34109;
assign x_34111 = x_2819 & x_2820;
assign x_34112 = x_2821 & x_2822;
assign x_34113 = x_34111 & x_34112;
assign x_34114 = x_2823 & x_2824;
assign x_34115 = x_2825 & x_2826;
assign x_34116 = x_34114 & x_34115;
assign x_34117 = x_34113 & x_34116;
assign x_34118 = x_34110 & x_34117;
assign x_34119 = x_2828 & x_2829;
assign x_34120 = x_2827 & x_34119;
assign x_34121 = x_2830 & x_2831;
assign x_34122 = x_2832 & x_2833;
assign x_34123 = x_34121 & x_34122;
assign x_34124 = x_34120 & x_34123;
assign x_34125 = x_2834 & x_2835;
assign x_34126 = x_2836 & x_2837;
assign x_34127 = x_34125 & x_34126;
assign x_34128 = x_2838 & x_2839;
assign x_34129 = x_2840 & x_2841;
assign x_34130 = x_34128 & x_34129;
assign x_34131 = x_34127 & x_34130;
assign x_34132 = x_34124 & x_34131;
assign x_34133 = x_34118 & x_34132;
assign x_34134 = x_2843 & x_2844;
assign x_34135 = x_2842 & x_34134;
assign x_34136 = x_2845 & x_2846;
assign x_34137 = x_2847 & x_2848;
assign x_34138 = x_34136 & x_34137;
assign x_34139 = x_34135 & x_34138;
assign x_34140 = x_2849 & x_2850;
assign x_34141 = x_2851 & x_2852;
assign x_34142 = x_34140 & x_34141;
assign x_34143 = x_2853 & x_2854;
assign x_34144 = x_2855 & x_2856;
assign x_34145 = x_34143 & x_34144;
assign x_34146 = x_34142 & x_34145;
assign x_34147 = x_34139 & x_34146;
assign x_34148 = x_2857 & x_2858;
assign x_34149 = x_2859 & x_2860;
assign x_34150 = x_34148 & x_34149;
assign x_34151 = x_2861 & x_2862;
assign x_34152 = x_2863 & x_2864;
assign x_34153 = x_34151 & x_34152;
assign x_34154 = x_34150 & x_34153;
assign x_34155 = x_2865 & x_2866;
assign x_34156 = x_2867 & x_2868;
assign x_34157 = x_34155 & x_34156;
assign x_34158 = x_2869 & x_2870;
assign x_34159 = x_2871 & x_2872;
assign x_34160 = x_34158 & x_34159;
assign x_34161 = x_34157 & x_34160;
assign x_34162 = x_34154 & x_34161;
assign x_34163 = x_34147 & x_34162;
assign x_34164 = x_34133 & x_34163;
assign x_34165 = x_2874 & x_2875;
assign x_34166 = x_2873 & x_34165;
assign x_34167 = x_2876 & x_2877;
assign x_34168 = x_2878 & x_2879;
assign x_34169 = x_34167 & x_34168;
assign x_34170 = x_34166 & x_34169;
assign x_34171 = x_2880 & x_2881;
assign x_34172 = x_2882 & x_2883;
assign x_34173 = x_34171 & x_34172;
assign x_34174 = x_2884 & x_2885;
assign x_34175 = x_2886 & x_2887;
assign x_34176 = x_34174 & x_34175;
assign x_34177 = x_34173 & x_34176;
assign x_34178 = x_34170 & x_34177;
assign x_34179 = x_2888 & x_2889;
assign x_34180 = x_2890 & x_2891;
assign x_34181 = x_34179 & x_34180;
assign x_34182 = x_2892 & x_2893;
assign x_34183 = x_2894 & x_2895;
assign x_34184 = x_34182 & x_34183;
assign x_34185 = x_34181 & x_34184;
assign x_34186 = x_2896 & x_2897;
assign x_34187 = x_2898 & x_2899;
assign x_34188 = x_34186 & x_34187;
assign x_34189 = x_2900 & x_2901;
assign x_34190 = x_2902 & x_2903;
assign x_34191 = x_34189 & x_34190;
assign x_34192 = x_34188 & x_34191;
assign x_34193 = x_34185 & x_34192;
assign x_34194 = x_34178 & x_34193;
assign x_34195 = x_2905 & x_2906;
assign x_34196 = x_2904 & x_34195;
assign x_34197 = x_2907 & x_2908;
assign x_34198 = x_2909 & x_2910;
assign x_34199 = x_34197 & x_34198;
assign x_34200 = x_34196 & x_34199;
assign x_34201 = x_2911 & x_2912;
assign x_34202 = x_2913 & x_2914;
assign x_34203 = x_34201 & x_34202;
assign x_34204 = x_2915 & x_2916;
assign x_34205 = x_2917 & x_2918;
assign x_34206 = x_34204 & x_34205;
assign x_34207 = x_34203 & x_34206;
assign x_34208 = x_34200 & x_34207;
assign x_34209 = x_2919 & x_2920;
assign x_34210 = x_2921 & x_2922;
assign x_34211 = x_34209 & x_34210;
assign x_34212 = x_2923 & x_2924;
assign x_34213 = x_2925 & x_2926;
assign x_34214 = x_34212 & x_34213;
assign x_34215 = x_34211 & x_34214;
assign x_34216 = x_2927 & x_2928;
assign x_34217 = x_2929 & x_2930;
assign x_34218 = x_34216 & x_34217;
assign x_34219 = x_2931 & x_2932;
assign x_34220 = x_2933 & x_2934;
assign x_34221 = x_34219 & x_34220;
assign x_34222 = x_34218 & x_34221;
assign x_34223 = x_34215 & x_34222;
assign x_34224 = x_34208 & x_34223;
assign x_34225 = x_34194 & x_34224;
assign x_34226 = x_34164 & x_34225;
assign x_34227 = x_34104 & x_34226;
assign x_34228 = x_33983 & x_34227;
assign x_34229 = x_33740 & x_34228;
assign x_34230 = x_2936 & x_2937;
assign x_34231 = x_2935 & x_34230;
assign x_34232 = x_2938 & x_2939;
assign x_34233 = x_2940 & x_2941;
assign x_34234 = x_34232 & x_34233;
assign x_34235 = x_34231 & x_34234;
assign x_34236 = x_2942 & x_2943;
assign x_34237 = x_2944 & x_2945;
assign x_34238 = x_34236 & x_34237;
assign x_34239 = x_2946 & x_2947;
assign x_34240 = x_2948 & x_2949;
assign x_34241 = x_34239 & x_34240;
assign x_34242 = x_34238 & x_34241;
assign x_34243 = x_34235 & x_34242;
assign x_34244 = x_2951 & x_2952;
assign x_34245 = x_2950 & x_34244;
assign x_34246 = x_2953 & x_2954;
assign x_34247 = x_2955 & x_2956;
assign x_34248 = x_34246 & x_34247;
assign x_34249 = x_34245 & x_34248;
assign x_34250 = x_2957 & x_2958;
assign x_34251 = x_2959 & x_2960;
assign x_34252 = x_34250 & x_34251;
assign x_34253 = x_2961 & x_2962;
assign x_34254 = x_2963 & x_2964;
assign x_34255 = x_34253 & x_34254;
assign x_34256 = x_34252 & x_34255;
assign x_34257 = x_34249 & x_34256;
assign x_34258 = x_34243 & x_34257;
assign x_34259 = x_2966 & x_2967;
assign x_34260 = x_2965 & x_34259;
assign x_34261 = x_2968 & x_2969;
assign x_34262 = x_2970 & x_2971;
assign x_34263 = x_34261 & x_34262;
assign x_34264 = x_34260 & x_34263;
assign x_34265 = x_2972 & x_2973;
assign x_34266 = x_2974 & x_2975;
assign x_34267 = x_34265 & x_34266;
assign x_34268 = x_2976 & x_2977;
assign x_34269 = x_2978 & x_2979;
assign x_34270 = x_34268 & x_34269;
assign x_34271 = x_34267 & x_34270;
assign x_34272 = x_34264 & x_34271;
assign x_34273 = x_2980 & x_2981;
assign x_34274 = x_2982 & x_2983;
assign x_34275 = x_34273 & x_34274;
assign x_34276 = x_2984 & x_2985;
assign x_34277 = x_2986 & x_2987;
assign x_34278 = x_34276 & x_34277;
assign x_34279 = x_34275 & x_34278;
assign x_34280 = x_2988 & x_2989;
assign x_34281 = x_2990 & x_2991;
assign x_34282 = x_34280 & x_34281;
assign x_34283 = x_2992 & x_2993;
assign x_34284 = x_2994 & x_2995;
assign x_34285 = x_34283 & x_34284;
assign x_34286 = x_34282 & x_34285;
assign x_34287 = x_34279 & x_34286;
assign x_34288 = x_34272 & x_34287;
assign x_34289 = x_34258 & x_34288;
assign x_34290 = x_2997 & x_2998;
assign x_34291 = x_2996 & x_34290;
assign x_34292 = x_2999 & x_3000;
assign x_34293 = x_3001 & x_3002;
assign x_34294 = x_34292 & x_34293;
assign x_34295 = x_34291 & x_34294;
assign x_34296 = x_3003 & x_3004;
assign x_34297 = x_3005 & x_3006;
assign x_34298 = x_34296 & x_34297;
assign x_34299 = x_3007 & x_3008;
assign x_34300 = x_3009 & x_3010;
assign x_34301 = x_34299 & x_34300;
assign x_34302 = x_34298 & x_34301;
assign x_34303 = x_34295 & x_34302;
assign x_34304 = x_3012 & x_3013;
assign x_34305 = x_3011 & x_34304;
assign x_34306 = x_3014 & x_3015;
assign x_34307 = x_3016 & x_3017;
assign x_34308 = x_34306 & x_34307;
assign x_34309 = x_34305 & x_34308;
assign x_34310 = x_3018 & x_3019;
assign x_34311 = x_3020 & x_3021;
assign x_34312 = x_34310 & x_34311;
assign x_34313 = x_3022 & x_3023;
assign x_34314 = x_3024 & x_3025;
assign x_34315 = x_34313 & x_34314;
assign x_34316 = x_34312 & x_34315;
assign x_34317 = x_34309 & x_34316;
assign x_34318 = x_34303 & x_34317;
assign x_34319 = x_3027 & x_3028;
assign x_34320 = x_3026 & x_34319;
assign x_34321 = x_3029 & x_3030;
assign x_34322 = x_3031 & x_3032;
assign x_34323 = x_34321 & x_34322;
assign x_34324 = x_34320 & x_34323;
assign x_34325 = x_3033 & x_3034;
assign x_34326 = x_3035 & x_3036;
assign x_34327 = x_34325 & x_34326;
assign x_34328 = x_3037 & x_3038;
assign x_34329 = x_3039 & x_3040;
assign x_34330 = x_34328 & x_34329;
assign x_34331 = x_34327 & x_34330;
assign x_34332 = x_34324 & x_34331;
assign x_34333 = x_3041 & x_3042;
assign x_34334 = x_3043 & x_3044;
assign x_34335 = x_34333 & x_34334;
assign x_34336 = x_3045 & x_3046;
assign x_34337 = x_3047 & x_3048;
assign x_34338 = x_34336 & x_34337;
assign x_34339 = x_34335 & x_34338;
assign x_34340 = x_3049 & x_3050;
assign x_34341 = x_3051 & x_3052;
assign x_34342 = x_34340 & x_34341;
assign x_34343 = x_3053 & x_3054;
assign x_34344 = x_3055 & x_3056;
assign x_34345 = x_34343 & x_34344;
assign x_34346 = x_34342 & x_34345;
assign x_34347 = x_34339 & x_34346;
assign x_34348 = x_34332 & x_34347;
assign x_34349 = x_34318 & x_34348;
assign x_34350 = x_34289 & x_34349;
assign x_34351 = x_3058 & x_3059;
assign x_34352 = x_3057 & x_34351;
assign x_34353 = x_3060 & x_3061;
assign x_34354 = x_3062 & x_3063;
assign x_34355 = x_34353 & x_34354;
assign x_34356 = x_34352 & x_34355;
assign x_34357 = x_3064 & x_3065;
assign x_34358 = x_3066 & x_3067;
assign x_34359 = x_34357 & x_34358;
assign x_34360 = x_3068 & x_3069;
assign x_34361 = x_3070 & x_3071;
assign x_34362 = x_34360 & x_34361;
assign x_34363 = x_34359 & x_34362;
assign x_34364 = x_34356 & x_34363;
assign x_34365 = x_3073 & x_3074;
assign x_34366 = x_3072 & x_34365;
assign x_34367 = x_3075 & x_3076;
assign x_34368 = x_3077 & x_3078;
assign x_34369 = x_34367 & x_34368;
assign x_34370 = x_34366 & x_34369;
assign x_34371 = x_3079 & x_3080;
assign x_34372 = x_3081 & x_3082;
assign x_34373 = x_34371 & x_34372;
assign x_34374 = x_3083 & x_3084;
assign x_34375 = x_3085 & x_3086;
assign x_34376 = x_34374 & x_34375;
assign x_34377 = x_34373 & x_34376;
assign x_34378 = x_34370 & x_34377;
assign x_34379 = x_34364 & x_34378;
assign x_34380 = x_3088 & x_3089;
assign x_34381 = x_3087 & x_34380;
assign x_34382 = x_3090 & x_3091;
assign x_34383 = x_3092 & x_3093;
assign x_34384 = x_34382 & x_34383;
assign x_34385 = x_34381 & x_34384;
assign x_34386 = x_3094 & x_3095;
assign x_34387 = x_3096 & x_3097;
assign x_34388 = x_34386 & x_34387;
assign x_34389 = x_3098 & x_3099;
assign x_34390 = x_3100 & x_3101;
assign x_34391 = x_34389 & x_34390;
assign x_34392 = x_34388 & x_34391;
assign x_34393 = x_34385 & x_34392;
assign x_34394 = x_3102 & x_3103;
assign x_34395 = x_3104 & x_3105;
assign x_34396 = x_34394 & x_34395;
assign x_34397 = x_3106 & x_3107;
assign x_34398 = x_3108 & x_3109;
assign x_34399 = x_34397 & x_34398;
assign x_34400 = x_34396 & x_34399;
assign x_34401 = x_3110 & x_3111;
assign x_34402 = x_3112 & x_3113;
assign x_34403 = x_34401 & x_34402;
assign x_34404 = x_3114 & x_3115;
assign x_34405 = x_3116 & x_3117;
assign x_34406 = x_34404 & x_34405;
assign x_34407 = x_34403 & x_34406;
assign x_34408 = x_34400 & x_34407;
assign x_34409 = x_34393 & x_34408;
assign x_34410 = x_34379 & x_34409;
assign x_34411 = x_3119 & x_3120;
assign x_34412 = x_3118 & x_34411;
assign x_34413 = x_3121 & x_3122;
assign x_34414 = x_3123 & x_3124;
assign x_34415 = x_34413 & x_34414;
assign x_34416 = x_34412 & x_34415;
assign x_34417 = x_3125 & x_3126;
assign x_34418 = x_3127 & x_3128;
assign x_34419 = x_34417 & x_34418;
assign x_34420 = x_3129 & x_3130;
assign x_34421 = x_3131 & x_3132;
assign x_34422 = x_34420 & x_34421;
assign x_34423 = x_34419 & x_34422;
assign x_34424 = x_34416 & x_34423;
assign x_34425 = x_3134 & x_3135;
assign x_34426 = x_3133 & x_34425;
assign x_34427 = x_3136 & x_3137;
assign x_34428 = x_3138 & x_3139;
assign x_34429 = x_34427 & x_34428;
assign x_34430 = x_34426 & x_34429;
assign x_34431 = x_3140 & x_3141;
assign x_34432 = x_3142 & x_3143;
assign x_34433 = x_34431 & x_34432;
assign x_34434 = x_3144 & x_3145;
assign x_34435 = x_3146 & x_3147;
assign x_34436 = x_34434 & x_34435;
assign x_34437 = x_34433 & x_34436;
assign x_34438 = x_34430 & x_34437;
assign x_34439 = x_34424 & x_34438;
assign x_34440 = x_3149 & x_3150;
assign x_34441 = x_3148 & x_34440;
assign x_34442 = x_3151 & x_3152;
assign x_34443 = x_3153 & x_3154;
assign x_34444 = x_34442 & x_34443;
assign x_34445 = x_34441 & x_34444;
assign x_34446 = x_3155 & x_3156;
assign x_34447 = x_3157 & x_3158;
assign x_34448 = x_34446 & x_34447;
assign x_34449 = x_3159 & x_3160;
assign x_34450 = x_3161 & x_3162;
assign x_34451 = x_34449 & x_34450;
assign x_34452 = x_34448 & x_34451;
assign x_34453 = x_34445 & x_34452;
assign x_34454 = x_3163 & x_3164;
assign x_34455 = x_3165 & x_3166;
assign x_34456 = x_34454 & x_34455;
assign x_34457 = x_3167 & x_3168;
assign x_34458 = x_3169 & x_3170;
assign x_34459 = x_34457 & x_34458;
assign x_34460 = x_34456 & x_34459;
assign x_34461 = x_3171 & x_3172;
assign x_34462 = x_3173 & x_3174;
assign x_34463 = x_34461 & x_34462;
assign x_34464 = x_3175 & x_3176;
assign x_34465 = x_3177 & x_3178;
assign x_34466 = x_34464 & x_34465;
assign x_34467 = x_34463 & x_34466;
assign x_34468 = x_34460 & x_34467;
assign x_34469 = x_34453 & x_34468;
assign x_34470 = x_34439 & x_34469;
assign x_34471 = x_34410 & x_34470;
assign x_34472 = x_34350 & x_34471;
assign x_34473 = x_3180 & x_3181;
assign x_34474 = x_3179 & x_34473;
assign x_34475 = x_3182 & x_3183;
assign x_34476 = x_3184 & x_3185;
assign x_34477 = x_34475 & x_34476;
assign x_34478 = x_34474 & x_34477;
assign x_34479 = x_3186 & x_3187;
assign x_34480 = x_3188 & x_3189;
assign x_34481 = x_34479 & x_34480;
assign x_34482 = x_3190 & x_3191;
assign x_34483 = x_3192 & x_3193;
assign x_34484 = x_34482 & x_34483;
assign x_34485 = x_34481 & x_34484;
assign x_34486 = x_34478 & x_34485;
assign x_34487 = x_3195 & x_3196;
assign x_34488 = x_3194 & x_34487;
assign x_34489 = x_3197 & x_3198;
assign x_34490 = x_3199 & x_3200;
assign x_34491 = x_34489 & x_34490;
assign x_34492 = x_34488 & x_34491;
assign x_34493 = x_3201 & x_3202;
assign x_34494 = x_3203 & x_3204;
assign x_34495 = x_34493 & x_34494;
assign x_34496 = x_3205 & x_3206;
assign x_34497 = x_3207 & x_3208;
assign x_34498 = x_34496 & x_34497;
assign x_34499 = x_34495 & x_34498;
assign x_34500 = x_34492 & x_34499;
assign x_34501 = x_34486 & x_34500;
assign x_34502 = x_3210 & x_3211;
assign x_34503 = x_3209 & x_34502;
assign x_34504 = x_3212 & x_3213;
assign x_34505 = x_3214 & x_3215;
assign x_34506 = x_34504 & x_34505;
assign x_34507 = x_34503 & x_34506;
assign x_34508 = x_3216 & x_3217;
assign x_34509 = x_3218 & x_3219;
assign x_34510 = x_34508 & x_34509;
assign x_34511 = x_3220 & x_3221;
assign x_34512 = x_3222 & x_3223;
assign x_34513 = x_34511 & x_34512;
assign x_34514 = x_34510 & x_34513;
assign x_34515 = x_34507 & x_34514;
assign x_34516 = x_3224 & x_3225;
assign x_34517 = x_3226 & x_3227;
assign x_34518 = x_34516 & x_34517;
assign x_34519 = x_3228 & x_3229;
assign x_34520 = x_3230 & x_3231;
assign x_34521 = x_34519 & x_34520;
assign x_34522 = x_34518 & x_34521;
assign x_34523 = x_3232 & x_3233;
assign x_34524 = x_3234 & x_3235;
assign x_34525 = x_34523 & x_34524;
assign x_34526 = x_3236 & x_3237;
assign x_34527 = x_3238 & x_3239;
assign x_34528 = x_34526 & x_34527;
assign x_34529 = x_34525 & x_34528;
assign x_34530 = x_34522 & x_34529;
assign x_34531 = x_34515 & x_34530;
assign x_34532 = x_34501 & x_34531;
assign x_34533 = x_3241 & x_3242;
assign x_34534 = x_3240 & x_34533;
assign x_34535 = x_3243 & x_3244;
assign x_34536 = x_3245 & x_3246;
assign x_34537 = x_34535 & x_34536;
assign x_34538 = x_34534 & x_34537;
assign x_34539 = x_3247 & x_3248;
assign x_34540 = x_3249 & x_3250;
assign x_34541 = x_34539 & x_34540;
assign x_34542 = x_3251 & x_3252;
assign x_34543 = x_3253 & x_3254;
assign x_34544 = x_34542 & x_34543;
assign x_34545 = x_34541 & x_34544;
assign x_34546 = x_34538 & x_34545;
assign x_34547 = x_3256 & x_3257;
assign x_34548 = x_3255 & x_34547;
assign x_34549 = x_3258 & x_3259;
assign x_34550 = x_3260 & x_3261;
assign x_34551 = x_34549 & x_34550;
assign x_34552 = x_34548 & x_34551;
assign x_34553 = x_3262 & x_3263;
assign x_34554 = x_3264 & x_3265;
assign x_34555 = x_34553 & x_34554;
assign x_34556 = x_3266 & x_3267;
assign x_34557 = x_3268 & x_3269;
assign x_34558 = x_34556 & x_34557;
assign x_34559 = x_34555 & x_34558;
assign x_34560 = x_34552 & x_34559;
assign x_34561 = x_34546 & x_34560;
assign x_34562 = x_3271 & x_3272;
assign x_34563 = x_3270 & x_34562;
assign x_34564 = x_3273 & x_3274;
assign x_34565 = x_3275 & x_3276;
assign x_34566 = x_34564 & x_34565;
assign x_34567 = x_34563 & x_34566;
assign x_34568 = x_3277 & x_3278;
assign x_34569 = x_3279 & x_3280;
assign x_34570 = x_34568 & x_34569;
assign x_34571 = x_3281 & x_3282;
assign x_34572 = x_3283 & x_3284;
assign x_34573 = x_34571 & x_34572;
assign x_34574 = x_34570 & x_34573;
assign x_34575 = x_34567 & x_34574;
assign x_34576 = x_3285 & x_3286;
assign x_34577 = x_3287 & x_3288;
assign x_34578 = x_34576 & x_34577;
assign x_34579 = x_3289 & x_3290;
assign x_34580 = x_3291 & x_3292;
assign x_34581 = x_34579 & x_34580;
assign x_34582 = x_34578 & x_34581;
assign x_34583 = x_3293 & x_3294;
assign x_34584 = x_3295 & x_3296;
assign x_34585 = x_34583 & x_34584;
assign x_34586 = x_3297 & x_3298;
assign x_34587 = x_3299 & x_3300;
assign x_34588 = x_34586 & x_34587;
assign x_34589 = x_34585 & x_34588;
assign x_34590 = x_34582 & x_34589;
assign x_34591 = x_34575 & x_34590;
assign x_34592 = x_34561 & x_34591;
assign x_34593 = x_34532 & x_34592;
assign x_34594 = x_3302 & x_3303;
assign x_34595 = x_3301 & x_34594;
assign x_34596 = x_3304 & x_3305;
assign x_34597 = x_3306 & x_3307;
assign x_34598 = x_34596 & x_34597;
assign x_34599 = x_34595 & x_34598;
assign x_34600 = x_3308 & x_3309;
assign x_34601 = x_3310 & x_3311;
assign x_34602 = x_34600 & x_34601;
assign x_34603 = x_3312 & x_3313;
assign x_34604 = x_3314 & x_3315;
assign x_34605 = x_34603 & x_34604;
assign x_34606 = x_34602 & x_34605;
assign x_34607 = x_34599 & x_34606;
assign x_34608 = x_3317 & x_3318;
assign x_34609 = x_3316 & x_34608;
assign x_34610 = x_3319 & x_3320;
assign x_34611 = x_3321 & x_3322;
assign x_34612 = x_34610 & x_34611;
assign x_34613 = x_34609 & x_34612;
assign x_34614 = x_3323 & x_3324;
assign x_34615 = x_3325 & x_3326;
assign x_34616 = x_34614 & x_34615;
assign x_34617 = x_3327 & x_3328;
assign x_34618 = x_3329 & x_3330;
assign x_34619 = x_34617 & x_34618;
assign x_34620 = x_34616 & x_34619;
assign x_34621 = x_34613 & x_34620;
assign x_34622 = x_34607 & x_34621;
assign x_34623 = x_3332 & x_3333;
assign x_34624 = x_3331 & x_34623;
assign x_34625 = x_3334 & x_3335;
assign x_34626 = x_3336 & x_3337;
assign x_34627 = x_34625 & x_34626;
assign x_34628 = x_34624 & x_34627;
assign x_34629 = x_3338 & x_3339;
assign x_34630 = x_3340 & x_3341;
assign x_34631 = x_34629 & x_34630;
assign x_34632 = x_3342 & x_3343;
assign x_34633 = x_3344 & x_3345;
assign x_34634 = x_34632 & x_34633;
assign x_34635 = x_34631 & x_34634;
assign x_34636 = x_34628 & x_34635;
assign x_34637 = x_3346 & x_3347;
assign x_34638 = x_3348 & x_3349;
assign x_34639 = x_34637 & x_34638;
assign x_34640 = x_3350 & x_3351;
assign x_34641 = x_3352 & x_3353;
assign x_34642 = x_34640 & x_34641;
assign x_34643 = x_34639 & x_34642;
assign x_34644 = x_3354 & x_3355;
assign x_34645 = x_3356 & x_3357;
assign x_34646 = x_34644 & x_34645;
assign x_34647 = x_3358 & x_3359;
assign x_34648 = x_3360 & x_3361;
assign x_34649 = x_34647 & x_34648;
assign x_34650 = x_34646 & x_34649;
assign x_34651 = x_34643 & x_34650;
assign x_34652 = x_34636 & x_34651;
assign x_34653 = x_34622 & x_34652;
assign x_34654 = x_3363 & x_3364;
assign x_34655 = x_3362 & x_34654;
assign x_34656 = x_3365 & x_3366;
assign x_34657 = x_3367 & x_3368;
assign x_34658 = x_34656 & x_34657;
assign x_34659 = x_34655 & x_34658;
assign x_34660 = x_3369 & x_3370;
assign x_34661 = x_3371 & x_3372;
assign x_34662 = x_34660 & x_34661;
assign x_34663 = x_3373 & x_3374;
assign x_34664 = x_3375 & x_3376;
assign x_34665 = x_34663 & x_34664;
assign x_34666 = x_34662 & x_34665;
assign x_34667 = x_34659 & x_34666;
assign x_34668 = x_3377 & x_3378;
assign x_34669 = x_3379 & x_3380;
assign x_34670 = x_34668 & x_34669;
assign x_34671 = x_3381 & x_3382;
assign x_34672 = x_3383 & x_3384;
assign x_34673 = x_34671 & x_34672;
assign x_34674 = x_34670 & x_34673;
assign x_34675 = x_3385 & x_3386;
assign x_34676 = x_3387 & x_3388;
assign x_34677 = x_34675 & x_34676;
assign x_34678 = x_3389 & x_3390;
assign x_34679 = x_3391 & x_3392;
assign x_34680 = x_34678 & x_34679;
assign x_34681 = x_34677 & x_34680;
assign x_34682 = x_34674 & x_34681;
assign x_34683 = x_34667 & x_34682;
assign x_34684 = x_3394 & x_3395;
assign x_34685 = x_3393 & x_34684;
assign x_34686 = x_3396 & x_3397;
assign x_34687 = x_3398 & x_3399;
assign x_34688 = x_34686 & x_34687;
assign x_34689 = x_34685 & x_34688;
assign x_34690 = x_3400 & x_3401;
assign x_34691 = x_3402 & x_3403;
assign x_34692 = x_34690 & x_34691;
assign x_34693 = x_3404 & x_3405;
assign x_34694 = x_3406 & x_3407;
assign x_34695 = x_34693 & x_34694;
assign x_34696 = x_34692 & x_34695;
assign x_34697 = x_34689 & x_34696;
assign x_34698 = x_3408 & x_3409;
assign x_34699 = x_3410 & x_3411;
assign x_34700 = x_34698 & x_34699;
assign x_34701 = x_3412 & x_3413;
assign x_34702 = x_3414 & x_3415;
assign x_34703 = x_34701 & x_34702;
assign x_34704 = x_34700 & x_34703;
assign x_34705 = x_3416 & x_3417;
assign x_34706 = x_3418 & x_3419;
assign x_34707 = x_34705 & x_34706;
assign x_34708 = x_3420 & x_3421;
assign x_34709 = x_3422 & x_3423;
assign x_34710 = x_34708 & x_34709;
assign x_34711 = x_34707 & x_34710;
assign x_34712 = x_34704 & x_34711;
assign x_34713 = x_34697 & x_34712;
assign x_34714 = x_34683 & x_34713;
assign x_34715 = x_34653 & x_34714;
assign x_34716 = x_34593 & x_34715;
assign x_34717 = x_34472 & x_34716;
assign x_34718 = x_3425 & x_3426;
assign x_34719 = x_3424 & x_34718;
assign x_34720 = x_3427 & x_3428;
assign x_34721 = x_3429 & x_3430;
assign x_34722 = x_34720 & x_34721;
assign x_34723 = x_34719 & x_34722;
assign x_34724 = x_3431 & x_3432;
assign x_34725 = x_3433 & x_3434;
assign x_34726 = x_34724 & x_34725;
assign x_34727 = x_3435 & x_3436;
assign x_34728 = x_3437 & x_3438;
assign x_34729 = x_34727 & x_34728;
assign x_34730 = x_34726 & x_34729;
assign x_34731 = x_34723 & x_34730;
assign x_34732 = x_3440 & x_3441;
assign x_34733 = x_3439 & x_34732;
assign x_34734 = x_3442 & x_3443;
assign x_34735 = x_3444 & x_3445;
assign x_34736 = x_34734 & x_34735;
assign x_34737 = x_34733 & x_34736;
assign x_34738 = x_3446 & x_3447;
assign x_34739 = x_3448 & x_3449;
assign x_34740 = x_34738 & x_34739;
assign x_34741 = x_3450 & x_3451;
assign x_34742 = x_3452 & x_3453;
assign x_34743 = x_34741 & x_34742;
assign x_34744 = x_34740 & x_34743;
assign x_34745 = x_34737 & x_34744;
assign x_34746 = x_34731 & x_34745;
assign x_34747 = x_3455 & x_3456;
assign x_34748 = x_3454 & x_34747;
assign x_34749 = x_3457 & x_3458;
assign x_34750 = x_3459 & x_3460;
assign x_34751 = x_34749 & x_34750;
assign x_34752 = x_34748 & x_34751;
assign x_34753 = x_3461 & x_3462;
assign x_34754 = x_3463 & x_3464;
assign x_34755 = x_34753 & x_34754;
assign x_34756 = x_3465 & x_3466;
assign x_34757 = x_3467 & x_3468;
assign x_34758 = x_34756 & x_34757;
assign x_34759 = x_34755 & x_34758;
assign x_34760 = x_34752 & x_34759;
assign x_34761 = x_3469 & x_3470;
assign x_34762 = x_3471 & x_3472;
assign x_34763 = x_34761 & x_34762;
assign x_34764 = x_3473 & x_3474;
assign x_34765 = x_3475 & x_3476;
assign x_34766 = x_34764 & x_34765;
assign x_34767 = x_34763 & x_34766;
assign x_34768 = x_3477 & x_3478;
assign x_34769 = x_3479 & x_3480;
assign x_34770 = x_34768 & x_34769;
assign x_34771 = x_3481 & x_3482;
assign x_34772 = x_3483 & x_3484;
assign x_34773 = x_34771 & x_34772;
assign x_34774 = x_34770 & x_34773;
assign x_34775 = x_34767 & x_34774;
assign x_34776 = x_34760 & x_34775;
assign x_34777 = x_34746 & x_34776;
assign x_34778 = x_3486 & x_3487;
assign x_34779 = x_3485 & x_34778;
assign x_34780 = x_3488 & x_3489;
assign x_34781 = x_3490 & x_3491;
assign x_34782 = x_34780 & x_34781;
assign x_34783 = x_34779 & x_34782;
assign x_34784 = x_3492 & x_3493;
assign x_34785 = x_3494 & x_3495;
assign x_34786 = x_34784 & x_34785;
assign x_34787 = x_3496 & x_3497;
assign x_34788 = x_3498 & x_3499;
assign x_34789 = x_34787 & x_34788;
assign x_34790 = x_34786 & x_34789;
assign x_34791 = x_34783 & x_34790;
assign x_34792 = x_3501 & x_3502;
assign x_34793 = x_3500 & x_34792;
assign x_34794 = x_3503 & x_3504;
assign x_34795 = x_3505 & x_3506;
assign x_34796 = x_34794 & x_34795;
assign x_34797 = x_34793 & x_34796;
assign x_34798 = x_3507 & x_3508;
assign x_34799 = x_3509 & x_3510;
assign x_34800 = x_34798 & x_34799;
assign x_34801 = x_3511 & x_3512;
assign x_34802 = x_3513 & x_3514;
assign x_34803 = x_34801 & x_34802;
assign x_34804 = x_34800 & x_34803;
assign x_34805 = x_34797 & x_34804;
assign x_34806 = x_34791 & x_34805;
assign x_34807 = x_3516 & x_3517;
assign x_34808 = x_3515 & x_34807;
assign x_34809 = x_3518 & x_3519;
assign x_34810 = x_3520 & x_3521;
assign x_34811 = x_34809 & x_34810;
assign x_34812 = x_34808 & x_34811;
assign x_34813 = x_3522 & x_3523;
assign x_34814 = x_3524 & x_3525;
assign x_34815 = x_34813 & x_34814;
assign x_34816 = x_3526 & x_3527;
assign x_34817 = x_3528 & x_3529;
assign x_34818 = x_34816 & x_34817;
assign x_34819 = x_34815 & x_34818;
assign x_34820 = x_34812 & x_34819;
assign x_34821 = x_3530 & x_3531;
assign x_34822 = x_3532 & x_3533;
assign x_34823 = x_34821 & x_34822;
assign x_34824 = x_3534 & x_3535;
assign x_34825 = x_3536 & x_3537;
assign x_34826 = x_34824 & x_34825;
assign x_34827 = x_34823 & x_34826;
assign x_34828 = x_3538 & x_3539;
assign x_34829 = x_3540 & x_3541;
assign x_34830 = x_34828 & x_34829;
assign x_34831 = x_3542 & x_3543;
assign x_34832 = x_3544 & x_3545;
assign x_34833 = x_34831 & x_34832;
assign x_34834 = x_34830 & x_34833;
assign x_34835 = x_34827 & x_34834;
assign x_34836 = x_34820 & x_34835;
assign x_34837 = x_34806 & x_34836;
assign x_34838 = x_34777 & x_34837;
assign x_34839 = x_3547 & x_3548;
assign x_34840 = x_3546 & x_34839;
assign x_34841 = x_3549 & x_3550;
assign x_34842 = x_3551 & x_3552;
assign x_34843 = x_34841 & x_34842;
assign x_34844 = x_34840 & x_34843;
assign x_34845 = x_3553 & x_3554;
assign x_34846 = x_3555 & x_3556;
assign x_34847 = x_34845 & x_34846;
assign x_34848 = x_3557 & x_3558;
assign x_34849 = x_3559 & x_3560;
assign x_34850 = x_34848 & x_34849;
assign x_34851 = x_34847 & x_34850;
assign x_34852 = x_34844 & x_34851;
assign x_34853 = x_3562 & x_3563;
assign x_34854 = x_3561 & x_34853;
assign x_34855 = x_3564 & x_3565;
assign x_34856 = x_3566 & x_3567;
assign x_34857 = x_34855 & x_34856;
assign x_34858 = x_34854 & x_34857;
assign x_34859 = x_3568 & x_3569;
assign x_34860 = x_3570 & x_3571;
assign x_34861 = x_34859 & x_34860;
assign x_34862 = x_3572 & x_3573;
assign x_34863 = x_3574 & x_3575;
assign x_34864 = x_34862 & x_34863;
assign x_34865 = x_34861 & x_34864;
assign x_34866 = x_34858 & x_34865;
assign x_34867 = x_34852 & x_34866;
assign x_34868 = x_3577 & x_3578;
assign x_34869 = x_3576 & x_34868;
assign x_34870 = x_3579 & x_3580;
assign x_34871 = x_3581 & x_3582;
assign x_34872 = x_34870 & x_34871;
assign x_34873 = x_34869 & x_34872;
assign x_34874 = x_3583 & x_3584;
assign x_34875 = x_3585 & x_3586;
assign x_34876 = x_34874 & x_34875;
assign x_34877 = x_3587 & x_3588;
assign x_34878 = x_3589 & x_3590;
assign x_34879 = x_34877 & x_34878;
assign x_34880 = x_34876 & x_34879;
assign x_34881 = x_34873 & x_34880;
assign x_34882 = x_3591 & x_3592;
assign x_34883 = x_3593 & x_3594;
assign x_34884 = x_34882 & x_34883;
assign x_34885 = x_3595 & x_3596;
assign x_34886 = x_3597 & x_3598;
assign x_34887 = x_34885 & x_34886;
assign x_34888 = x_34884 & x_34887;
assign x_34889 = x_3599 & x_3600;
assign x_34890 = x_3601 & x_3602;
assign x_34891 = x_34889 & x_34890;
assign x_34892 = x_3603 & x_3604;
assign x_34893 = x_3605 & x_3606;
assign x_34894 = x_34892 & x_34893;
assign x_34895 = x_34891 & x_34894;
assign x_34896 = x_34888 & x_34895;
assign x_34897 = x_34881 & x_34896;
assign x_34898 = x_34867 & x_34897;
assign x_34899 = x_3608 & x_3609;
assign x_34900 = x_3607 & x_34899;
assign x_34901 = x_3610 & x_3611;
assign x_34902 = x_3612 & x_3613;
assign x_34903 = x_34901 & x_34902;
assign x_34904 = x_34900 & x_34903;
assign x_34905 = x_3614 & x_3615;
assign x_34906 = x_3616 & x_3617;
assign x_34907 = x_34905 & x_34906;
assign x_34908 = x_3618 & x_3619;
assign x_34909 = x_3620 & x_3621;
assign x_34910 = x_34908 & x_34909;
assign x_34911 = x_34907 & x_34910;
assign x_34912 = x_34904 & x_34911;
assign x_34913 = x_3623 & x_3624;
assign x_34914 = x_3622 & x_34913;
assign x_34915 = x_3625 & x_3626;
assign x_34916 = x_3627 & x_3628;
assign x_34917 = x_34915 & x_34916;
assign x_34918 = x_34914 & x_34917;
assign x_34919 = x_3629 & x_3630;
assign x_34920 = x_3631 & x_3632;
assign x_34921 = x_34919 & x_34920;
assign x_34922 = x_3633 & x_3634;
assign x_34923 = x_3635 & x_3636;
assign x_34924 = x_34922 & x_34923;
assign x_34925 = x_34921 & x_34924;
assign x_34926 = x_34918 & x_34925;
assign x_34927 = x_34912 & x_34926;
assign x_34928 = x_3638 & x_3639;
assign x_34929 = x_3637 & x_34928;
assign x_34930 = x_3640 & x_3641;
assign x_34931 = x_3642 & x_3643;
assign x_34932 = x_34930 & x_34931;
assign x_34933 = x_34929 & x_34932;
assign x_34934 = x_3644 & x_3645;
assign x_34935 = x_3646 & x_3647;
assign x_34936 = x_34934 & x_34935;
assign x_34937 = x_3648 & x_3649;
assign x_34938 = x_3650 & x_3651;
assign x_34939 = x_34937 & x_34938;
assign x_34940 = x_34936 & x_34939;
assign x_34941 = x_34933 & x_34940;
assign x_34942 = x_3652 & x_3653;
assign x_34943 = x_3654 & x_3655;
assign x_34944 = x_34942 & x_34943;
assign x_34945 = x_3656 & x_3657;
assign x_34946 = x_3658 & x_3659;
assign x_34947 = x_34945 & x_34946;
assign x_34948 = x_34944 & x_34947;
assign x_34949 = x_3660 & x_3661;
assign x_34950 = x_3662 & x_3663;
assign x_34951 = x_34949 & x_34950;
assign x_34952 = x_3664 & x_3665;
assign x_34953 = x_3666 & x_3667;
assign x_34954 = x_34952 & x_34953;
assign x_34955 = x_34951 & x_34954;
assign x_34956 = x_34948 & x_34955;
assign x_34957 = x_34941 & x_34956;
assign x_34958 = x_34927 & x_34957;
assign x_34959 = x_34898 & x_34958;
assign x_34960 = x_34838 & x_34959;
assign x_34961 = x_3669 & x_3670;
assign x_34962 = x_3668 & x_34961;
assign x_34963 = x_3671 & x_3672;
assign x_34964 = x_3673 & x_3674;
assign x_34965 = x_34963 & x_34964;
assign x_34966 = x_34962 & x_34965;
assign x_34967 = x_3675 & x_3676;
assign x_34968 = x_3677 & x_3678;
assign x_34969 = x_34967 & x_34968;
assign x_34970 = x_3679 & x_3680;
assign x_34971 = x_3681 & x_3682;
assign x_34972 = x_34970 & x_34971;
assign x_34973 = x_34969 & x_34972;
assign x_34974 = x_34966 & x_34973;
assign x_34975 = x_3684 & x_3685;
assign x_34976 = x_3683 & x_34975;
assign x_34977 = x_3686 & x_3687;
assign x_34978 = x_3688 & x_3689;
assign x_34979 = x_34977 & x_34978;
assign x_34980 = x_34976 & x_34979;
assign x_34981 = x_3690 & x_3691;
assign x_34982 = x_3692 & x_3693;
assign x_34983 = x_34981 & x_34982;
assign x_34984 = x_3694 & x_3695;
assign x_34985 = x_3696 & x_3697;
assign x_34986 = x_34984 & x_34985;
assign x_34987 = x_34983 & x_34986;
assign x_34988 = x_34980 & x_34987;
assign x_34989 = x_34974 & x_34988;
assign x_34990 = x_3699 & x_3700;
assign x_34991 = x_3698 & x_34990;
assign x_34992 = x_3701 & x_3702;
assign x_34993 = x_3703 & x_3704;
assign x_34994 = x_34992 & x_34993;
assign x_34995 = x_34991 & x_34994;
assign x_34996 = x_3705 & x_3706;
assign x_34997 = x_3707 & x_3708;
assign x_34998 = x_34996 & x_34997;
assign x_34999 = x_3709 & x_3710;
assign x_35000 = x_3711 & x_3712;
assign x_35001 = x_34999 & x_35000;
assign x_35002 = x_34998 & x_35001;
assign x_35003 = x_34995 & x_35002;
assign x_35004 = x_3713 & x_3714;
assign x_35005 = x_3715 & x_3716;
assign x_35006 = x_35004 & x_35005;
assign x_35007 = x_3717 & x_3718;
assign x_35008 = x_3719 & x_3720;
assign x_35009 = x_35007 & x_35008;
assign x_35010 = x_35006 & x_35009;
assign x_35011 = x_3721 & x_3722;
assign x_35012 = x_3723 & x_3724;
assign x_35013 = x_35011 & x_35012;
assign x_35014 = x_3725 & x_3726;
assign x_35015 = x_3727 & x_3728;
assign x_35016 = x_35014 & x_35015;
assign x_35017 = x_35013 & x_35016;
assign x_35018 = x_35010 & x_35017;
assign x_35019 = x_35003 & x_35018;
assign x_35020 = x_34989 & x_35019;
assign x_35021 = x_3730 & x_3731;
assign x_35022 = x_3729 & x_35021;
assign x_35023 = x_3732 & x_3733;
assign x_35024 = x_3734 & x_3735;
assign x_35025 = x_35023 & x_35024;
assign x_35026 = x_35022 & x_35025;
assign x_35027 = x_3736 & x_3737;
assign x_35028 = x_3738 & x_3739;
assign x_35029 = x_35027 & x_35028;
assign x_35030 = x_3740 & x_3741;
assign x_35031 = x_3742 & x_3743;
assign x_35032 = x_35030 & x_35031;
assign x_35033 = x_35029 & x_35032;
assign x_35034 = x_35026 & x_35033;
assign x_35035 = x_3745 & x_3746;
assign x_35036 = x_3744 & x_35035;
assign x_35037 = x_3747 & x_3748;
assign x_35038 = x_3749 & x_3750;
assign x_35039 = x_35037 & x_35038;
assign x_35040 = x_35036 & x_35039;
assign x_35041 = x_3751 & x_3752;
assign x_35042 = x_3753 & x_3754;
assign x_35043 = x_35041 & x_35042;
assign x_35044 = x_3755 & x_3756;
assign x_35045 = x_3757 & x_3758;
assign x_35046 = x_35044 & x_35045;
assign x_35047 = x_35043 & x_35046;
assign x_35048 = x_35040 & x_35047;
assign x_35049 = x_35034 & x_35048;
assign x_35050 = x_3760 & x_3761;
assign x_35051 = x_3759 & x_35050;
assign x_35052 = x_3762 & x_3763;
assign x_35053 = x_3764 & x_3765;
assign x_35054 = x_35052 & x_35053;
assign x_35055 = x_35051 & x_35054;
assign x_35056 = x_3766 & x_3767;
assign x_35057 = x_3768 & x_3769;
assign x_35058 = x_35056 & x_35057;
assign x_35059 = x_3770 & x_3771;
assign x_35060 = x_3772 & x_3773;
assign x_35061 = x_35059 & x_35060;
assign x_35062 = x_35058 & x_35061;
assign x_35063 = x_35055 & x_35062;
assign x_35064 = x_3774 & x_3775;
assign x_35065 = x_3776 & x_3777;
assign x_35066 = x_35064 & x_35065;
assign x_35067 = x_3778 & x_3779;
assign x_35068 = x_3780 & x_3781;
assign x_35069 = x_35067 & x_35068;
assign x_35070 = x_35066 & x_35069;
assign x_35071 = x_3782 & x_3783;
assign x_35072 = x_3784 & x_3785;
assign x_35073 = x_35071 & x_35072;
assign x_35074 = x_3786 & x_3787;
assign x_35075 = x_3788 & x_3789;
assign x_35076 = x_35074 & x_35075;
assign x_35077 = x_35073 & x_35076;
assign x_35078 = x_35070 & x_35077;
assign x_35079 = x_35063 & x_35078;
assign x_35080 = x_35049 & x_35079;
assign x_35081 = x_35020 & x_35080;
assign x_35082 = x_3791 & x_3792;
assign x_35083 = x_3790 & x_35082;
assign x_35084 = x_3793 & x_3794;
assign x_35085 = x_3795 & x_3796;
assign x_35086 = x_35084 & x_35085;
assign x_35087 = x_35083 & x_35086;
assign x_35088 = x_3797 & x_3798;
assign x_35089 = x_3799 & x_3800;
assign x_35090 = x_35088 & x_35089;
assign x_35091 = x_3801 & x_3802;
assign x_35092 = x_3803 & x_3804;
assign x_35093 = x_35091 & x_35092;
assign x_35094 = x_35090 & x_35093;
assign x_35095 = x_35087 & x_35094;
assign x_35096 = x_3806 & x_3807;
assign x_35097 = x_3805 & x_35096;
assign x_35098 = x_3808 & x_3809;
assign x_35099 = x_3810 & x_3811;
assign x_35100 = x_35098 & x_35099;
assign x_35101 = x_35097 & x_35100;
assign x_35102 = x_3812 & x_3813;
assign x_35103 = x_3814 & x_3815;
assign x_35104 = x_35102 & x_35103;
assign x_35105 = x_3816 & x_3817;
assign x_35106 = x_3818 & x_3819;
assign x_35107 = x_35105 & x_35106;
assign x_35108 = x_35104 & x_35107;
assign x_35109 = x_35101 & x_35108;
assign x_35110 = x_35095 & x_35109;
assign x_35111 = x_3821 & x_3822;
assign x_35112 = x_3820 & x_35111;
assign x_35113 = x_3823 & x_3824;
assign x_35114 = x_3825 & x_3826;
assign x_35115 = x_35113 & x_35114;
assign x_35116 = x_35112 & x_35115;
assign x_35117 = x_3827 & x_3828;
assign x_35118 = x_3829 & x_3830;
assign x_35119 = x_35117 & x_35118;
assign x_35120 = x_3831 & x_3832;
assign x_35121 = x_3833 & x_3834;
assign x_35122 = x_35120 & x_35121;
assign x_35123 = x_35119 & x_35122;
assign x_35124 = x_35116 & x_35123;
assign x_35125 = x_3835 & x_3836;
assign x_35126 = x_3837 & x_3838;
assign x_35127 = x_35125 & x_35126;
assign x_35128 = x_3839 & x_3840;
assign x_35129 = x_3841 & x_3842;
assign x_35130 = x_35128 & x_35129;
assign x_35131 = x_35127 & x_35130;
assign x_35132 = x_3843 & x_3844;
assign x_35133 = x_3845 & x_3846;
assign x_35134 = x_35132 & x_35133;
assign x_35135 = x_3847 & x_3848;
assign x_35136 = x_3849 & x_3850;
assign x_35137 = x_35135 & x_35136;
assign x_35138 = x_35134 & x_35137;
assign x_35139 = x_35131 & x_35138;
assign x_35140 = x_35124 & x_35139;
assign x_35141 = x_35110 & x_35140;
assign x_35142 = x_3852 & x_3853;
assign x_35143 = x_3851 & x_35142;
assign x_35144 = x_3854 & x_3855;
assign x_35145 = x_3856 & x_3857;
assign x_35146 = x_35144 & x_35145;
assign x_35147 = x_35143 & x_35146;
assign x_35148 = x_3858 & x_3859;
assign x_35149 = x_3860 & x_3861;
assign x_35150 = x_35148 & x_35149;
assign x_35151 = x_3862 & x_3863;
assign x_35152 = x_3864 & x_3865;
assign x_35153 = x_35151 & x_35152;
assign x_35154 = x_35150 & x_35153;
assign x_35155 = x_35147 & x_35154;
assign x_35156 = x_3866 & x_3867;
assign x_35157 = x_3868 & x_3869;
assign x_35158 = x_35156 & x_35157;
assign x_35159 = x_3870 & x_3871;
assign x_35160 = x_3872 & x_3873;
assign x_35161 = x_35159 & x_35160;
assign x_35162 = x_35158 & x_35161;
assign x_35163 = x_3874 & x_3875;
assign x_35164 = x_3876 & x_3877;
assign x_35165 = x_35163 & x_35164;
assign x_35166 = x_3878 & x_3879;
assign x_35167 = x_3880 & x_3881;
assign x_35168 = x_35166 & x_35167;
assign x_35169 = x_35165 & x_35168;
assign x_35170 = x_35162 & x_35169;
assign x_35171 = x_35155 & x_35170;
assign x_35172 = x_3883 & x_3884;
assign x_35173 = x_3882 & x_35172;
assign x_35174 = x_3885 & x_3886;
assign x_35175 = x_3887 & x_3888;
assign x_35176 = x_35174 & x_35175;
assign x_35177 = x_35173 & x_35176;
assign x_35178 = x_3889 & x_3890;
assign x_35179 = x_3891 & x_3892;
assign x_35180 = x_35178 & x_35179;
assign x_35181 = x_3893 & x_3894;
assign x_35182 = x_3895 & x_3896;
assign x_35183 = x_35181 & x_35182;
assign x_35184 = x_35180 & x_35183;
assign x_35185 = x_35177 & x_35184;
assign x_35186 = x_3897 & x_3898;
assign x_35187 = x_3899 & x_3900;
assign x_35188 = x_35186 & x_35187;
assign x_35189 = x_3901 & x_3902;
assign x_35190 = x_3903 & x_3904;
assign x_35191 = x_35189 & x_35190;
assign x_35192 = x_35188 & x_35191;
assign x_35193 = x_3905 & x_3906;
assign x_35194 = x_3907 & x_3908;
assign x_35195 = x_35193 & x_35194;
assign x_35196 = x_3909 & x_3910;
assign x_35197 = x_3911 & x_3912;
assign x_35198 = x_35196 & x_35197;
assign x_35199 = x_35195 & x_35198;
assign x_35200 = x_35192 & x_35199;
assign x_35201 = x_35185 & x_35200;
assign x_35202 = x_35171 & x_35201;
assign x_35203 = x_35141 & x_35202;
assign x_35204 = x_35081 & x_35203;
assign x_35205 = x_34960 & x_35204;
assign x_35206 = x_34717 & x_35205;
assign x_35207 = x_34229 & x_35206;
assign x_35208 = x_33252 & x_35207;
assign x_35209 = x_3914 & x_3915;
assign x_35210 = x_3913 & x_35209;
assign x_35211 = x_3916 & x_3917;
assign x_35212 = x_3918 & x_3919;
assign x_35213 = x_35211 & x_35212;
assign x_35214 = x_35210 & x_35213;
assign x_35215 = x_3920 & x_3921;
assign x_35216 = x_3922 & x_3923;
assign x_35217 = x_35215 & x_35216;
assign x_35218 = x_3924 & x_3925;
assign x_35219 = x_3926 & x_3927;
assign x_35220 = x_35218 & x_35219;
assign x_35221 = x_35217 & x_35220;
assign x_35222 = x_35214 & x_35221;
assign x_35223 = x_3929 & x_3930;
assign x_35224 = x_3928 & x_35223;
assign x_35225 = x_3931 & x_3932;
assign x_35226 = x_3933 & x_3934;
assign x_35227 = x_35225 & x_35226;
assign x_35228 = x_35224 & x_35227;
assign x_35229 = x_3935 & x_3936;
assign x_35230 = x_3937 & x_3938;
assign x_35231 = x_35229 & x_35230;
assign x_35232 = x_3939 & x_3940;
assign x_35233 = x_3941 & x_3942;
assign x_35234 = x_35232 & x_35233;
assign x_35235 = x_35231 & x_35234;
assign x_35236 = x_35228 & x_35235;
assign x_35237 = x_35222 & x_35236;
assign x_35238 = x_3944 & x_3945;
assign x_35239 = x_3943 & x_35238;
assign x_35240 = x_3946 & x_3947;
assign x_35241 = x_3948 & x_3949;
assign x_35242 = x_35240 & x_35241;
assign x_35243 = x_35239 & x_35242;
assign x_35244 = x_3950 & x_3951;
assign x_35245 = x_3952 & x_3953;
assign x_35246 = x_35244 & x_35245;
assign x_35247 = x_3954 & x_3955;
assign x_35248 = x_3956 & x_3957;
assign x_35249 = x_35247 & x_35248;
assign x_35250 = x_35246 & x_35249;
assign x_35251 = x_35243 & x_35250;
assign x_35252 = x_3958 & x_3959;
assign x_35253 = x_3960 & x_3961;
assign x_35254 = x_35252 & x_35253;
assign x_35255 = x_3962 & x_3963;
assign x_35256 = x_3964 & x_3965;
assign x_35257 = x_35255 & x_35256;
assign x_35258 = x_35254 & x_35257;
assign x_35259 = x_3966 & x_3967;
assign x_35260 = x_3968 & x_3969;
assign x_35261 = x_35259 & x_35260;
assign x_35262 = x_3970 & x_3971;
assign x_35263 = x_3972 & x_3973;
assign x_35264 = x_35262 & x_35263;
assign x_35265 = x_35261 & x_35264;
assign x_35266 = x_35258 & x_35265;
assign x_35267 = x_35251 & x_35266;
assign x_35268 = x_35237 & x_35267;
assign x_35269 = x_3975 & x_3976;
assign x_35270 = x_3974 & x_35269;
assign x_35271 = x_3977 & x_3978;
assign x_35272 = x_3979 & x_3980;
assign x_35273 = x_35271 & x_35272;
assign x_35274 = x_35270 & x_35273;
assign x_35275 = x_3981 & x_3982;
assign x_35276 = x_3983 & x_3984;
assign x_35277 = x_35275 & x_35276;
assign x_35278 = x_3985 & x_3986;
assign x_35279 = x_3987 & x_3988;
assign x_35280 = x_35278 & x_35279;
assign x_35281 = x_35277 & x_35280;
assign x_35282 = x_35274 & x_35281;
assign x_35283 = x_3990 & x_3991;
assign x_35284 = x_3989 & x_35283;
assign x_35285 = x_3992 & x_3993;
assign x_35286 = x_3994 & x_3995;
assign x_35287 = x_35285 & x_35286;
assign x_35288 = x_35284 & x_35287;
assign x_35289 = x_3996 & x_3997;
assign x_35290 = x_3998 & x_3999;
assign x_35291 = x_35289 & x_35290;
assign x_35292 = x_4000 & x_4001;
assign x_35293 = x_4002 & x_4003;
assign x_35294 = x_35292 & x_35293;
assign x_35295 = x_35291 & x_35294;
assign x_35296 = x_35288 & x_35295;
assign x_35297 = x_35282 & x_35296;
assign x_35298 = x_4005 & x_4006;
assign x_35299 = x_4004 & x_35298;
assign x_35300 = x_4007 & x_4008;
assign x_35301 = x_4009 & x_4010;
assign x_35302 = x_35300 & x_35301;
assign x_35303 = x_35299 & x_35302;
assign x_35304 = x_4011 & x_4012;
assign x_35305 = x_4013 & x_4014;
assign x_35306 = x_35304 & x_35305;
assign x_35307 = x_4015 & x_4016;
assign x_35308 = x_4017 & x_4018;
assign x_35309 = x_35307 & x_35308;
assign x_35310 = x_35306 & x_35309;
assign x_35311 = x_35303 & x_35310;
assign x_35312 = x_4019 & x_4020;
assign x_35313 = x_4021 & x_4022;
assign x_35314 = x_35312 & x_35313;
assign x_35315 = x_4023 & x_4024;
assign x_35316 = x_4025 & x_4026;
assign x_35317 = x_35315 & x_35316;
assign x_35318 = x_35314 & x_35317;
assign x_35319 = x_4027 & x_4028;
assign x_35320 = x_4029 & x_4030;
assign x_35321 = x_35319 & x_35320;
assign x_35322 = x_4031 & x_4032;
assign x_35323 = x_4033 & x_4034;
assign x_35324 = x_35322 & x_35323;
assign x_35325 = x_35321 & x_35324;
assign x_35326 = x_35318 & x_35325;
assign x_35327 = x_35311 & x_35326;
assign x_35328 = x_35297 & x_35327;
assign x_35329 = x_35268 & x_35328;
assign x_35330 = x_4036 & x_4037;
assign x_35331 = x_4035 & x_35330;
assign x_35332 = x_4038 & x_4039;
assign x_35333 = x_4040 & x_4041;
assign x_35334 = x_35332 & x_35333;
assign x_35335 = x_35331 & x_35334;
assign x_35336 = x_4042 & x_4043;
assign x_35337 = x_4044 & x_4045;
assign x_35338 = x_35336 & x_35337;
assign x_35339 = x_4046 & x_4047;
assign x_35340 = x_4048 & x_4049;
assign x_35341 = x_35339 & x_35340;
assign x_35342 = x_35338 & x_35341;
assign x_35343 = x_35335 & x_35342;
assign x_35344 = x_4051 & x_4052;
assign x_35345 = x_4050 & x_35344;
assign x_35346 = x_4053 & x_4054;
assign x_35347 = x_4055 & x_4056;
assign x_35348 = x_35346 & x_35347;
assign x_35349 = x_35345 & x_35348;
assign x_35350 = x_4057 & x_4058;
assign x_35351 = x_4059 & x_4060;
assign x_35352 = x_35350 & x_35351;
assign x_35353 = x_4061 & x_4062;
assign x_35354 = x_4063 & x_4064;
assign x_35355 = x_35353 & x_35354;
assign x_35356 = x_35352 & x_35355;
assign x_35357 = x_35349 & x_35356;
assign x_35358 = x_35343 & x_35357;
assign x_35359 = x_4066 & x_4067;
assign x_35360 = x_4065 & x_35359;
assign x_35361 = x_4068 & x_4069;
assign x_35362 = x_4070 & x_4071;
assign x_35363 = x_35361 & x_35362;
assign x_35364 = x_35360 & x_35363;
assign x_35365 = x_4072 & x_4073;
assign x_35366 = x_4074 & x_4075;
assign x_35367 = x_35365 & x_35366;
assign x_35368 = x_4076 & x_4077;
assign x_35369 = x_4078 & x_4079;
assign x_35370 = x_35368 & x_35369;
assign x_35371 = x_35367 & x_35370;
assign x_35372 = x_35364 & x_35371;
assign x_35373 = x_4080 & x_4081;
assign x_35374 = x_4082 & x_4083;
assign x_35375 = x_35373 & x_35374;
assign x_35376 = x_4084 & x_4085;
assign x_35377 = x_4086 & x_4087;
assign x_35378 = x_35376 & x_35377;
assign x_35379 = x_35375 & x_35378;
assign x_35380 = x_4088 & x_4089;
assign x_35381 = x_4090 & x_4091;
assign x_35382 = x_35380 & x_35381;
assign x_35383 = x_4092 & x_4093;
assign x_35384 = x_4094 & x_4095;
assign x_35385 = x_35383 & x_35384;
assign x_35386 = x_35382 & x_35385;
assign x_35387 = x_35379 & x_35386;
assign x_35388 = x_35372 & x_35387;
assign x_35389 = x_35358 & x_35388;
assign x_35390 = x_4097 & x_4098;
assign x_35391 = x_4096 & x_35390;
assign x_35392 = x_4099 & x_4100;
assign x_35393 = x_4101 & x_4102;
assign x_35394 = x_35392 & x_35393;
assign x_35395 = x_35391 & x_35394;
assign x_35396 = x_4103 & x_4104;
assign x_35397 = x_4105 & x_4106;
assign x_35398 = x_35396 & x_35397;
assign x_35399 = x_4107 & x_4108;
assign x_35400 = x_4109 & x_4110;
assign x_35401 = x_35399 & x_35400;
assign x_35402 = x_35398 & x_35401;
assign x_35403 = x_35395 & x_35402;
assign x_35404 = x_4112 & x_4113;
assign x_35405 = x_4111 & x_35404;
assign x_35406 = x_4114 & x_4115;
assign x_35407 = x_4116 & x_4117;
assign x_35408 = x_35406 & x_35407;
assign x_35409 = x_35405 & x_35408;
assign x_35410 = x_4118 & x_4119;
assign x_35411 = x_4120 & x_4121;
assign x_35412 = x_35410 & x_35411;
assign x_35413 = x_4122 & x_4123;
assign x_35414 = x_4124 & x_4125;
assign x_35415 = x_35413 & x_35414;
assign x_35416 = x_35412 & x_35415;
assign x_35417 = x_35409 & x_35416;
assign x_35418 = x_35403 & x_35417;
assign x_35419 = x_4127 & x_4128;
assign x_35420 = x_4126 & x_35419;
assign x_35421 = x_4129 & x_4130;
assign x_35422 = x_4131 & x_4132;
assign x_35423 = x_35421 & x_35422;
assign x_35424 = x_35420 & x_35423;
assign x_35425 = x_4133 & x_4134;
assign x_35426 = x_4135 & x_4136;
assign x_35427 = x_35425 & x_35426;
assign x_35428 = x_4137 & x_4138;
assign x_35429 = x_4139 & x_4140;
assign x_35430 = x_35428 & x_35429;
assign x_35431 = x_35427 & x_35430;
assign x_35432 = x_35424 & x_35431;
assign x_35433 = x_4141 & x_4142;
assign x_35434 = x_4143 & x_4144;
assign x_35435 = x_35433 & x_35434;
assign x_35436 = x_4145 & x_4146;
assign x_35437 = x_4147 & x_4148;
assign x_35438 = x_35436 & x_35437;
assign x_35439 = x_35435 & x_35438;
assign x_35440 = x_4149 & x_4150;
assign x_35441 = x_4151 & x_4152;
assign x_35442 = x_35440 & x_35441;
assign x_35443 = x_4153 & x_4154;
assign x_35444 = x_4155 & x_4156;
assign x_35445 = x_35443 & x_35444;
assign x_35446 = x_35442 & x_35445;
assign x_35447 = x_35439 & x_35446;
assign x_35448 = x_35432 & x_35447;
assign x_35449 = x_35418 & x_35448;
assign x_35450 = x_35389 & x_35449;
assign x_35451 = x_35329 & x_35450;
assign x_35452 = x_4158 & x_4159;
assign x_35453 = x_4157 & x_35452;
assign x_35454 = x_4160 & x_4161;
assign x_35455 = x_4162 & x_4163;
assign x_35456 = x_35454 & x_35455;
assign x_35457 = x_35453 & x_35456;
assign x_35458 = x_4164 & x_4165;
assign x_35459 = x_4166 & x_4167;
assign x_35460 = x_35458 & x_35459;
assign x_35461 = x_4168 & x_4169;
assign x_35462 = x_4170 & x_4171;
assign x_35463 = x_35461 & x_35462;
assign x_35464 = x_35460 & x_35463;
assign x_35465 = x_35457 & x_35464;
assign x_35466 = x_4173 & x_4174;
assign x_35467 = x_4172 & x_35466;
assign x_35468 = x_4175 & x_4176;
assign x_35469 = x_4177 & x_4178;
assign x_35470 = x_35468 & x_35469;
assign x_35471 = x_35467 & x_35470;
assign x_35472 = x_4179 & x_4180;
assign x_35473 = x_4181 & x_4182;
assign x_35474 = x_35472 & x_35473;
assign x_35475 = x_4183 & x_4184;
assign x_35476 = x_4185 & x_4186;
assign x_35477 = x_35475 & x_35476;
assign x_35478 = x_35474 & x_35477;
assign x_35479 = x_35471 & x_35478;
assign x_35480 = x_35465 & x_35479;
assign x_35481 = x_4188 & x_4189;
assign x_35482 = x_4187 & x_35481;
assign x_35483 = x_4190 & x_4191;
assign x_35484 = x_4192 & x_4193;
assign x_35485 = x_35483 & x_35484;
assign x_35486 = x_35482 & x_35485;
assign x_35487 = x_4194 & x_4195;
assign x_35488 = x_4196 & x_4197;
assign x_35489 = x_35487 & x_35488;
assign x_35490 = x_4198 & x_4199;
assign x_35491 = x_4200 & x_4201;
assign x_35492 = x_35490 & x_35491;
assign x_35493 = x_35489 & x_35492;
assign x_35494 = x_35486 & x_35493;
assign x_35495 = x_4202 & x_4203;
assign x_35496 = x_4204 & x_4205;
assign x_35497 = x_35495 & x_35496;
assign x_35498 = x_4206 & x_4207;
assign x_35499 = x_4208 & x_4209;
assign x_35500 = x_35498 & x_35499;
assign x_35501 = x_35497 & x_35500;
assign x_35502 = x_4210 & x_4211;
assign x_35503 = x_4212 & x_4213;
assign x_35504 = x_35502 & x_35503;
assign x_35505 = x_4214 & x_4215;
assign x_35506 = x_4216 & x_4217;
assign x_35507 = x_35505 & x_35506;
assign x_35508 = x_35504 & x_35507;
assign x_35509 = x_35501 & x_35508;
assign x_35510 = x_35494 & x_35509;
assign x_35511 = x_35480 & x_35510;
assign x_35512 = x_4219 & x_4220;
assign x_35513 = x_4218 & x_35512;
assign x_35514 = x_4221 & x_4222;
assign x_35515 = x_4223 & x_4224;
assign x_35516 = x_35514 & x_35515;
assign x_35517 = x_35513 & x_35516;
assign x_35518 = x_4225 & x_4226;
assign x_35519 = x_4227 & x_4228;
assign x_35520 = x_35518 & x_35519;
assign x_35521 = x_4229 & x_4230;
assign x_35522 = x_4231 & x_4232;
assign x_35523 = x_35521 & x_35522;
assign x_35524 = x_35520 & x_35523;
assign x_35525 = x_35517 & x_35524;
assign x_35526 = x_4234 & x_4235;
assign x_35527 = x_4233 & x_35526;
assign x_35528 = x_4236 & x_4237;
assign x_35529 = x_4238 & x_4239;
assign x_35530 = x_35528 & x_35529;
assign x_35531 = x_35527 & x_35530;
assign x_35532 = x_4240 & x_4241;
assign x_35533 = x_4242 & x_4243;
assign x_35534 = x_35532 & x_35533;
assign x_35535 = x_4244 & x_4245;
assign x_35536 = x_4246 & x_4247;
assign x_35537 = x_35535 & x_35536;
assign x_35538 = x_35534 & x_35537;
assign x_35539 = x_35531 & x_35538;
assign x_35540 = x_35525 & x_35539;
assign x_35541 = x_4249 & x_4250;
assign x_35542 = x_4248 & x_35541;
assign x_35543 = x_4251 & x_4252;
assign x_35544 = x_4253 & x_4254;
assign x_35545 = x_35543 & x_35544;
assign x_35546 = x_35542 & x_35545;
assign x_35547 = x_4255 & x_4256;
assign x_35548 = x_4257 & x_4258;
assign x_35549 = x_35547 & x_35548;
assign x_35550 = x_4259 & x_4260;
assign x_35551 = x_4261 & x_4262;
assign x_35552 = x_35550 & x_35551;
assign x_35553 = x_35549 & x_35552;
assign x_35554 = x_35546 & x_35553;
assign x_35555 = x_4263 & x_4264;
assign x_35556 = x_4265 & x_4266;
assign x_35557 = x_35555 & x_35556;
assign x_35558 = x_4267 & x_4268;
assign x_35559 = x_4269 & x_4270;
assign x_35560 = x_35558 & x_35559;
assign x_35561 = x_35557 & x_35560;
assign x_35562 = x_4271 & x_4272;
assign x_35563 = x_4273 & x_4274;
assign x_35564 = x_35562 & x_35563;
assign x_35565 = x_4275 & x_4276;
assign x_35566 = x_4277 & x_4278;
assign x_35567 = x_35565 & x_35566;
assign x_35568 = x_35564 & x_35567;
assign x_35569 = x_35561 & x_35568;
assign x_35570 = x_35554 & x_35569;
assign x_35571 = x_35540 & x_35570;
assign x_35572 = x_35511 & x_35571;
assign x_35573 = x_4280 & x_4281;
assign x_35574 = x_4279 & x_35573;
assign x_35575 = x_4282 & x_4283;
assign x_35576 = x_4284 & x_4285;
assign x_35577 = x_35575 & x_35576;
assign x_35578 = x_35574 & x_35577;
assign x_35579 = x_4286 & x_4287;
assign x_35580 = x_4288 & x_4289;
assign x_35581 = x_35579 & x_35580;
assign x_35582 = x_4290 & x_4291;
assign x_35583 = x_4292 & x_4293;
assign x_35584 = x_35582 & x_35583;
assign x_35585 = x_35581 & x_35584;
assign x_35586 = x_35578 & x_35585;
assign x_35587 = x_4295 & x_4296;
assign x_35588 = x_4294 & x_35587;
assign x_35589 = x_4297 & x_4298;
assign x_35590 = x_4299 & x_4300;
assign x_35591 = x_35589 & x_35590;
assign x_35592 = x_35588 & x_35591;
assign x_35593 = x_4301 & x_4302;
assign x_35594 = x_4303 & x_4304;
assign x_35595 = x_35593 & x_35594;
assign x_35596 = x_4305 & x_4306;
assign x_35597 = x_4307 & x_4308;
assign x_35598 = x_35596 & x_35597;
assign x_35599 = x_35595 & x_35598;
assign x_35600 = x_35592 & x_35599;
assign x_35601 = x_35586 & x_35600;
assign x_35602 = x_4310 & x_4311;
assign x_35603 = x_4309 & x_35602;
assign x_35604 = x_4312 & x_4313;
assign x_35605 = x_4314 & x_4315;
assign x_35606 = x_35604 & x_35605;
assign x_35607 = x_35603 & x_35606;
assign x_35608 = x_4316 & x_4317;
assign x_35609 = x_4318 & x_4319;
assign x_35610 = x_35608 & x_35609;
assign x_35611 = x_4320 & x_4321;
assign x_35612 = x_4322 & x_4323;
assign x_35613 = x_35611 & x_35612;
assign x_35614 = x_35610 & x_35613;
assign x_35615 = x_35607 & x_35614;
assign x_35616 = x_4324 & x_4325;
assign x_35617 = x_4326 & x_4327;
assign x_35618 = x_35616 & x_35617;
assign x_35619 = x_4328 & x_4329;
assign x_35620 = x_4330 & x_4331;
assign x_35621 = x_35619 & x_35620;
assign x_35622 = x_35618 & x_35621;
assign x_35623 = x_4332 & x_4333;
assign x_35624 = x_4334 & x_4335;
assign x_35625 = x_35623 & x_35624;
assign x_35626 = x_4336 & x_4337;
assign x_35627 = x_4338 & x_4339;
assign x_35628 = x_35626 & x_35627;
assign x_35629 = x_35625 & x_35628;
assign x_35630 = x_35622 & x_35629;
assign x_35631 = x_35615 & x_35630;
assign x_35632 = x_35601 & x_35631;
assign x_35633 = x_4341 & x_4342;
assign x_35634 = x_4340 & x_35633;
assign x_35635 = x_4343 & x_4344;
assign x_35636 = x_4345 & x_4346;
assign x_35637 = x_35635 & x_35636;
assign x_35638 = x_35634 & x_35637;
assign x_35639 = x_4347 & x_4348;
assign x_35640 = x_4349 & x_4350;
assign x_35641 = x_35639 & x_35640;
assign x_35642 = x_4351 & x_4352;
assign x_35643 = x_4353 & x_4354;
assign x_35644 = x_35642 & x_35643;
assign x_35645 = x_35641 & x_35644;
assign x_35646 = x_35638 & x_35645;
assign x_35647 = x_4355 & x_4356;
assign x_35648 = x_4357 & x_4358;
assign x_35649 = x_35647 & x_35648;
assign x_35650 = x_4359 & x_4360;
assign x_35651 = x_4361 & x_4362;
assign x_35652 = x_35650 & x_35651;
assign x_35653 = x_35649 & x_35652;
assign x_35654 = x_4363 & x_4364;
assign x_35655 = x_4365 & x_4366;
assign x_35656 = x_35654 & x_35655;
assign x_35657 = x_4367 & x_4368;
assign x_35658 = x_4369 & x_4370;
assign x_35659 = x_35657 & x_35658;
assign x_35660 = x_35656 & x_35659;
assign x_35661 = x_35653 & x_35660;
assign x_35662 = x_35646 & x_35661;
assign x_35663 = x_4372 & x_4373;
assign x_35664 = x_4371 & x_35663;
assign x_35665 = x_4374 & x_4375;
assign x_35666 = x_4376 & x_4377;
assign x_35667 = x_35665 & x_35666;
assign x_35668 = x_35664 & x_35667;
assign x_35669 = x_4378 & x_4379;
assign x_35670 = x_4380 & x_4381;
assign x_35671 = x_35669 & x_35670;
assign x_35672 = x_4382 & x_4383;
assign x_35673 = x_4384 & x_4385;
assign x_35674 = x_35672 & x_35673;
assign x_35675 = x_35671 & x_35674;
assign x_35676 = x_35668 & x_35675;
assign x_35677 = x_4386 & x_4387;
assign x_35678 = x_4388 & x_4389;
assign x_35679 = x_35677 & x_35678;
assign x_35680 = x_4390 & x_4391;
assign x_35681 = x_4392 & x_4393;
assign x_35682 = x_35680 & x_35681;
assign x_35683 = x_35679 & x_35682;
assign x_35684 = x_4394 & x_4395;
assign x_35685 = x_4396 & x_4397;
assign x_35686 = x_35684 & x_35685;
assign x_35687 = x_4398 & x_4399;
assign x_35688 = x_4400 & x_4401;
assign x_35689 = x_35687 & x_35688;
assign x_35690 = x_35686 & x_35689;
assign x_35691 = x_35683 & x_35690;
assign x_35692 = x_35676 & x_35691;
assign x_35693 = x_35662 & x_35692;
assign x_35694 = x_35632 & x_35693;
assign x_35695 = x_35572 & x_35694;
assign x_35696 = x_35451 & x_35695;
assign x_35697 = x_4403 & x_4404;
assign x_35698 = x_4402 & x_35697;
assign x_35699 = x_4405 & x_4406;
assign x_35700 = x_4407 & x_4408;
assign x_35701 = x_35699 & x_35700;
assign x_35702 = x_35698 & x_35701;
assign x_35703 = x_4409 & x_4410;
assign x_35704 = x_4411 & x_4412;
assign x_35705 = x_35703 & x_35704;
assign x_35706 = x_4413 & x_4414;
assign x_35707 = x_4415 & x_4416;
assign x_35708 = x_35706 & x_35707;
assign x_35709 = x_35705 & x_35708;
assign x_35710 = x_35702 & x_35709;
assign x_35711 = x_4418 & x_4419;
assign x_35712 = x_4417 & x_35711;
assign x_35713 = x_4420 & x_4421;
assign x_35714 = x_4422 & x_4423;
assign x_35715 = x_35713 & x_35714;
assign x_35716 = x_35712 & x_35715;
assign x_35717 = x_4424 & x_4425;
assign x_35718 = x_4426 & x_4427;
assign x_35719 = x_35717 & x_35718;
assign x_35720 = x_4428 & x_4429;
assign x_35721 = x_4430 & x_4431;
assign x_35722 = x_35720 & x_35721;
assign x_35723 = x_35719 & x_35722;
assign x_35724 = x_35716 & x_35723;
assign x_35725 = x_35710 & x_35724;
assign x_35726 = x_4433 & x_4434;
assign x_35727 = x_4432 & x_35726;
assign x_35728 = x_4435 & x_4436;
assign x_35729 = x_4437 & x_4438;
assign x_35730 = x_35728 & x_35729;
assign x_35731 = x_35727 & x_35730;
assign x_35732 = x_4439 & x_4440;
assign x_35733 = x_4441 & x_4442;
assign x_35734 = x_35732 & x_35733;
assign x_35735 = x_4443 & x_4444;
assign x_35736 = x_4445 & x_4446;
assign x_35737 = x_35735 & x_35736;
assign x_35738 = x_35734 & x_35737;
assign x_35739 = x_35731 & x_35738;
assign x_35740 = x_4447 & x_4448;
assign x_35741 = x_4449 & x_4450;
assign x_35742 = x_35740 & x_35741;
assign x_35743 = x_4451 & x_4452;
assign x_35744 = x_4453 & x_4454;
assign x_35745 = x_35743 & x_35744;
assign x_35746 = x_35742 & x_35745;
assign x_35747 = x_4455 & x_4456;
assign x_35748 = x_4457 & x_4458;
assign x_35749 = x_35747 & x_35748;
assign x_35750 = x_4459 & x_4460;
assign x_35751 = x_4461 & x_4462;
assign x_35752 = x_35750 & x_35751;
assign x_35753 = x_35749 & x_35752;
assign x_35754 = x_35746 & x_35753;
assign x_35755 = x_35739 & x_35754;
assign x_35756 = x_35725 & x_35755;
assign x_35757 = x_4464 & x_4465;
assign x_35758 = x_4463 & x_35757;
assign x_35759 = x_4466 & x_4467;
assign x_35760 = x_4468 & x_4469;
assign x_35761 = x_35759 & x_35760;
assign x_35762 = x_35758 & x_35761;
assign x_35763 = x_4470 & x_4471;
assign x_35764 = x_4472 & x_4473;
assign x_35765 = x_35763 & x_35764;
assign x_35766 = x_4474 & x_4475;
assign x_35767 = x_4476 & x_4477;
assign x_35768 = x_35766 & x_35767;
assign x_35769 = x_35765 & x_35768;
assign x_35770 = x_35762 & x_35769;
assign x_35771 = x_4479 & x_4480;
assign x_35772 = x_4478 & x_35771;
assign x_35773 = x_4481 & x_4482;
assign x_35774 = x_4483 & x_4484;
assign x_35775 = x_35773 & x_35774;
assign x_35776 = x_35772 & x_35775;
assign x_35777 = x_4485 & x_4486;
assign x_35778 = x_4487 & x_4488;
assign x_35779 = x_35777 & x_35778;
assign x_35780 = x_4489 & x_4490;
assign x_35781 = x_4491 & x_4492;
assign x_35782 = x_35780 & x_35781;
assign x_35783 = x_35779 & x_35782;
assign x_35784 = x_35776 & x_35783;
assign x_35785 = x_35770 & x_35784;
assign x_35786 = x_4494 & x_4495;
assign x_35787 = x_4493 & x_35786;
assign x_35788 = x_4496 & x_4497;
assign x_35789 = x_4498 & x_4499;
assign x_35790 = x_35788 & x_35789;
assign x_35791 = x_35787 & x_35790;
assign x_35792 = x_4500 & x_4501;
assign x_35793 = x_4502 & x_4503;
assign x_35794 = x_35792 & x_35793;
assign x_35795 = x_4504 & x_4505;
assign x_35796 = x_4506 & x_4507;
assign x_35797 = x_35795 & x_35796;
assign x_35798 = x_35794 & x_35797;
assign x_35799 = x_35791 & x_35798;
assign x_35800 = x_4508 & x_4509;
assign x_35801 = x_4510 & x_4511;
assign x_35802 = x_35800 & x_35801;
assign x_35803 = x_4512 & x_4513;
assign x_35804 = x_4514 & x_4515;
assign x_35805 = x_35803 & x_35804;
assign x_35806 = x_35802 & x_35805;
assign x_35807 = x_4516 & x_4517;
assign x_35808 = x_4518 & x_4519;
assign x_35809 = x_35807 & x_35808;
assign x_35810 = x_4520 & x_4521;
assign x_35811 = x_4522 & x_4523;
assign x_35812 = x_35810 & x_35811;
assign x_35813 = x_35809 & x_35812;
assign x_35814 = x_35806 & x_35813;
assign x_35815 = x_35799 & x_35814;
assign x_35816 = x_35785 & x_35815;
assign x_35817 = x_35756 & x_35816;
assign x_35818 = x_4525 & x_4526;
assign x_35819 = x_4524 & x_35818;
assign x_35820 = x_4527 & x_4528;
assign x_35821 = x_4529 & x_4530;
assign x_35822 = x_35820 & x_35821;
assign x_35823 = x_35819 & x_35822;
assign x_35824 = x_4531 & x_4532;
assign x_35825 = x_4533 & x_4534;
assign x_35826 = x_35824 & x_35825;
assign x_35827 = x_4535 & x_4536;
assign x_35828 = x_4537 & x_4538;
assign x_35829 = x_35827 & x_35828;
assign x_35830 = x_35826 & x_35829;
assign x_35831 = x_35823 & x_35830;
assign x_35832 = x_4540 & x_4541;
assign x_35833 = x_4539 & x_35832;
assign x_35834 = x_4542 & x_4543;
assign x_35835 = x_4544 & x_4545;
assign x_35836 = x_35834 & x_35835;
assign x_35837 = x_35833 & x_35836;
assign x_35838 = x_4546 & x_4547;
assign x_35839 = x_4548 & x_4549;
assign x_35840 = x_35838 & x_35839;
assign x_35841 = x_4550 & x_4551;
assign x_35842 = x_4552 & x_4553;
assign x_35843 = x_35841 & x_35842;
assign x_35844 = x_35840 & x_35843;
assign x_35845 = x_35837 & x_35844;
assign x_35846 = x_35831 & x_35845;
assign x_35847 = x_4555 & x_4556;
assign x_35848 = x_4554 & x_35847;
assign x_35849 = x_4557 & x_4558;
assign x_35850 = x_4559 & x_4560;
assign x_35851 = x_35849 & x_35850;
assign x_35852 = x_35848 & x_35851;
assign x_35853 = x_4561 & x_4562;
assign x_35854 = x_4563 & x_4564;
assign x_35855 = x_35853 & x_35854;
assign x_35856 = x_4565 & x_4566;
assign x_35857 = x_4567 & x_4568;
assign x_35858 = x_35856 & x_35857;
assign x_35859 = x_35855 & x_35858;
assign x_35860 = x_35852 & x_35859;
assign x_35861 = x_4569 & x_4570;
assign x_35862 = x_4571 & x_4572;
assign x_35863 = x_35861 & x_35862;
assign x_35864 = x_4573 & x_4574;
assign x_35865 = x_4575 & x_4576;
assign x_35866 = x_35864 & x_35865;
assign x_35867 = x_35863 & x_35866;
assign x_35868 = x_4577 & x_4578;
assign x_35869 = x_4579 & x_4580;
assign x_35870 = x_35868 & x_35869;
assign x_35871 = x_4581 & x_4582;
assign x_35872 = x_4583 & x_4584;
assign x_35873 = x_35871 & x_35872;
assign x_35874 = x_35870 & x_35873;
assign x_35875 = x_35867 & x_35874;
assign x_35876 = x_35860 & x_35875;
assign x_35877 = x_35846 & x_35876;
assign x_35878 = x_4586 & x_4587;
assign x_35879 = x_4585 & x_35878;
assign x_35880 = x_4588 & x_4589;
assign x_35881 = x_4590 & x_4591;
assign x_35882 = x_35880 & x_35881;
assign x_35883 = x_35879 & x_35882;
assign x_35884 = x_4592 & x_4593;
assign x_35885 = x_4594 & x_4595;
assign x_35886 = x_35884 & x_35885;
assign x_35887 = x_4596 & x_4597;
assign x_35888 = x_4598 & x_4599;
assign x_35889 = x_35887 & x_35888;
assign x_35890 = x_35886 & x_35889;
assign x_35891 = x_35883 & x_35890;
assign x_35892 = x_4601 & x_4602;
assign x_35893 = x_4600 & x_35892;
assign x_35894 = x_4603 & x_4604;
assign x_35895 = x_4605 & x_4606;
assign x_35896 = x_35894 & x_35895;
assign x_35897 = x_35893 & x_35896;
assign x_35898 = x_4607 & x_4608;
assign x_35899 = x_4609 & x_4610;
assign x_35900 = x_35898 & x_35899;
assign x_35901 = x_4611 & x_4612;
assign x_35902 = x_4613 & x_4614;
assign x_35903 = x_35901 & x_35902;
assign x_35904 = x_35900 & x_35903;
assign x_35905 = x_35897 & x_35904;
assign x_35906 = x_35891 & x_35905;
assign x_35907 = x_4616 & x_4617;
assign x_35908 = x_4615 & x_35907;
assign x_35909 = x_4618 & x_4619;
assign x_35910 = x_4620 & x_4621;
assign x_35911 = x_35909 & x_35910;
assign x_35912 = x_35908 & x_35911;
assign x_35913 = x_4622 & x_4623;
assign x_35914 = x_4624 & x_4625;
assign x_35915 = x_35913 & x_35914;
assign x_35916 = x_4626 & x_4627;
assign x_35917 = x_4628 & x_4629;
assign x_35918 = x_35916 & x_35917;
assign x_35919 = x_35915 & x_35918;
assign x_35920 = x_35912 & x_35919;
assign x_35921 = x_4630 & x_4631;
assign x_35922 = x_4632 & x_4633;
assign x_35923 = x_35921 & x_35922;
assign x_35924 = x_4634 & x_4635;
assign x_35925 = x_4636 & x_4637;
assign x_35926 = x_35924 & x_35925;
assign x_35927 = x_35923 & x_35926;
assign x_35928 = x_4638 & x_4639;
assign x_35929 = x_4640 & x_4641;
assign x_35930 = x_35928 & x_35929;
assign x_35931 = x_4642 & x_4643;
assign x_35932 = x_4644 & x_4645;
assign x_35933 = x_35931 & x_35932;
assign x_35934 = x_35930 & x_35933;
assign x_35935 = x_35927 & x_35934;
assign x_35936 = x_35920 & x_35935;
assign x_35937 = x_35906 & x_35936;
assign x_35938 = x_35877 & x_35937;
assign x_35939 = x_35817 & x_35938;
assign x_35940 = x_4647 & x_4648;
assign x_35941 = x_4646 & x_35940;
assign x_35942 = x_4649 & x_4650;
assign x_35943 = x_4651 & x_4652;
assign x_35944 = x_35942 & x_35943;
assign x_35945 = x_35941 & x_35944;
assign x_35946 = x_4653 & x_4654;
assign x_35947 = x_4655 & x_4656;
assign x_35948 = x_35946 & x_35947;
assign x_35949 = x_4657 & x_4658;
assign x_35950 = x_4659 & x_4660;
assign x_35951 = x_35949 & x_35950;
assign x_35952 = x_35948 & x_35951;
assign x_35953 = x_35945 & x_35952;
assign x_35954 = x_4662 & x_4663;
assign x_35955 = x_4661 & x_35954;
assign x_35956 = x_4664 & x_4665;
assign x_35957 = x_4666 & x_4667;
assign x_35958 = x_35956 & x_35957;
assign x_35959 = x_35955 & x_35958;
assign x_35960 = x_4668 & x_4669;
assign x_35961 = x_4670 & x_4671;
assign x_35962 = x_35960 & x_35961;
assign x_35963 = x_4672 & x_4673;
assign x_35964 = x_4674 & x_4675;
assign x_35965 = x_35963 & x_35964;
assign x_35966 = x_35962 & x_35965;
assign x_35967 = x_35959 & x_35966;
assign x_35968 = x_35953 & x_35967;
assign x_35969 = x_4677 & x_4678;
assign x_35970 = x_4676 & x_35969;
assign x_35971 = x_4679 & x_4680;
assign x_35972 = x_4681 & x_4682;
assign x_35973 = x_35971 & x_35972;
assign x_35974 = x_35970 & x_35973;
assign x_35975 = x_4683 & x_4684;
assign x_35976 = x_4685 & x_4686;
assign x_35977 = x_35975 & x_35976;
assign x_35978 = x_4687 & x_4688;
assign x_35979 = x_4689 & x_4690;
assign x_35980 = x_35978 & x_35979;
assign x_35981 = x_35977 & x_35980;
assign x_35982 = x_35974 & x_35981;
assign x_35983 = x_4691 & x_4692;
assign x_35984 = x_4693 & x_4694;
assign x_35985 = x_35983 & x_35984;
assign x_35986 = x_4695 & x_4696;
assign x_35987 = x_4697 & x_4698;
assign x_35988 = x_35986 & x_35987;
assign x_35989 = x_35985 & x_35988;
assign x_35990 = x_4699 & x_4700;
assign x_35991 = x_4701 & x_4702;
assign x_35992 = x_35990 & x_35991;
assign x_35993 = x_4703 & x_4704;
assign x_35994 = x_4705 & x_4706;
assign x_35995 = x_35993 & x_35994;
assign x_35996 = x_35992 & x_35995;
assign x_35997 = x_35989 & x_35996;
assign x_35998 = x_35982 & x_35997;
assign x_35999 = x_35968 & x_35998;
assign x_36000 = x_4708 & x_4709;
assign x_36001 = x_4707 & x_36000;
assign x_36002 = x_4710 & x_4711;
assign x_36003 = x_4712 & x_4713;
assign x_36004 = x_36002 & x_36003;
assign x_36005 = x_36001 & x_36004;
assign x_36006 = x_4714 & x_4715;
assign x_36007 = x_4716 & x_4717;
assign x_36008 = x_36006 & x_36007;
assign x_36009 = x_4718 & x_4719;
assign x_36010 = x_4720 & x_4721;
assign x_36011 = x_36009 & x_36010;
assign x_36012 = x_36008 & x_36011;
assign x_36013 = x_36005 & x_36012;
assign x_36014 = x_4723 & x_4724;
assign x_36015 = x_4722 & x_36014;
assign x_36016 = x_4725 & x_4726;
assign x_36017 = x_4727 & x_4728;
assign x_36018 = x_36016 & x_36017;
assign x_36019 = x_36015 & x_36018;
assign x_36020 = x_4729 & x_4730;
assign x_36021 = x_4731 & x_4732;
assign x_36022 = x_36020 & x_36021;
assign x_36023 = x_4733 & x_4734;
assign x_36024 = x_4735 & x_4736;
assign x_36025 = x_36023 & x_36024;
assign x_36026 = x_36022 & x_36025;
assign x_36027 = x_36019 & x_36026;
assign x_36028 = x_36013 & x_36027;
assign x_36029 = x_4738 & x_4739;
assign x_36030 = x_4737 & x_36029;
assign x_36031 = x_4740 & x_4741;
assign x_36032 = x_4742 & x_4743;
assign x_36033 = x_36031 & x_36032;
assign x_36034 = x_36030 & x_36033;
assign x_36035 = x_4744 & x_4745;
assign x_36036 = x_4746 & x_4747;
assign x_36037 = x_36035 & x_36036;
assign x_36038 = x_4748 & x_4749;
assign x_36039 = x_4750 & x_4751;
assign x_36040 = x_36038 & x_36039;
assign x_36041 = x_36037 & x_36040;
assign x_36042 = x_36034 & x_36041;
assign x_36043 = x_4752 & x_4753;
assign x_36044 = x_4754 & x_4755;
assign x_36045 = x_36043 & x_36044;
assign x_36046 = x_4756 & x_4757;
assign x_36047 = x_4758 & x_4759;
assign x_36048 = x_36046 & x_36047;
assign x_36049 = x_36045 & x_36048;
assign x_36050 = x_4760 & x_4761;
assign x_36051 = x_4762 & x_4763;
assign x_36052 = x_36050 & x_36051;
assign x_36053 = x_4764 & x_4765;
assign x_36054 = x_4766 & x_4767;
assign x_36055 = x_36053 & x_36054;
assign x_36056 = x_36052 & x_36055;
assign x_36057 = x_36049 & x_36056;
assign x_36058 = x_36042 & x_36057;
assign x_36059 = x_36028 & x_36058;
assign x_36060 = x_35999 & x_36059;
assign x_36061 = x_4769 & x_4770;
assign x_36062 = x_4768 & x_36061;
assign x_36063 = x_4771 & x_4772;
assign x_36064 = x_4773 & x_4774;
assign x_36065 = x_36063 & x_36064;
assign x_36066 = x_36062 & x_36065;
assign x_36067 = x_4775 & x_4776;
assign x_36068 = x_4777 & x_4778;
assign x_36069 = x_36067 & x_36068;
assign x_36070 = x_4779 & x_4780;
assign x_36071 = x_4781 & x_4782;
assign x_36072 = x_36070 & x_36071;
assign x_36073 = x_36069 & x_36072;
assign x_36074 = x_36066 & x_36073;
assign x_36075 = x_4784 & x_4785;
assign x_36076 = x_4783 & x_36075;
assign x_36077 = x_4786 & x_4787;
assign x_36078 = x_4788 & x_4789;
assign x_36079 = x_36077 & x_36078;
assign x_36080 = x_36076 & x_36079;
assign x_36081 = x_4790 & x_4791;
assign x_36082 = x_4792 & x_4793;
assign x_36083 = x_36081 & x_36082;
assign x_36084 = x_4794 & x_4795;
assign x_36085 = x_4796 & x_4797;
assign x_36086 = x_36084 & x_36085;
assign x_36087 = x_36083 & x_36086;
assign x_36088 = x_36080 & x_36087;
assign x_36089 = x_36074 & x_36088;
assign x_36090 = x_4799 & x_4800;
assign x_36091 = x_4798 & x_36090;
assign x_36092 = x_4801 & x_4802;
assign x_36093 = x_4803 & x_4804;
assign x_36094 = x_36092 & x_36093;
assign x_36095 = x_36091 & x_36094;
assign x_36096 = x_4805 & x_4806;
assign x_36097 = x_4807 & x_4808;
assign x_36098 = x_36096 & x_36097;
assign x_36099 = x_4809 & x_4810;
assign x_36100 = x_4811 & x_4812;
assign x_36101 = x_36099 & x_36100;
assign x_36102 = x_36098 & x_36101;
assign x_36103 = x_36095 & x_36102;
assign x_36104 = x_4813 & x_4814;
assign x_36105 = x_4815 & x_4816;
assign x_36106 = x_36104 & x_36105;
assign x_36107 = x_4817 & x_4818;
assign x_36108 = x_4819 & x_4820;
assign x_36109 = x_36107 & x_36108;
assign x_36110 = x_36106 & x_36109;
assign x_36111 = x_4821 & x_4822;
assign x_36112 = x_4823 & x_4824;
assign x_36113 = x_36111 & x_36112;
assign x_36114 = x_4825 & x_4826;
assign x_36115 = x_4827 & x_4828;
assign x_36116 = x_36114 & x_36115;
assign x_36117 = x_36113 & x_36116;
assign x_36118 = x_36110 & x_36117;
assign x_36119 = x_36103 & x_36118;
assign x_36120 = x_36089 & x_36119;
assign x_36121 = x_4830 & x_4831;
assign x_36122 = x_4829 & x_36121;
assign x_36123 = x_4832 & x_4833;
assign x_36124 = x_4834 & x_4835;
assign x_36125 = x_36123 & x_36124;
assign x_36126 = x_36122 & x_36125;
assign x_36127 = x_4836 & x_4837;
assign x_36128 = x_4838 & x_4839;
assign x_36129 = x_36127 & x_36128;
assign x_36130 = x_4840 & x_4841;
assign x_36131 = x_4842 & x_4843;
assign x_36132 = x_36130 & x_36131;
assign x_36133 = x_36129 & x_36132;
assign x_36134 = x_36126 & x_36133;
assign x_36135 = x_4844 & x_4845;
assign x_36136 = x_4846 & x_4847;
assign x_36137 = x_36135 & x_36136;
assign x_36138 = x_4848 & x_4849;
assign x_36139 = x_4850 & x_4851;
assign x_36140 = x_36138 & x_36139;
assign x_36141 = x_36137 & x_36140;
assign x_36142 = x_4852 & x_4853;
assign x_36143 = x_4854 & x_4855;
assign x_36144 = x_36142 & x_36143;
assign x_36145 = x_4856 & x_4857;
assign x_36146 = x_4858 & x_4859;
assign x_36147 = x_36145 & x_36146;
assign x_36148 = x_36144 & x_36147;
assign x_36149 = x_36141 & x_36148;
assign x_36150 = x_36134 & x_36149;
assign x_36151 = x_4861 & x_4862;
assign x_36152 = x_4860 & x_36151;
assign x_36153 = x_4863 & x_4864;
assign x_36154 = x_4865 & x_4866;
assign x_36155 = x_36153 & x_36154;
assign x_36156 = x_36152 & x_36155;
assign x_36157 = x_4867 & x_4868;
assign x_36158 = x_4869 & x_4870;
assign x_36159 = x_36157 & x_36158;
assign x_36160 = x_4871 & x_4872;
assign x_36161 = x_4873 & x_4874;
assign x_36162 = x_36160 & x_36161;
assign x_36163 = x_36159 & x_36162;
assign x_36164 = x_36156 & x_36163;
assign x_36165 = x_4875 & x_4876;
assign x_36166 = x_4877 & x_4878;
assign x_36167 = x_36165 & x_36166;
assign x_36168 = x_4879 & x_4880;
assign x_36169 = x_4881 & x_4882;
assign x_36170 = x_36168 & x_36169;
assign x_36171 = x_36167 & x_36170;
assign x_36172 = x_4883 & x_4884;
assign x_36173 = x_4885 & x_4886;
assign x_36174 = x_36172 & x_36173;
assign x_36175 = x_4887 & x_4888;
assign x_36176 = x_4889 & x_4890;
assign x_36177 = x_36175 & x_36176;
assign x_36178 = x_36174 & x_36177;
assign x_36179 = x_36171 & x_36178;
assign x_36180 = x_36164 & x_36179;
assign x_36181 = x_36150 & x_36180;
assign x_36182 = x_36120 & x_36181;
assign x_36183 = x_36060 & x_36182;
assign x_36184 = x_35939 & x_36183;
assign x_36185 = x_35696 & x_36184;
assign x_36186 = x_4892 & x_4893;
assign x_36187 = x_4891 & x_36186;
assign x_36188 = x_4894 & x_4895;
assign x_36189 = x_4896 & x_4897;
assign x_36190 = x_36188 & x_36189;
assign x_36191 = x_36187 & x_36190;
assign x_36192 = x_4898 & x_4899;
assign x_36193 = x_4900 & x_4901;
assign x_36194 = x_36192 & x_36193;
assign x_36195 = x_4902 & x_4903;
assign x_36196 = x_4904 & x_4905;
assign x_36197 = x_36195 & x_36196;
assign x_36198 = x_36194 & x_36197;
assign x_36199 = x_36191 & x_36198;
assign x_36200 = x_4907 & x_4908;
assign x_36201 = x_4906 & x_36200;
assign x_36202 = x_4909 & x_4910;
assign x_36203 = x_4911 & x_4912;
assign x_36204 = x_36202 & x_36203;
assign x_36205 = x_36201 & x_36204;
assign x_36206 = x_4913 & x_4914;
assign x_36207 = x_4915 & x_4916;
assign x_36208 = x_36206 & x_36207;
assign x_36209 = x_4917 & x_4918;
assign x_36210 = x_4919 & x_4920;
assign x_36211 = x_36209 & x_36210;
assign x_36212 = x_36208 & x_36211;
assign x_36213 = x_36205 & x_36212;
assign x_36214 = x_36199 & x_36213;
assign x_36215 = x_4922 & x_4923;
assign x_36216 = x_4921 & x_36215;
assign x_36217 = x_4924 & x_4925;
assign x_36218 = x_4926 & x_4927;
assign x_36219 = x_36217 & x_36218;
assign x_36220 = x_36216 & x_36219;
assign x_36221 = x_4928 & x_4929;
assign x_36222 = x_4930 & x_4931;
assign x_36223 = x_36221 & x_36222;
assign x_36224 = x_4932 & x_4933;
assign x_36225 = x_4934 & x_4935;
assign x_36226 = x_36224 & x_36225;
assign x_36227 = x_36223 & x_36226;
assign x_36228 = x_36220 & x_36227;
assign x_36229 = x_4936 & x_4937;
assign x_36230 = x_4938 & x_4939;
assign x_36231 = x_36229 & x_36230;
assign x_36232 = x_4940 & x_4941;
assign x_36233 = x_4942 & x_4943;
assign x_36234 = x_36232 & x_36233;
assign x_36235 = x_36231 & x_36234;
assign x_36236 = x_4944 & x_4945;
assign x_36237 = x_4946 & x_4947;
assign x_36238 = x_36236 & x_36237;
assign x_36239 = x_4948 & x_4949;
assign x_36240 = x_4950 & x_4951;
assign x_36241 = x_36239 & x_36240;
assign x_36242 = x_36238 & x_36241;
assign x_36243 = x_36235 & x_36242;
assign x_36244 = x_36228 & x_36243;
assign x_36245 = x_36214 & x_36244;
assign x_36246 = x_4953 & x_4954;
assign x_36247 = x_4952 & x_36246;
assign x_36248 = x_4955 & x_4956;
assign x_36249 = x_4957 & x_4958;
assign x_36250 = x_36248 & x_36249;
assign x_36251 = x_36247 & x_36250;
assign x_36252 = x_4959 & x_4960;
assign x_36253 = x_4961 & x_4962;
assign x_36254 = x_36252 & x_36253;
assign x_36255 = x_4963 & x_4964;
assign x_36256 = x_4965 & x_4966;
assign x_36257 = x_36255 & x_36256;
assign x_36258 = x_36254 & x_36257;
assign x_36259 = x_36251 & x_36258;
assign x_36260 = x_4968 & x_4969;
assign x_36261 = x_4967 & x_36260;
assign x_36262 = x_4970 & x_4971;
assign x_36263 = x_4972 & x_4973;
assign x_36264 = x_36262 & x_36263;
assign x_36265 = x_36261 & x_36264;
assign x_36266 = x_4974 & x_4975;
assign x_36267 = x_4976 & x_4977;
assign x_36268 = x_36266 & x_36267;
assign x_36269 = x_4978 & x_4979;
assign x_36270 = x_4980 & x_4981;
assign x_36271 = x_36269 & x_36270;
assign x_36272 = x_36268 & x_36271;
assign x_36273 = x_36265 & x_36272;
assign x_36274 = x_36259 & x_36273;
assign x_36275 = x_4983 & x_4984;
assign x_36276 = x_4982 & x_36275;
assign x_36277 = x_4985 & x_4986;
assign x_36278 = x_4987 & x_4988;
assign x_36279 = x_36277 & x_36278;
assign x_36280 = x_36276 & x_36279;
assign x_36281 = x_4989 & x_4990;
assign x_36282 = x_4991 & x_4992;
assign x_36283 = x_36281 & x_36282;
assign x_36284 = x_4993 & x_4994;
assign x_36285 = x_4995 & x_4996;
assign x_36286 = x_36284 & x_36285;
assign x_36287 = x_36283 & x_36286;
assign x_36288 = x_36280 & x_36287;
assign x_36289 = x_4997 & x_4998;
assign x_36290 = x_4999 & x_5000;
assign x_36291 = x_36289 & x_36290;
assign x_36292 = x_5001 & x_5002;
assign x_36293 = x_5003 & x_5004;
assign x_36294 = x_36292 & x_36293;
assign x_36295 = x_36291 & x_36294;
assign x_36296 = x_5005 & x_5006;
assign x_36297 = x_5007 & x_5008;
assign x_36298 = x_36296 & x_36297;
assign x_36299 = x_5009 & x_5010;
assign x_36300 = x_5011 & x_5012;
assign x_36301 = x_36299 & x_36300;
assign x_36302 = x_36298 & x_36301;
assign x_36303 = x_36295 & x_36302;
assign x_36304 = x_36288 & x_36303;
assign x_36305 = x_36274 & x_36304;
assign x_36306 = x_36245 & x_36305;
assign x_36307 = x_5014 & x_5015;
assign x_36308 = x_5013 & x_36307;
assign x_36309 = x_5016 & x_5017;
assign x_36310 = x_5018 & x_5019;
assign x_36311 = x_36309 & x_36310;
assign x_36312 = x_36308 & x_36311;
assign x_36313 = x_5020 & x_5021;
assign x_36314 = x_5022 & x_5023;
assign x_36315 = x_36313 & x_36314;
assign x_36316 = x_5024 & x_5025;
assign x_36317 = x_5026 & x_5027;
assign x_36318 = x_36316 & x_36317;
assign x_36319 = x_36315 & x_36318;
assign x_36320 = x_36312 & x_36319;
assign x_36321 = x_5029 & x_5030;
assign x_36322 = x_5028 & x_36321;
assign x_36323 = x_5031 & x_5032;
assign x_36324 = x_5033 & x_5034;
assign x_36325 = x_36323 & x_36324;
assign x_36326 = x_36322 & x_36325;
assign x_36327 = x_5035 & x_5036;
assign x_36328 = x_5037 & x_5038;
assign x_36329 = x_36327 & x_36328;
assign x_36330 = x_5039 & x_5040;
assign x_36331 = x_5041 & x_5042;
assign x_36332 = x_36330 & x_36331;
assign x_36333 = x_36329 & x_36332;
assign x_36334 = x_36326 & x_36333;
assign x_36335 = x_36320 & x_36334;
assign x_36336 = x_5044 & x_5045;
assign x_36337 = x_5043 & x_36336;
assign x_36338 = x_5046 & x_5047;
assign x_36339 = x_5048 & x_5049;
assign x_36340 = x_36338 & x_36339;
assign x_36341 = x_36337 & x_36340;
assign x_36342 = x_5050 & x_5051;
assign x_36343 = x_5052 & x_5053;
assign x_36344 = x_36342 & x_36343;
assign x_36345 = x_5054 & x_5055;
assign x_36346 = x_5056 & x_5057;
assign x_36347 = x_36345 & x_36346;
assign x_36348 = x_36344 & x_36347;
assign x_36349 = x_36341 & x_36348;
assign x_36350 = x_5058 & x_5059;
assign x_36351 = x_5060 & x_5061;
assign x_36352 = x_36350 & x_36351;
assign x_36353 = x_5062 & x_5063;
assign x_36354 = x_5064 & x_5065;
assign x_36355 = x_36353 & x_36354;
assign x_36356 = x_36352 & x_36355;
assign x_36357 = x_5066 & x_5067;
assign x_36358 = x_5068 & x_5069;
assign x_36359 = x_36357 & x_36358;
assign x_36360 = x_5070 & x_5071;
assign x_36361 = x_5072 & x_5073;
assign x_36362 = x_36360 & x_36361;
assign x_36363 = x_36359 & x_36362;
assign x_36364 = x_36356 & x_36363;
assign x_36365 = x_36349 & x_36364;
assign x_36366 = x_36335 & x_36365;
assign x_36367 = x_5075 & x_5076;
assign x_36368 = x_5074 & x_36367;
assign x_36369 = x_5077 & x_5078;
assign x_36370 = x_5079 & x_5080;
assign x_36371 = x_36369 & x_36370;
assign x_36372 = x_36368 & x_36371;
assign x_36373 = x_5081 & x_5082;
assign x_36374 = x_5083 & x_5084;
assign x_36375 = x_36373 & x_36374;
assign x_36376 = x_5085 & x_5086;
assign x_36377 = x_5087 & x_5088;
assign x_36378 = x_36376 & x_36377;
assign x_36379 = x_36375 & x_36378;
assign x_36380 = x_36372 & x_36379;
assign x_36381 = x_5090 & x_5091;
assign x_36382 = x_5089 & x_36381;
assign x_36383 = x_5092 & x_5093;
assign x_36384 = x_5094 & x_5095;
assign x_36385 = x_36383 & x_36384;
assign x_36386 = x_36382 & x_36385;
assign x_36387 = x_5096 & x_5097;
assign x_36388 = x_5098 & x_5099;
assign x_36389 = x_36387 & x_36388;
assign x_36390 = x_5100 & x_5101;
assign x_36391 = x_5102 & x_5103;
assign x_36392 = x_36390 & x_36391;
assign x_36393 = x_36389 & x_36392;
assign x_36394 = x_36386 & x_36393;
assign x_36395 = x_36380 & x_36394;
assign x_36396 = x_5105 & x_5106;
assign x_36397 = x_5104 & x_36396;
assign x_36398 = x_5107 & x_5108;
assign x_36399 = x_5109 & x_5110;
assign x_36400 = x_36398 & x_36399;
assign x_36401 = x_36397 & x_36400;
assign x_36402 = x_5111 & x_5112;
assign x_36403 = x_5113 & x_5114;
assign x_36404 = x_36402 & x_36403;
assign x_36405 = x_5115 & x_5116;
assign x_36406 = x_5117 & x_5118;
assign x_36407 = x_36405 & x_36406;
assign x_36408 = x_36404 & x_36407;
assign x_36409 = x_36401 & x_36408;
assign x_36410 = x_5119 & x_5120;
assign x_36411 = x_5121 & x_5122;
assign x_36412 = x_36410 & x_36411;
assign x_36413 = x_5123 & x_5124;
assign x_36414 = x_5125 & x_5126;
assign x_36415 = x_36413 & x_36414;
assign x_36416 = x_36412 & x_36415;
assign x_36417 = x_5127 & x_5128;
assign x_36418 = x_5129 & x_5130;
assign x_36419 = x_36417 & x_36418;
assign x_36420 = x_5131 & x_5132;
assign x_36421 = x_5133 & x_5134;
assign x_36422 = x_36420 & x_36421;
assign x_36423 = x_36419 & x_36422;
assign x_36424 = x_36416 & x_36423;
assign x_36425 = x_36409 & x_36424;
assign x_36426 = x_36395 & x_36425;
assign x_36427 = x_36366 & x_36426;
assign x_36428 = x_36306 & x_36427;
assign x_36429 = x_5136 & x_5137;
assign x_36430 = x_5135 & x_36429;
assign x_36431 = x_5138 & x_5139;
assign x_36432 = x_5140 & x_5141;
assign x_36433 = x_36431 & x_36432;
assign x_36434 = x_36430 & x_36433;
assign x_36435 = x_5142 & x_5143;
assign x_36436 = x_5144 & x_5145;
assign x_36437 = x_36435 & x_36436;
assign x_36438 = x_5146 & x_5147;
assign x_36439 = x_5148 & x_5149;
assign x_36440 = x_36438 & x_36439;
assign x_36441 = x_36437 & x_36440;
assign x_36442 = x_36434 & x_36441;
assign x_36443 = x_5151 & x_5152;
assign x_36444 = x_5150 & x_36443;
assign x_36445 = x_5153 & x_5154;
assign x_36446 = x_5155 & x_5156;
assign x_36447 = x_36445 & x_36446;
assign x_36448 = x_36444 & x_36447;
assign x_36449 = x_5157 & x_5158;
assign x_36450 = x_5159 & x_5160;
assign x_36451 = x_36449 & x_36450;
assign x_36452 = x_5161 & x_5162;
assign x_36453 = x_5163 & x_5164;
assign x_36454 = x_36452 & x_36453;
assign x_36455 = x_36451 & x_36454;
assign x_36456 = x_36448 & x_36455;
assign x_36457 = x_36442 & x_36456;
assign x_36458 = x_5166 & x_5167;
assign x_36459 = x_5165 & x_36458;
assign x_36460 = x_5168 & x_5169;
assign x_36461 = x_5170 & x_5171;
assign x_36462 = x_36460 & x_36461;
assign x_36463 = x_36459 & x_36462;
assign x_36464 = x_5172 & x_5173;
assign x_36465 = x_5174 & x_5175;
assign x_36466 = x_36464 & x_36465;
assign x_36467 = x_5176 & x_5177;
assign x_36468 = x_5178 & x_5179;
assign x_36469 = x_36467 & x_36468;
assign x_36470 = x_36466 & x_36469;
assign x_36471 = x_36463 & x_36470;
assign x_36472 = x_5180 & x_5181;
assign x_36473 = x_5182 & x_5183;
assign x_36474 = x_36472 & x_36473;
assign x_36475 = x_5184 & x_5185;
assign x_36476 = x_5186 & x_5187;
assign x_36477 = x_36475 & x_36476;
assign x_36478 = x_36474 & x_36477;
assign x_36479 = x_5188 & x_5189;
assign x_36480 = x_5190 & x_5191;
assign x_36481 = x_36479 & x_36480;
assign x_36482 = x_5192 & x_5193;
assign x_36483 = x_5194 & x_5195;
assign x_36484 = x_36482 & x_36483;
assign x_36485 = x_36481 & x_36484;
assign x_36486 = x_36478 & x_36485;
assign x_36487 = x_36471 & x_36486;
assign x_36488 = x_36457 & x_36487;
assign x_36489 = x_5197 & x_5198;
assign x_36490 = x_5196 & x_36489;
assign x_36491 = x_5199 & x_5200;
assign x_36492 = x_5201 & x_5202;
assign x_36493 = x_36491 & x_36492;
assign x_36494 = x_36490 & x_36493;
assign x_36495 = x_5203 & x_5204;
assign x_36496 = x_5205 & x_5206;
assign x_36497 = x_36495 & x_36496;
assign x_36498 = x_5207 & x_5208;
assign x_36499 = x_5209 & x_5210;
assign x_36500 = x_36498 & x_36499;
assign x_36501 = x_36497 & x_36500;
assign x_36502 = x_36494 & x_36501;
assign x_36503 = x_5212 & x_5213;
assign x_36504 = x_5211 & x_36503;
assign x_36505 = x_5214 & x_5215;
assign x_36506 = x_5216 & x_5217;
assign x_36507 = x_36505 & x_36506;
assign x_36508 = x_36504 & x_36507;
assign x_36509 = x_5218 & x_5219;
assign x_36510 = x_5220 & x_5221;
assign x_36511 = x_36509 & x_36510;
assign x_36512 = x_5222 & x_5223;
assign x_36513 = x_5224 & x_5225;
assign x_36514 = x_36512 & x_36513;
assign x_36515 = x_36511 & x_36514;
assign x_36516 = x_36508 & x_36515;
assign x_36517 = x_36502 & x_36516;
assign x_36518 = x_5227 & x_5228;
assign x_36519 = x_5226 & x_36518;
assign x_36520 = x_5229 & x_5230;
assign x_36521 = x_5231 & x_5232;
assign x_36522 = x_36520 & x_36521;
assign x_36523 = x_36519 & x_36522;
assign x_36524 = x_5233 & x_5234;
assign x_36525 = x_5235 & x_5236;
assign x_36526 = x_36524 & x_36525;
assign x_36527 = x_5237 & x_5238;
assign x_36528 = x_5239 & x_5240;
assign x_36529 = x_36527 & x_36528;
assign x_36530 = x_36526 & x_36529;
assign x_36531 = x_36523 & x_36530;
assign x_36532 = x_5241 & x_5242;
assign x_36533 = x_5243 & x_5244;
assign x_36534 = x_36532 & x_36533;
assign x_36535 = x_5245 & x_5246;
assign x_36536 = x_5247 & x_5248;
assign x_36537 = x_36535 & x_36536;
assign x_36538 = x_36534 & x_36537;
assign x_36539 = x_5249 & x_5250;
assign x_36540 = x_5251 & x_5252;
assign x_36541 = x_36539 & x_36540;
assign x_36542 = x_5253 & x_5254;
assign x_36543 = x_5255 & x_5256;
assign x_36544 = x_36542 & x_36543;
assign x_36545 = x_36541 & x_36544;
assign x_36546 = x_36538 & x_36545;
assign x_36547 = x_36531 & x_36546;
assign x_36548 = x_36517 & x_36547;
assign x_36549 = x_36488 & x_36548;
assign x_36550 = x_5258 & x_5259;
assign x_36551 = x_5257 & x_36550;
assign x_36552 = x_5260 & x_5261;
assign x_36553 = x_5262 & x_5263;
assign x_36554 = x_36552 & x_36553;
assign x_36555 = x_36551 & x_36554;
assign x_36556 = x_5264 & x_5265;
assign x_36557 = x_5266 & x_5267;
assign x_36558 = x_36556 & x_36557;
assign x_36559 = x_5268 & x_5269;
assign x_36560 = x_5270 & x_5271;
assign x_36561 = x_36559 & x_36560;
assign x_36562 = x_36558 & x_36561;
assign x_36563 = x_36555 & x_36562;
assign x_36564 = x_5273 & x_5274;
assign x_36565 = x_5272 & x_36564;
assign x_36566 = x_5275 & x_5276;
assign x_36567 = x_5277 & x_5278;
assign x_36568 = x_36566 & x_36567;
assign x_36569 = x_36565 & x_36568;
assign x_36570 = x_5279 & x_5280;
assign x_36571 = x_5281 & x_5282;
assign x_36572 = x_36570 & x_36571;
assign x_36573 = x_5283 & x_5284;
assign x_36574 = x_5285 & x_5286;
assign x_36575 = x_36573 & x_36574;
assign x_36576 = x_36572 & x_36575;
assign x_36577 = x_36569 & x_36576;
assign x_36578 = x_36563 & x_36577;
assign x_36579 = x_5288 & x_5289;
assign x_36580 = x_5287 & x_36579;
assign x_36581 = x_5290 & x_5291;
assign x_36582 = x_5292 & x_5293;
assign x_36583 = x_36581 & x_36582;
assign x_36584 = x_36580 & x_36583;
assign x_36585 = x_5294 & x_5295;
assign x_36586 = x_5296 & x_5297;
assign x_36587 = x_36585 & x_36586;
assign x_36588 = x_5298 & x_5299;
assign x_36589 = x_5300 & x_5301;
assign x_36590 = x_36588 & x_36589;
assign x_36591 = x_36587 & x_36590;
assign x_36592 = x_36584 & x_36591;
assign x_36593 = x_5302 & x_5303;
assign x_36594 = x_5304 & x_5305;
assign x_36595 = x_36593 & x_36594;
assign x_36596 = x_5306 & x_5307;
assign x_36597 = x_5308 & x_5309;
assign x_36598 = x_36596 & x_36597;
assign x_36599 = x_36595 & x_36598;
assign x_36600 = x_5310 & x_5311;
assign x_36601 = x_5312 & x_5313;
assign x_36602 = x_36600 & x_36601;
assign x_36603 = x_5314 & x_5315;
assign x_36604 = x_5316 & x_5317;
assign x_36605 = x_36603 & x_36604;
assign x_36606 = x_36602 & x_36605;
assign x_36607 = x_36599 & x_36606;
assign x_36608 = x_36592 & x_36607;
assign x_36609 = x_36578 & x_36608;
assign x_36610 = x_5319 & x_5320;
assign x_36611 = x_5318 & x_36610;
assign x_36612 = x_5321 & x_5322;
assign x_36613 = x_5323 & x_5324;
assign x_36614 = x_36612 & x_36613;
assign x_36615 = x_36611 & x_36614;
assign x_36616 = x_5325 & x_5326;
assign x_36617 = x_5327 & x_5328;
assign x_36618 = x_36616 & x_36617;
assign x_36619 = x_5329 & x_5330;
assign x_36620 = x_5331 & x_5332;
assign x_36621 = x_36619 & x_36620;
assign x_36622 = x_36618 & x_36621;
assign x_36623 = x_36615 & x_36622;
assign x_36624 = x_5333 & x_5334;
assign x_36625 = x_5335 & x_5336;
assign x_36626 = x_36624 & x_36625;
assign x_36627 = x_5337 & x_5338;
assign x_36628 = x_5339 & x_5340;
assign x_36629 = x_36627 & x_36628;
assign x_36630 = x_36626 & x_36629;
assign x_36631 = x_5341 & x_5342;
assign x_36632 = x_5343 & x_5344;
assign x_36633 = x_36631 & x_36632;
assign x_36634 = x_5345 & x_5346;
assign x_36635 = x_5347 & x_5348;
assign x_36636 = x_36634 & x_36635;
assign x_36637 = x_36633 & x_36636;
assign x_36638 = x_36630 & x_36637;
assign x_36639 = x_36623 & x_36638;
assign x_36640 = x_5350 & x_5351;
assign x_36641 = x_5349 & x_36640;
assign x_36642 = x_5352 & x_5353;
assign x_36643 = x_5354 & x_5355;
assign x_36644 = x_36642 & x_36643;
assign x_36645 = x_36641 & x_36644;
assign x_36646 = x_5356 & x_5357;
assign x_36647 = x_5358 & x_5359;
assign x_36648 = x_36646 & x_36647;
assign x_36649 = x_5360 & x_5361;
assign x_36650 = x_5362 & x_5363;
assign x_36651 = x_36649 & x_36650;
assign x_36652 = x_36648 & x_36651;
assign x_36653 = x_36645 & x_36652;
assign x_36654 = x_5364 & x_5365;
assign x_36655 = x_5366 & x_5367;
assign x_36656 = x_36654 & x_36655;
assign x_36657 = x_5368 & x_5369;
assign x_36658 = x_5370 & x_5371;
assign x_36659 = x_36657 & x_36658;
assign x_36660 = x_36656 & x_36659;
assign x_36661 = x_5372 & x_5373;
assign x_36662 = x_5374 & x_5375;
assign x_36663 = x_36661 & x_36662;
assign x_36664 = x_5376 & x_5377;
assign x_36665 = x_5378 & x_5379;
assign x_36666 = x_36664 & x_36665;
assign x_36667 = x_36663 & x_36666;
assign x_36668 = x_36660 & x_36667;
assign x_36669 = x_36653 & x_36668;
assign x_36670 = x_36639 & x_36669;
assign x_36671 = x_36609 & x_36670;
assign x_36672 = x_36549 & x_36671;
assign x_36673 = x_36428 & x_36672;
assign x_36674 = x_5381 & x_5382;
assign x_36675 = x_5380 & x_36674;
assign x_36676 = x_5383 & x_5384;
assign x_36677 = x_5385 & x_5386;
assign x_36678 = x_36676 & x_36677;
assign x_36679 = x_36675 & x_36678;
assign x_36680 = x_5387 & x_5388;
assign x_36681 = x_5389 & x_5390;
assign x_36682 = x_36680 & x_36681;
assign x_36683 = x_5391 & x_5392;
assign x_36684 = x_5393 & x_5394;
assign x_36685 = x_36683 & x_36684;
assign x_36686 = x_36682 & x_36685;
assign x_36687 = x_36679 & x_36686;
assign x_36688 = x_5396 & x_5397;
assign x_36689 = x_5395 & x_36688;
assign x_36690 = x_5398 & x_5399;
assign x_36691 = x_5400 & x_5401;
assign x_36692 = x_36690 & x_36691;
assign x_36693 = x_36689 & x_36692;
assign x_36694 = x_5402 & x_5403;
assign x_36695 = x_5404 & x_5405;
assign x_36696 = x_36694 & x_36695;
assign x_36697 = x_5406 & x_5407;
assign x_36698 = x_5408 & x_5409;
assign x_36699 = x_36697 & x_36698;
assign x_36700 = x_36696 & x_36699;
assign x_36701 = x_36693 & x_36700;
assign x_36702 = x_36687 & x_36701;
assign x_36703 = x_5411 & x_5412;
assign x_36704 = x_5410 & x_36703;
assign x_36705 = x_5413 & x_5414;
assign x_36706 = x_5415 & x_5416;
assign x_36707 = x_36705 & x_36706;
assign x_36708 = x_36704 & x_36707;
assign x_36709 = x_5417 & x_5418;
assign x_36710 = x_5419 & x_5420;
assign x_36711 = x_36709 & x_36710;
assign x_36712 = x_5421 & x_5422;
assign x_36713 = x_5423 & x_5424;
assign x_36714 = x_36712 & x_36713;
assign x_36715 = x_36711 & x_36714;
assign x_36716 = x_36708 & x_36715;
assign x_36717 = x_5425 & x_5426;
assign x_36718 = x_5427 & x_5428;
assign x_36719 = x_36717 & x_36718;
assign x_36720 = x_5429 & x_5430;
assign x_36721 = x_5431 & x_5432;
assign x_36722 = x_36720 & x_36721;
assign x_36723 = x_36719 & x_36722;
assign x_36724 = x_5433 & x_5434;
assign x_36725 = x_5435 & x_5436;
assign x_36726 = x_36724 & x_36725;
assign x_36727 = x_5437 & x_5438;
assign x_36728 = x_5439 & x_5440;
assign x_36729 = x_36727 & x_36728;
assign x_36730 = x_36726 & x_36729;
assign x_36731 = x_36723 & x_36730;
assign x_36732 = x_36716 & x_36731;
assign x_36733 = x_36702 & x_36732;
assign x_36734 = x_5442 & x_5443;
assign x_36735 = x_5441 & x_36734;
assign x_36736 = x_5444 & x_5445;
assign x_36737 = x_5446 & x_5447;
assign x_36738 = x_36736 & x_36737;
assign x_36739 = x_36735 & x_36738;
assign x_36740 = x_5448 & x_5449;
assign x_36741 = x_5450 & x_5451;
assign x_36742 = x_36740 & x_36741;
assign x_36743 = x_5452 & x_5453;
assign x_36744 = x_5454 & x_5455;
assign x_36745 = x_36743 & x_36744;
assign x_36746 = x_36742 & x_36745;
assign x_36747 = x_36739 & x_36746;
assign x_36748 = x_5457 & x_5458;
assign x_36749 = x_5456 & x_36748;
assign x_36750 = x_5459 & x_5460;
assign x_36751 = x_5461 & x_5462;
assign x_36752 = x_36750 & x_36751;
assign x_36753 = x_36749 & x_36752;
assign x_36754 = x_5463 & x_5464;
assign x_36755 = x_5465 & x_5466;
assign x_36756 = x_36754 & x_36755;
assign x_36757 = x_5467 & x_5468;
assign x_36758 = x_5469 & x_5470;
assign x_36759 = x_36757 & x_36758;
assign x_36760 = x_36756 & x_36759;
assign x_36761 = x_36753 & x_36760;
assign x_36762 = x_36747 & x_36761;
assign x_36763 = x_5472 & x_5473;
assign x_36764 = x_5471 & x_36763;
assign x_36765 = x_5474 & x_5475;
assign x_36766 = x_5476 & x_5477;
assign x_36767 = x_36765 & x_36766;
assign x_36768 = x_36764 & x_36767;
assign x_36769 = x_5478 & x_5479;
assign x_36770 = x_5480 & x_5481;
assign x_36771 = x_36769 & x_36770;
assign x_36772 = x_5482 & x_5483;
assign x_36773 = x_5484 & x_5485;
assign x_36774 = x_36772 & x_36773;
assign x_36775 = x_36771 & x_36774;
assign x_36776 = x_36768 & x_36775;
assign x_36777 = x_5486 & x_5487;
assign x_36778 = x_5488 & x_5489;
assign x_36779 = x_36777 & x_36778;
assign x_36780 = x_5490 & x_5491;
assign x_36781 = x_5492 & x_5493;
assign x_36782 = x_36780 & x_36781;
assign x_36783 = x_36779 & x_36782;
assign x_36784 = x_5494 & x_5495;
assign x_36785 = x_5496 & x_5497;
assign x_36786 = x_36784 & x_36785;
assign x_36787 = x_5498 & x_5499;
assign x_36788 = x_5500 & x_5501;
assign x_36789 = x_36787 & x_36788;
assign x_36790 = x_36786 & x_36789;
assign x_36791 = x_36783 & x_36790;
assign x_36792 = x_36776 & x_36791;
assign x_36793 = x_36762 & x_36792;
assign x_36794 = x_36733 & x_36793;
assign x_36795 = x_5503 & x_5504;
assign x_36796 = x_5502 & x_36795;
assign x_36797 = x_5505 & x_5506;
assign x_36798 = x_5507 & x_5508;
assign x_36799 = x_36797 & x_36798;
assign x_36800 = x_36796 & x_36799;
assign x_36801 = x_5509 & x_5510;
assign x_36802 = x_5511 & x_5512;
assign x_36803 = x_36801 & x_36802;
assign x_36804 = x_5513 & x_5514;
assign x_36805 = x_5515 & x_5516;
assign x_36806 = x_36804 & x_36805;
assign x_36807 = x_36803 & x_36806;
assign x_36808 = x_36800 & x_36807;
assign x_36809 = x_5518 & x_5519;
assign x_36810 = x_5517 & x_36809;
assign x_36811 = x_5520 & x_5521;
assign x_36812 = x_5522 & x_5523;
assign x_36813 = x_36811 & x_36812;
assign x_36814 = x_36810 & x_36813;
assign x_36815 = x_5524 & x_5525;
assign x_36816 = x_5526 & x_5527;
assign x_36817 = x_36815 & x_36816;
assign x_36818 = x_5528 & x_5529;
assign x_36819 = x_5530 & x_5531;
assign x_36820 = x_36818 & x_36819;
assign x_36821 = x_36817 & x_36820;
assign x_36822 = x_36814 & x_36821;
assign x_36823 = x_36808 & x_36822;
assign x_36824 = x_5533 & x_5534;
assign x_36825 = x_5532 & x_36824;
assign x_36826 = x_5535 & x_5536;
assign x_36827 = x_5537 & x_5538;
assign x_36828 = x_36826 & x_36827;
assign x_36829 = x_36825 & x_36828;
assign x_36830 = x_5539 & x_5540;
assign x_36831 = x_5541 & x_5542;
assign x_36832 = x_36830 & x_36831;
assign x_36833 = x_5543 & x_5544;
assign x_36834 = x_5545 & x_5546;
assign x_36835 = x_36833 & x_36834;
assign x_36836 = x_36832 & x_36835;
assign x_36837 = x_36829 & x_36836;
assign x_36838 = x_5547 & x_5548;
assign x_36839 = x_5549 & x_5550;
assign x_36840 = x_36838 & x_36839;
assign x_36841 = x_5551 & x_5552;
assign x_36842 = x_5553 & x_5554;
assign x_36843 = x_36841 & x_36842;
assign x_36844 = x_36840 & x_36843;
assign x_36845 = x_5555 & x_5556;
assign x_36846 = x_5557 & x_5558;
assign x_36847 = x_36845 & x_36846;
assign x_36848 = x_5559 & x_5560;
assign x_36849 = x_5561 & x_5562;
assign x_36850 = x_36848 & x_36849;
assign x_36851 = x_36847 & x_36850;
assign x_36852 = x_36844 & x_36851;
assign x_36853 = x_36837 & x_36852;
assign x_36854 = x_36823 & x_36853;
assign x_36855 = x_5564 & x_5565;
assign x_36856 = x_5563 & x_36855;
assign x_36857 = x_5566 & x_5567;
assign x_36858 = x_5568 & x_5569;
assign x_36859 = x_36857 & x_36858;
assign x_36860 = x_36856 & x_36859;
assign x_36861 = x_5570 & x_5571;
assign x_36862 = x_5572 & x_5573;
assign x_36863 = x_36861 & x_36862;
assign x_36864 = x_5574 & x_5575;
assign x_36865 = x_5576 & x_5577;
assign x_36866 = x_36864 & x_36865;
assign x_36867 = x_36863 & x_36866;
assign x_36868 = x_36860 & x_36867;
assign x_36869 = x_5579 & x_5580;
assign x_36870 = x_5578 & x_36869;
assign x_36871 = x_5581 & x_5582;
assign x_36872 = x_5583 & x_5584;
assign x_36873 = x_36871 & x_36872;
assign x_36874 = x_36870 & x_36873;
assign x_36875 = x_5585 & x_5586;
assign x_36876 = x_5587 & x_5588;
assign x_36877 = x_36875 & x_36876;
assign x_36878 = x_5589 & x_5590;
assign x_36879 = x_5591 & x_5592;
assign x_36880 = x_36878 & x_36879;
assign x_36881 = x_36877 & x_36880;
assign x_36882 = x_36874 & x_36881;
assign x_36883 = x_36868 & x_36882;
assign x_36884 = x_5594 & x_5595;
assign x_36885 = x_5593 & x_36884;
assign x_36886 = x_5596 & x_5597;
assign x_36887 = x_5598 & x_5599;
assign x_36888 = x_36886 & x_36887;
assign x_36889 = x_36885 & x_36888;
assign x_36890 = x_5600 & x_5601;
assign x_36891 = x_5602 & x_5603;
assign x_36892 = x_36890 & x_36891;
assign x_36893 = x_5604 & x_5605;
assign x_36894 = x_5606 & x_5607;
assign x_36895 = x_36893 & x_36894;
assign x_36896 = x_36892 & x_36895;
assign x_36897 = x_36889 & x_36896;
assign x_36898 = x_5608 & x_5609;
assign x_36899 = x_5610 & x_5611;
assign x_36900 = x_36898 & x_36899;
assign x_36901 = x_5612 & x_5613;
assign x_36902 = x_5614 & x_5615;
assign x_36903 = x_36901 & x_36902;
assign x_36904 = x_36900 & x_36903;
assign x_36905 = x_5616 & x_5617;
assign x_36906 = x_5618 & x_5619;
assign x_36907 = x_36905 & x_36906;
assign x_36908 = x_5620 & x_5621;
assign x_36909 = x_5622 & x_5623;
assign x_36910 = x_36908 & x_36909;
assign x_36911 = x_36907 & x_36910;
assign x_36912 = x_36904 & x_36911;
assign x_36913 = x_36897 & x_36912;
assign x_36914 = x_36883 & x_36913;
assign x_36915 = x_36854 & x_36914;
assign x_36916 = x_36794 & x_36915;
assign x_36917 = x_5625 & x_5626;
assign x_36918 = x_5624 & x_36917;
assign x_36919 = x_5627 & x_5628;
assign x_36920 = x_5629 & x_5630;
assign x_36921 = x_36919 & x_36920;
assign x_36922 = x_36918 & x_36921;
assign x_36923 = x_5631 & x_5632;
assign x_36924 = x_5633 & x_5634;
assign x_36925 = x_36923 & x_36924;
assign x_36926 = x_5635 & x_5636;
assign x_36927 = x_5637 & x_5638;
assign x_36928 = x_36926 & x_36927;
assign x_36929 = x_36925 & x_36928;
assign x_36930 = x_36922 & x_36929;
assign x_36931 = x_5640 & x_5641;
assign x_36932 = x_5639 & x_36931;
assign x_36933 = x_5642 & x_5643;
assign x_36934 = x_5644 & x_5645;
assign x_36935 = x_36933 & x_36934;
assign x_36936 = x_36932 & x_36935;
assign x_36937 = x_5646 & x_5647;
assign x_36938 = x_5648 & x_5649;
assign x_36939 = x_36937 & x_36938;
assign x_36940 = x_5650 & x_5651;
assign x_36941 = x_5652 & x_5653;
assign x_36942 = x_36940 & x_36941;
assign x_36943 = x_36939 & x_36942;
assign x_36944 = x_36936 & x_36943;
assign x_36945 = x_36930 & x_36944;
assign x_36946 = x_5655 & x_5656;
assign x_36947 = x_5654 & x_36946;
assign x_36948 = x_5657 & x_5658;
assign x_36949 = x_5659 & x_5660;
assign x_36950 = x_36948 & x_36949;
assign x_36951 = x_36947 & x_36950;
assign x_36952 = x_5661 & x_5662;
assign x_36953 = x_5663 & x_5664;
assign x_36954 = x_36952 & x_36953;
assign x_36955 = x_5665 & x_5666;
assign x_36956 = x_5667 & x_5668;
assign x_36957 = x_36955 & x_36956;
assign x_36958 = x_36954 & x_36957;
assign x_36959 = x_36951 & x_36958;
assign x_36960 = x_5669 & x_5670;
assign x_36961 = x_5671 & x_5672;
assign x_36962 = x_36960 & x_36961;
assign x_36963 = x_5673 & x_5674;
assign x_36964 = x_5675 & x_5676;
assign x_36965 = x_36963 & x_36964;
assign x_36966 = x_36962 & x_36965;
assign x_36967 = x_5677 & x_5678;
assign x_36968 = x_5679 & x_5680;
assign x_36969 = x_36967 & x_36968;
assign x_36970 = x_5681 & x_5682;
assign x_36971 = x_5683 & x_5684;
assign x_36972 = x_36970 & x_36971;
assign x_36973 = x_36969 & x_36972;
assign x_36974 = x_36966 & x_36973;
assign x_36975 = x_36959 & x_36974;
assign x_36976 = x_36945 & x_36975;
assign x_36977 = x_5686 & x_5687;
assign x_36978 = x_5685 & x_36977;
assign x_36979 = x_5688 & x_5689;
assign x_36980 = x_5690 & x_5691;
assign x_36981 = x_36979 & x_36980;
assign x_36982 = x_36978 & x_36981;
assign x_36983 = x_5692 & x_5693;
assign x_36984 = x_5694 & x_5695;
assign x_36985 = x_36983 & x_36984;
assign x_36986 = x_5696 & x_5697;
assign x_36987 = x_5698 & x_5699;
assign x_36988 = x_36986 & x_36987;
assign x_36989 = x_36985 & x_36988;
assign x_36990 = x_36982 & x_36989;
assign x_36991 = x_5701 & x_5702;
assign x_36992 = x_5700 & x_36991;
assign x_36993 = x_5703 & x_5704;
assign x_36994 = x_5705 & x_5706;
assign x_36995 = x_36993 & x_36994;
assign x_36996 = x_36992 & x_36995;
assign x_36997 = x_5707 & x_5708;
assign x_36998 = x_5709 & x_5710;
assign x_36999 = x_36997 & x_36998;
assign x_37000 = x_5711 & x_5712;
assign x_37001 = x_5713 & x_5714;
assign x_37002 = x_37000 & x_37001;
assign x_37003 = x_36999 & x_37002;
assign x_37004 = x_36996 & x_37003;
assign x_37005 = x_36990 & x_37004;
assign x_37006 = x_5716 & x_5717;
assign x_37007 = x_5715 & x_37006;
assign x_37008 = x_5718 & x_5719;
assign x_37009 = x_5720 & x_5721;
assign x_37010 = x_37008 & x_37009;
assign x_37011 = x_37007 & x_37010;
assign x_37012 = x_5722 & x_5723;
assign x_37013 = x_5724 & x_5725;
assign x_37014 = x_37012 & x_37013;
assign x_37015 = x_5726 & x_5727;
assign x_37016 = x_5728 & x_5729;
assign x_37017 = x_37015 & x_37016;
assign x_37018 = x_37014 & x_37017;
assign x_37019 = x_37011 & x_37018;
assign x_37020 = x_5730 & x_5731;
assign x_37021 = x_5732 & x_5733;
assign x_37022 = x_37020 & x_37021;
assign x_37023 = x_5734 & x_5735;
assign x_37024 = x_5736 & x_5737;
assign x_37025 = x_37023 & x_37024;
assign x_37026 = x_37022 & x_37025;
assign x_37027 = x_5738 & x_5739;
assign x_37028 = x_5740 & x_5741;
assign x_37029 = x_37027 & x_37028;
assign x_37030 = x_5742 & x_5743;
assign x_37031 = x_5744 & x_5745;
assign x_37032 = x_37030 & x_37031;
assign x_37033 = x_37029 & x_37032;
assign x_37034 = x_37026 & x_37033;
assign x_37035 = x_37019 & x_37034;
assign x_37036 = x_37005 & x_37035;
assign x_37037 = x_36976 & x_37036;
assign x_37038 = x_5747 & x_5748;
assign x_37039 = x_5746 & x_37038;
assign x_37040 = x_5749 & x_5750;
assign x_37041 = x_5751 & x_5752;
assign x_37042 = x_37040 & x_37041;
assign x_37043 = x_37039 & x_37042;
assign x_37044 = x_5753 & x_5754;
assign x_37045 = x_5755 & x_5756;
assign x_37046 = x_37044 & x_37045;
assign x_37047 = x_5757 & x_5758;
assign x_37048 = x_5759 & x_5760;
assign x_37049 = x_37047 & x_37048;
assign x_37050 = x_37046 & x_37049;
assign x_37051 = x_37043 & x_37050;
assign x_37052 = x_5762 & x_5763;
assign x_37053 = x_5761 & x_37052;
assign x_37054 = x_5764 & x_5765;
assign x_37055 = x_5766 & x_5767;
assign x_37056 = x_37054 & x_37055;
assign x_37057 = x_37053 & x_37056;
assign x_37058 = x_5768 & x_5769;
assign x_37059 = x_5770 & x_5771;
assign x_37060 = x_37058 & x_37059;
assign x_37061 = x_5772 & x_5773;
assign x_37062 = x_5774 & x_5775;
assign x_37063 = x_37061 & x_37062;
assign x_37064 = x_37060 & x_37063;
assign x_37065 = x_37057 & x_37064;
assign x_37066 = x_37051 & x_37065;
assign x_37067 = x_5777 & x_5778;
assign x_37068 = x_5776 & x_37067;
assign x_37069 = x_5779 & x_5780;
assign x_37070 = x_5781 & x_5782;
assign x_37071 = x_37069 & x_37070;
assign x_37072 = x_37068 & x_37071;
assign x_37073 = x_5783 & x_5784;
assign x_37074 = x_5785 & x_5786;
assign x_37075 = x_37073 & x_37074;
assign x_37076 = x_5787 & x_5788;
assign x_37077 = x_5789 & x_5790;
assign x_37078 = x_37076 & x_37077;
assign x_37079 = x_37075 & x_37078;
assign x_37080 = x_37072 & x_37079;
assign x_37081 = x_5791 & x_5792;
assign x_37082 = x_5793 & x_5794;
assign x_37083 = x_37081 & x_37082;
assign x_37084 = x_5795 & x_5796;
assign x_37085 = x_5797 & x_5798;
assign x_37086 = x_37084 & x_37085;
assign x_37087 = x_37083 & x_37086;
assign x_37088 = x_5799 & x_5800;
assign x_37089 = x_5801 & x_5802;
assign x_37090 = x_37088 & x_37089;
assign x_37091 = x_5803 & x_5804;
assign x_37092 = x_5805 & x_5806;
assign x_37093 = x_37091 & x_37092;
assign x_37094 = x_37090 & x_37093;
assign x_37095 = x_37087 & x_37094;
assign x_37096 = x_37080 & x_37095;
assign x_37097 = x_37066 & x_37096;
assign x_37098 = x_5808 & x_5809;
assign x_37099 = x_5807 & x_37098;
assign x_37100 = x_5810 & x_5811;
assign x_37101 = x_5812 & x_5813;
assign x_37102 = x_37100 & x_37101;
assign x_37103 = x_37099 & x_37102;
assign x_37104 = x_5814 & x_5815;
assign x_37105 = x_5816 & x_5817;
assign x_37106 = x_37104 & x_37105;
assign x_37107 = x_5818 & x_5819;
assign x_37108 = x_5820 & x_5821;
assign x_37109 = x_37107 & x_37108;
assign x_37110 = x_37106 & x_37109;
assign x_37111 = x_37103 & x_37110;
assign x_37112 = x_5822 & x_5823;
assign x_37113 = x_5824 & x_5825;
assign x_37114 = x_37112 & x_37113;
assign x_37115 = x_5826 & x_5827;
assign x_37116 = x_5828 & x_5829;
assign x_37117 = x_37115 & x_37116;
assign x_37118 = x_37114 & x_37117;
assign x_37119 = x_5830 & x_5831;
assign x_37120 = x_5832 & x_5833;
assign x_37121 = x_37119 & x_37120;
assign x_37122 = x_5834 & x_5835;
assign x_37123 = x_5836 & x_5837;
assign x_37124 = x_37122 & x_37123;
assign x_37125 = x_37121 & x_37124;
assign x_37126 = x_37118 & x_37125;
assign x_37127 = x_37111 & x_37126;
assign x_37128 = x_5839 & x_5840;
assign x_37129 = x_5838 & x_37128;
assign x_37130 = x_5841 & x_5842;
assign x_37131 = x_5843 & x_5844;
assign x_37132 = x_37130 & x_37131;
assign x_37133 = x_37129 & x_37132;
assign x_37134 = x_5845 & x_5846;
assign x_37135 = x_5847 & x_5848;
assign x_37136 = x_37134 & x_37135;
assign x_37137 = x_5849 & x_5850;
assign x_37138 = x_5851 & x_5852;
assign x_37139 = x_37137 & x_37138;
assign x_37140 = x_37136 & x_37139;
assign x_37141 = x_37133 & x_37140;
assign x_37142 = x_5853 & x_5854;
assign x_37143 = x_5855 & x_5856;
assign x_37144 = x_37142 & x_37143;
assign x_37145 = x_5857 & x_5858;
assign x_37146 = x_5859 & x_5860;
assign x_37147 = x_37145 & x_37146;
assign x_37148 = x_37144 & x_37147;
assign x_37149 = x_5861 & x_5862;
assign x_37150 = x_5863 & x_5864;
assign x_37151 = x_37149 & x_37150;
assign x_37152 = x_5865 & x_5866;
assign x_37153 = x_5867 & x_5868;
assign x_37154 = x_37152 & x_37153;
assign x_37155 = x_37151 & x_37154;
assign x_37156 = x_37148 & x_37155;
assign x_37157 = x_37141 & x_37156;
assign x_37158 = x_37127 & x_37157;
assign x_37159 = x_37097 & x_37158;
assign x_37160 = x_37037 & x_37159;
assign x_37161 = x_36916 & x_37160;
assign x_37162 = x_36673 & x_37161;
assign x_37163 = x_36185 & x_37162;
assign x_37164 = x_5870 & x_5871;
assign x_37165 = x_5869 & x_37164;
assign x_37166 = x_5872 & x_5873;
assign x_37167 = x_5874 & x_5875;
assign x_37168 = x_37166 & x_37167;
assign x_37169 = x_37165 & x_37168;
assign x_37170 = x_5876 & x_5877;
assign x_37171 = x_5878 & x_5879;
assign x_37172 = x_37170 & x_37171;
assign x_37173 = x_5880 & x_5881;
assign x_37174 = x_5882 & x_5883;
assign x_37175 = x_37173 & x_37174;
assign x_37176 = x_37172 & x_37175;
assign x_37177 = x_37169 & x_37176;
assign x_37178 = x_5885 & x_5886;
assign x_37179 = x_5884 & x_37178;
assign x_37180 = x_5887 & x_5888;
assign x_37181 = x_5889 & x_5890;
assign x_37182 = x_37180 & x_37181;
assign x_37183 = x_37179 & x_37182;
assign x_37184 = x_5891 & x_5892;
assign x_37185 = x_5893 & x_5894;
assign x_37186 = x_37184 & x_37185;
assign x_37187 = x_5895 & x_5896;
assign x_37188 = x_5897 & x_5898;
assign x_37189 = x_37187 & x_37188;
assign x_37190 = x_37186 & x_37189;
assign x_37191 = x_37183 & x_37190;
assign x_37192 = x_37177 & x_37191;
assign x_37193 = x_5900 & x_5901;
assign x_37194 = x_5899 & x_37193;
assign x_37195 = x_5902 & x_5903;
assign x_37196 = x_5904 & x_5905;
assign x_37197 = x_37195 & x_37196;
assign x_37198 = x_37194 & x_37197;
assign x_37199 = x_5906 & x_5907;
assign x_37200 = x_5908 & x_5909;
assign x_37201 = x_37199 & x_37200;
assign x_37202 = x_5910 & x_5911;
assign x_37203 = x_5912 & x_5913;
assign x_37204 = x_37202 & x_37203;
assign x_37205 = x_37201 & x_37204;
assign x_37206 = x_37198 & x_37205;
assign x_37207 = x_5914 & x_5915;
assign x_37208 = x_5916 & x_5917;
assign x_37209 = x_37207 & x_37208;
assign x_37210 = x_5918 & x_5919;
assign x_37211 = x_5920 & x_5921;
assign x_37212 = x_37210 & x_37211;
assign x_37213 = x_37209 & x_37212;
assign x_37214 = x_5922 & x_5923;
assign x_37215 = x_5924 & x_5925;
assign x_37216 = x_37214 & x_37215;
assign x_37217 = x_5926 & x_5927;
assign x_37218 = x_5928 & x_5929;
assign x_37219 = x_37217 & x_37218;
assign x_37220 = x_37216 & x_37219;
assign x_37221 = x_37213 & x_37220;
assign x_37222 = x_37206 & x_37221;
assign x_37223 = x_37192 & x_37222;
assign x_37224 = x_5931 & x_5932;
assign x_37225 = x_5930 & x_37224;
assign x_37226 = x_5933 & x_5934;
assign x_37227 = x_5935 & x_5936;
assign x_37228 = x_37226 & x_37227;
assign x_37229 = x_37225 & x_37228;
assign x_37230 = x_5937 & x_5938;
assign x_37231 = x_5939 & x_5940;
assign x_37232 = x_37230 & x_37231;
assign x_37233 = x_5941 & x_5942;
assign x_37234 = x_5943 & x_5944;
assign x_37235 = x_37233 & x_37234;
assign x_37236 = x_37232 & x_37235;
assign x_37237 = x_37229 & x_37236;
assign x_37238 = x_5946 & x_5947;
assign x_37239 = x_5945 & x_37238;
assign x_37240 = x_5948 & x_5949;
assign x_37241 = x_5950 & x_5951;
assign x_37242 = x_37240 & x_37241;
assign x_37243 = x_37239 & x_37242;
assign x_37244 = x_5952 & x_5953;
assign x_37245 = x_5954 & x_5955;
assign x_37246 = x_37244 & x_37245;
assign x_37247 = x_5956 & x_5957;
assign x_37248 = x_5958 & x_5959;
assign x_37249 = x_37247 & x_37248;
assign x_37250 = x_37246 & x_37249;
assign x_37251 = x_37243 & x_37250;
assign x_37252 = x_37237 & x_37251;
assign x_37253 = x_5961 & x_5962;
assign x_37254 = x_5960 & x_37253;
assign x_37255 = x_5963 & x_5964;
assign x_37256 = x_5965 & x_5966;
assign x_37257 = x_37255 & x_37256;
assign x_37258 = x_37254 & x_37257;
assign x_37259 = x_5967 & x_5968;
assign x_37260 = x_5969 & x_5970;
assign x_37261 = x_37259 & x_37260;
assign x_37262 = x_5971 & x_5972;
assign x_37263 = x_5973 & x_5974;
assign x_37264 = x_37262 & x_37263;
assign x_37265 = x_37261 & x_37264;
assign x_37266 = x_37258 & x_37265;
assign x_37267 = x_5975 & x_5976;
assign x_37268 = x_5977 & x_5978;
assign x_37269 = x_37267 & x_37268;
assign x_37270 = x_5979 & x_5980;
assign x_37271 = x_5981 & x_5982;
assign x_37272 = x_37270 & x_37271;
assign x_37273 = x_37269 & x_37272;
assign x_37274 = x_5983 & x_5984;
assign x_37275 = x_5985 & x_5986;
assign x_37276 = x_37274 & x_37275;
assign x_37277 = x_5987 & x_5988;
assign x_37278 = x_5989 & x_5990;
assign x_37279 = x_37277 & x_37278;
assign x_37280 = x_37276 & x_37279;
assign x_37281 = x_37273 & x_37280;
assign x_37282 = x_37266 & x_37281;
assign x_37283 = x_37252 & x_37282;
assign x_37284 = x_37223 & x_37283;
assign x_37285 = x_5992 & x_5993;
assign x_37286 = x_5991 & x_37285;
assign x_37287 = x_5994 & x_5995;
assign x_37288 = x_5996 & x_5997;
assign x_37289 = x_37287 & x_37288;
assign x_37290 = x_37286 & x_37289;
assign x_37291 = x_5998 & x_5999;
assign x_37292 = x_6000 & x_6001;
assign x_37293 = x_37291 & x_37292;
assign x_37294 = x_6002 & x_6003;
assign x_37295 = x_6004 & x_6005;
assign x_37296 = x_37294 & x_37295;
assign x_37297 = x_37293 & x_37296;
assign x_37298 = x_37290 & x_37297;
assign x_37299 = x_6007 & x_6008;
assign x_37300 = x_6006 & x_37299;
assign x_37301 = x_6009 & x_6010;
assign x_37302 = x_6011 & x_6012;
assign x_37303 = x_37301 & x_37302;
assign x_37304 = x_37300 & x_37303;
assign x_37305 = x_6013 & x_6014;
assign x_37306 = x_6015 & x_6016;
assign x_37307 = x_37305 & x_37306;
assign x_37308 = x_6017 & x_6018;
assign x_37309 = x_6019 & x_6020;
assign x_37310 = x_37308 & x_37309;
assign x_37311 = x_37307 & x_37310;
assign x_37312 = x_37304 & x_37311;
assign x_37313 = x_37298 & x_37312;
assign x_37314 = x_6022 & x_6023;
assign x_37315 = x_6021 & x_37314;
assign x_37316 = x_6024 & x_6025;
assign x_37317 = x_6026 & x_6027;
assign x_37318 = x_37316 & x_37317;
assign x_37319 = x_37315 & x_37318;
assign x_37320 = x_6028 & x_6029;
assign x_37321 = x_6030 & x_6031;
assign x_37322 = x_37320 & x_37321;
assign x_37323 = x_6032 & x_6033;
assign x_37324 = x_6034 & x_6035;
assign x_37325 = x_37323 & x_37324;
assign x_37326 = x_37322 & x_37325;
assign x_37327 = x_37319 & x_37326;
assign x_37328 = x_6036 & x_6037;
assign x_37329 = x_6038 & x_6039;
assign x_37330 = x_37328 & x_37329;
assign x_37331 = x_6040 & x_6041;
assign x_37332 = x_6042 & x_6043;
assign x_37333 = x_37331 & x_37332;
assign x_37334 = x_37330 & x_37333;
assign x_37335 = x_6044 & x_6045;
assign x_37336 = x_6046 & x_6047;
assign x_37337 = x_37335 & x_37336;
assign x_37338 = x_6048 & x_6049;
assign x_37339 = x_6050 & x_6051;
assign x_37340 = x_37338 & x_37339;
assign x_37341 = x_37337 & x_37340;
assign x_37342 = x_37334 & x_37341;
assign x_37343 = x_37327 & x_37342;
assign x_37344 = x_37313 & x_37343;
assign x_37345 = x_6053 & x_6054;
assign x_37346 = x_6052 & x_37345;
assign x_37347 = x_6055 & x_6056;
assign x_37348 = x_6057 & x_6058;
assign x_37349 = x_37347 & x_37348;
assign x_37350 = x_37346 & x_37349;
assign x_37351 = x_6059 & x_6060;
assign x_37352 = x_6061 & x_6062;
assign x_37353 = x_37351 & x_37352;
assign x_37354 = x_6063 & x_6064;
assign x_37355 = x_6065 & x_6066;
assign x_37356 = x_37354 & x_37355;
assign x_37357 = x_37353 & x_37356;
assign x_37358 = x_37350 & x_37357;
assign x_37359 = x_6068 & x_6069;
assign x_37360 = x_6067 & x_37359;
assign x_37361 = x_6070 & x_6071;
assign x_37362 = x_6072 & x_6073;
assign x_37363 = x_37361 & x_37362;
assign x_37364 = x_37360 & x_37363;
assign x_37365 = x_6074 & x_6075;
assign x_37366 = x_6076 & x_6077;
assign x_37367 = x_37365 & x_37366;
assign x_37368 = x_6078 & x_6079;
assign x_37369 = x_6080 & x_6081;
assign x_37370 = x_37368 & x_37369;
assign x_37371 = x_37367 & x_37370;
assign x_37372 = x_37364 & x_37371;
assign x_37373 = x_37358 & x_37372;
assign x_37374 = x_6083 & x_6084;
assign x_37375 = x_6082 & x_37374;
assign x_37376 = x_6085 & x_6086;
assign x_37377 = x_6087 & x_6088;
assign x_37378 = x_37376 & x_37377;
assign x_37379 = x_37375 & x_37378;
assign x_37380 = x_6089 & x_6090;
assign x_37381 = x_6091 & x_6092;
assign x_37382 = x_37380 & x_37381;
assign x_37383 = x_6093 & x_6094;
assign x_37384 = x_6095 & x_6096;
assign x_37385 = x_37383 & x_37384;
assign x_37386 = x_37382 & x_37385;
assign x_37387 = x_37379 & x_37386;
assign x_37388 = x_6097 & x_6098;
assign x_37389 = x_6099 & x_6100;
assign x_37390 = x_37388 & x_37389;
assign x_37391 = x_6101 & x_6102;
assign x_37392 = x_6103 & x_6104;
assign x_37393 = x_37391 & x_37392;
assign x_37394 = x_37390 & x_37393;
assign x_37395 = x_6105 & x_6106;
assign x_37396 = x_6107 & x_6108;
assign x_37397 = x_37395 & x_37396;
assign x_37398 = x_6109 & x_6110;
assign x_37399 = x_6111 & x_6112;
assign x_37400 = x_37398 & x_37399;
assign x_37401 = x_37397 & x_37400;
assign x_37402 = x_37394 & x_37401;
assign x_37403 = x_37387 & x_37402;
assign x_37404 = x_37373 & x_37403;
assign x_37405 = x_37344 & x_37404;
assign x_37406 = x_37284 & x_37405;
assign x_37407 = x_6114 & x_6115;
assign x_37408 = x_6113 & x_37407;
assign x_37409 = x_6116 & x_6117;
assign x_37410 = x_6118 & x_6119;
assign x_37411 = x_37409 & x_37410;
assign x_37412 = x_37408 & x_37411;
assign x_37413 = x_6120 & x_6121;
assign x_37414 = x_6122 & x_6123;
assign x_37415 = x_37413 & x_37414;
assign x_37416 = x_6124 & x_6125;
assign x_37417 = x_6126 & x_6127;
assign x_37418 = x_37416 & x_37417;
assign x_37419 = x_37415 & x_37418;
assign x_37420 = x_37412 & x_37419;
assign x_37421 = x_6129 & x_6130;
assign x_37422 = x_6128 & x_37421;
assign x_37423 = x_6131 & x_6132;
assign x_37424 = x_6133 & x_6134;
assign x_37425 = x_37423 & x_37424;
assign x_37426 = x_37422 & x_37425;
assign x_37427 = x_6135 & x_6136;
assign x_37428 = x_6137 & x_6138;
assign x_37429 = x_37427 & x_37428;
assign x_37430 = x_6139 & x_6140;
assign x_37431 = x_6141 & x_6142;
assign x_37432 = x_37430 & x_37431;
assign x_37433 = x_37429 & x_37432;
assign x_37434 = x_37426 & x_37433;
assign x_37435 = x_37420 & x_37434;
assign x_37436 = x_6144 & x_6145;
assign x_37437 = x_6143 & x_37436;
assign x_37438 = x_6146 & x_6147;
assign x_37439 = x_6148 & x_6149;
assign x_37440 = x_37438 & x_37439;
assign x_37441 = x_37437 & x_37440;
assign x_37442 = x_6150 & x_6151;
assign x_37443 = x_6152 & x_6153;
assign x_37444 = x_37442 & x_37443;
assign x_37445 = x_6154 & x_6155;
assign x_37446 = x_6156 & x_6157;
assign x_37447 = x_37445 & x_37446;
assign x_37448 = x_37444 & x_37447;
assign x_37449 = x_37441 & x_37448;
assign x_37450 = x_6158 & x_6159;
assign x_37451 = x_6160 & x_6161;
assign x_37452 = x_37450 & x_37451;
assign x_37453 = x_6162 & x_6163;
assign x_37454 = x_6164 & x_6165;
assign x_37455 = x_37453 & x_37454;
assign x_37456 = x_37452 & x_37455;
assign x_37457 = x_6166 & x_6167;
assign x_37458 = x_6168 & x_6169;
assign x_37459 = x_37457 & x_37458;
assign x_37460 = x_6170 & x_6171;
assign x_37461 = x_6172 & x_6173;
assign x_37462 = x_37460 & x_37461;
assign x_37463 = x_37459 & x_37462;
assign x_37464 = x_37456 & x_37463;
assign x_37465 = x_37449 & x_37464;
assign x_37466 = x_37435 & x_37465;
assign x_37467 = x_6175 & x_6176;
assign x_37468 = x_6174 & x_37467;
assign x_37469 = x_6177 & x_6178;
assign x_37470 = x_6179 & x_6180;
assign x_37471 = x_37469 & x_37470;
assign x_37472 = x_37468 & x_37471;
assign x_37473 = x_6181 & x_6182;
assign x_37474 = x_6183 & x_6184;
assign x_37475 = x_37473 & x_37474;
assign x_37476 = x_6185 & x_6186;
assign x_37477 = x_6187 & x_6188;
assign x_37478 = x_37476 & x_37477;
assign x_37479 = x_37475 & x_37478;
assign x_37480 = x_37472 & x_37479;
assign x_37481 = x_6190 & x_6191;
assign x_37482 = x_6189 & x_37481;
assign x_37483 = x_6192 & x_6193;
assign x_37484 = x_6194 & x_6195;
assign x_37485 = x_37483 & x_37484;
assign x_37486 = x_37482 & x_37485;
assign x_37487 = x_6196 & x_6197;
assign x_37488 = x_6198 & x_6199;
assign x_37489 = x_37487 & x_37488;
assign x_37490 = x_6200 & x_6201;
assign x_37491 = x_6202 & x_6203;
assign x_37492 = x_37490 & x_37491;
assign x_37493 = x_37489 & x_37492;
assign x_37494 = x_37486 & x_37493;
assign x_37495 = x_37480 & x_37494;
assign x_37496 = x_6205 & x_6206;
assign x_37497 = x_6204 & x_37496;
assign x_37498 = x_6207 & x_6208;
assign x_37499 = x_6209 & x_6210;
assign x_37500 = x_37498 & x_37499;
assign x_37501 = x_37497 & x_37500;
assign x_37502 = x_6211 & x_6212;
assign x_37503 = x_6213 & x_6214;
assign x_37504 = x_37502 & x_37503;
assign x_37505 = x_6215 & x_6216;
assign x_37506 = x_6217 & x_6218;
assign x_37507 = x_37505 & x_37506;
assign x_37508 = x_37504 & x_37507;
assign x_37509 = x_37501 & x_37508;
assign x_37510 = x_6219 & x_6220;
assign x_37511 = x_6221 & x_6222;
assign x_37512 = x_37510 & x_37511;
assign x_37513 = x_6223 & x_6224;
assign x_37514 = x_6225 & x_6226;
assign x_37515 = x_37513 & x_37514;
assign x_37516 = x_37512 & x_37515;
assign x_37517 = x_6227 & x_6228;
assign x_37518 = x_6229 & x_6230;
assign x_37519 = x_37517 & x_37518;
assign x_37520 = x_6231 & x_6232;
assign x_37521 = x_6233 & x_6234;
assign x_37522 = x_37520 & x_37521;
assign x_37523 = x_37519 & x_37522;
assign x_37524 = x_37516 & x_37523;
assign x_37525 = x_37509 & x_37524;
assign x_37526 = x_37495 & x_37525;
assign x_37527 = x_37466 & x_37526;
assign x_37528 = x_6236 & x_6237;
assign x_37529 = x_6235 & x_37528;
assign x_37530 = x_6238 & x_6239;
assign x_37531 = x_6240 & x_6241;
assign x_37532 = x_37530 & x_37531;
assign x_37533 = x_37529 & x_37532;
assign x_37534 = x_6242 & x_6243;
assign x_37535 = x_6244 & x_6245;
assign x_37536 = x_37534 & x_37535;
assign x_37537 = x_6246 & x_6247;
assign x_37538 = x_6248 & x_6249;
assign x_37539 = x_37537 & x_37538;
assign x_37540 = x_37536 & x_37539;
assign x_37541 = x_37533 & x_37540;
assign x_37542 = x_6251 & x_6252;
assign x_37543 = x_6250 & x_37542;
assign x_37544 = x_6253 & x_6254;
assign x_37545 = x_6255 & x_6256;
assign x_37546 = x_37544 & x_37545;
assign x_37547 = x_37543 & x_37546;
assign x_37548 = x_6257 & x_6258;
assign x_37549 = x_6259 & x_6260;
assign x_37550 = x_37548 & x_37549;
assign x_37551 = x_6261 & x_6262;
assign x_37552 = x_6263 & x_6264;
assign x_37553 = x_37551 & x_37552;
assign x_37554 = x_37550 & x_37553;
assign x_37555 = x_37547 & x_37554;
assign x_37556 = x_37541 & x_37555;
assign x_37557 = x_6266 & x_6267;
assign x_37558 = x_6265 & x_37557;
assign x_37559 = x_6268 & x_6269;
assign x_37560 = x_6270 & x_6271;
assign x_37561 = x_37559 & x_37560;
assign x_37562 = x_37558 & x_37561;
assign x_37563 = x_6272 & x_6273;
assign x_37564 = x_6274 & x_6275;
assign x_37565 = x_37563 & x_37564;
assign x_37566 = x_6276 & x_6277;
assign x_37567 = x_6278 & x_6279;
assign x_37568 = x_37566 & x_37567;
assign x_37569 = x_37565 & x_37568;
assign x_37570 = x_37562 & x_37569;
assign x_37571 = x_6280 & x_6281;
assign x_37572 = x_6282 & x_6283;
assign x_37573 = x_37571 & x_37572;
assign x_37574 = x_6284 & x_6285;
assign x_37575 = x_6286 & x_6287;
assign x_37576 = x_37574 & x_37575;
assign x_37577 = x_37573 & x_37576;
assign x_37578 = x_6288 & x_6289;
assign x_37579 = x_6290 & x_6291;
assign x_37580 = x_37578 & x_37579;
assign x_37581 = x_6292 & x_6293;
assign x_37582 = x_6294 & x_6295;
assign x_37583 = x_37581 & x_37582;
assign x_37584 = x_37580 & x_37583;
assign x_37585 = x_37577 & x_37584;
assign x_37586 = x_37570 & x_37585;
assign x_37587 = x_37556 & x_37586;
assign x_37588 = x_6297 & x_6298;
assign x_37589 = x_6296 & x_37588;
assign x_37590 = x_6299 & x_6300;
assign x_37591 = x_6301 & x_6302;
assign x_37592 = x_37590 & x_37591;
assign x_37593 = x_37589 & x_37592;
assign x_37594 = x_6303 & x_6304;
assign x_37595 = x_6305 & x_6306;
assign x_37596 = x_37594 & x_37595;
assign x_37597 = x_6307 & x_6308;
assign x_37598 = x_6309 & x_6310;
assign x_37599 = x_37597 & x_37598;
assign x_37600 = x_37596 & x_37599;
assign x_37601 = x_37593 & x_37600;
assign x_37602 = x_6311 & x_6312;
assign x_37603 = x_6313 & x_6314;
assign x_37604 = x_37602 & x_37603;
assign x_37605 = x_6315 & x_6316;
assign x_37606 = x_6317 & x_6318;
assign x_37607 = x_37605 & x_37606;
assign x_37608 = x_37604 & x_37607;
assign x_37609 = x_6319 & x_6320;
assign x_37610 = x_6321 & x_6322;
assign x_37611 = x_37609 & x_37610;
assign x_37612 = x_6323 & x_6324;
assign x_37613 = x_6325 & x_6326;
assign x_37614 = x_37612 & x_37613;
assign x_37615 = x_37611 & x_37614;
assign x_37616 = x_37608 & x_37615;
assign x_37617 = x_37601 & x_37616;
assign x_37618 = x_6328 & x_6329;
assign x_37619 = x_6327 & x_37618;
assign x_37620 = x_6330 & x_6331;
assign x_37621 = x_6332 & x_6333;
assign x_37622 = x_37620 & x_37621;
assign x_37623 = x_37619 & x_37622;
assign x_37624 = x_6334 & x_6335;
assign x_37625 = x_6336 & x_6337;
assign x_37626 = x_37624 & x_37625;
assign x_37627 = x_6338 & x_6339;
assign x_37628 = x_6340 & x_6341;
assign x_37629 = x_37627 & x_37628;
assign x_37630 = x_37626 & x_37629;
assign x_37631 = x_37623 & x_37630;
assign x_37632 = x_6342 & x_6343;
assign x_37633 = x_6344 & x_6345;
assign x_37634 = x_37632 & x_37633;
assign x_37635 = x_6346 & x_6347;
assign x_37636 = x_6348 & x_6349;
assign x_37637 = x_37635 & x_37636;
assign x_37638 = x_37634 & x_37637;
assign x_37639 = x_6350 & x_6351;
assign x_37640 = x_6352 & x_6353;
assign x_37641 = x_37639 & x_37640;
assign x_37642 = x_6354 & x_6355;
assign x_37643 = x_6356 & x_6357;
assign x_37644 = x_37642 & x_37643;
assign x_37645 = x_37641 & x_37644;
assign x_37646 = x_37638 & x_37645;
assign x_37647 = x_37631 & x_37646;
assign x_37648 = x_37617 & x_37647;
assign x_37649 = x_37587 & x_37648;
assign x_37650 = x_37527 & x_37649;
assign x_37651 = x_37406 & x_37650;
assign x_37652 = x_6359 & x_6360;
assign x_37653 = x_6358 & x_37652;
assign x_37654 = x_6361 & x_6362;
assign x_37655 = x_6363 & x_6364;
assign x_37656 = x_37654 & x_37655;
assign x_37657 = x_37653 & x_37656;
assign x_37658 = x_6365 & x_6366;
assign x_37659 = x_6367 & x_6368;
assign x_37660 = x_37658 & x_37659;
assign x_37661 = x_6369 & x_6370;
assign x_37662 = x_6371 & x_6372;
assign x_37663 = x_37661 & x_37662;
assign x_37664 = x_37660 & x_37663;
assign x_37665 = x_37657 & x_37664;
assign x_37666 = x_6374 & x_6375;
assign x_37667 = x_6373 & x_37666;
assign x_37668 = x_6376 & x_6377;
assign x_37669 = x_6378 & x_6379;
assign x_37670 = x_37668 & x_37669;
assign x_37671 = x_37667 & x_37670;
assign x_37672 = x_6380 & x_6381;
assign x_37673 = x_6382 & x_6383;
assign x_37674 = x_37672 & x_37673;
assign x_37675 = x_6384 & x_6385;
assign x_37676 = x_6386 & x_6387;
assign x_37677 = x_37675 & x_37676;
assign x_37678 = x_37674 & x_37677;
assign x_37679 = x_37671 & x_37678;
assign x_37680 = x_37665 & x_37679;
assign x_37681 = x_6389 & x_6390;
assign x_37682 = x_6388 & x_37681;
assign x_37683 = x_6391 & x_6392;
assign x_37684 = x_6393 & x_6394;
assign x_37685 = x_37683 & x_37684;
assign x_37686 = x_37682 & x_37685;
assign x_37687 = x_6395 & x_6396;
assign x_37688 = x_6397 & x_6398;
assign x_37689 = x_37687 & x_37688;
assign x_37690 = x_6399 & x_6400;
assign x_37691 = x_6401 & x_6402;
assign x_37692 = x_37690 & x_37691;
assign x_37693 = x_37689 & x_37692;
assign x_37694 = x_37686 & x_37693;
assign x_37695 = x_6403 & x_6404;
assign x_37696 = x_6405 & x_6406;
assign x_37697 = x_37695 & x_37696;
assign x_37698 = x_6407 & x_6408;
assign x_37699 = x_6409 & x_6410;
assign x_37700 = x_37698 & x_37699;
assign x_37701 = x_37697 & x_37700;
assign x_37702 = x_6411 & x_6412;
assign x_37703 = x_6413 & x_6414;
assign x_37704 = x_37702 & x_37703;
assign x_37705 = x_6415 & x_6416;
assign x_37706 = x_6417 & x_6418;
assign x_37707 = x_37705 & x_37706;
assign x_37708 = x_37704 & x_37707;
assign x_37709 = x_37701 & x_37708;
assign x_37710 = x_37694 & x_37709;
assign x_37711 = x_37680 & x_37710;
assign x_37712 = x_6420 & x_6421;
assign x_37713 = x_6419 & x_37712;
assign x_37714 = x_6422 & x_6423;
assign x_37715 = x_6424 & x_6425;
assign x_37716 = x_37714 & x_37715;
assign x_37717 = x_37713 & x_37716;
assign x_37718 = x_6426 & x_6427;
assign x_37719 = x_6428 & x_6429;
assign x_37720 = x_37718 & x_37719;
assign x_37721 = x_6430 & x_6431;
assign x_37722 = x_6432 & x_6433;
assign x_37723 = x_37721 & x_37722;
assign x_37724 = x_37720 & x_37723;
assign x_37725 = x_37717 & x_37724;
assign x_37726 = x_6435 & x_6436;
assign x_37727 = x_6434 & x_37726;
assign x_37728 = x_6437 & x_6438;
assign x_37729 = x_6439 & x_6440;
assign x_37730 = x_37728 & x_37729;
assign x_37731 = x_37727 & x_37730;
assign x_37732 = x_6441 & x_6442;
assign x_37733 = x_6443 & x_6444;
assign x_37734 = x_37732 & x_37733;
assign x_37735 = x_6445 & x_6446;
assign x_37736 = x_6447 & x_6448;
assign x_37737 = x_37735 & x_37736;
assign x_37738 = x_37734 & x_37737;
assign x_37739 = x_37731 & x_37738;
assign x_37740 = x_37725 & x_37739;
assign x_37741 = x_6450 & x_6451;
assign x_37742 = x_6449 & x_37741;
assign x_37743 = x_6452 & x_6453;
assign x_37744 = x_6454 & x_6455;
assign x_37745 = x_37743 & x_37744;
assign x_37746 = x_37742 & x_37745;
assign x_37747 = x_6456 & x_6457;
assign x_37748 = x_6458 & x_6459;
assign x_37749 = x_37747 & x_37748;
assign x_37750 = x_6460 & x_6461;
assign x_37751 = x_6462 & x_6463;
assign x_37752 = x_37750 & x_37751;
assign x_37753 = x_37749 & x_37752;
assign x_37754 = x_37746 & x_37753;
assign x_37755 = x_6464 & x_6465;
assign x_37756 = x_6466 & x_6467;
assign x_37757 = x_37755 & x_37756;
assign x_37758 = x_6468 & x_6469;
assign x_37759 = x_6470 & x_6471;
assign x_37760 = x_37758 & x_37759;
assign x_37761 = x_37757 & x_37760;
assign x_37762 = x_6472 & x_6473;
assign x_37763 = x_6474 & x_6475;
assign x_37764 = x_37762 & x_37763;
assign x_37765 = x_6476 & x_6477;
assign x_37766 = x_6478 & x_6479;
assign x_37767 = x_37765 & x_37766;
assign x_37768 = x_37764 & x_37767;
assign x_37769 = x_37761 & x_37768;
assign x_37770 = x_37754 & x_37769;
assign x_37771 = x_37740 & x_37770;
assign x_37772 = x_37711 & x_37771;
assign x_37773 = x_6481 & x_6482;
assign x_37774 = x_6480 & x_37773;
assign x_37775 = x_6483 & x_6484;
assign x_37776 = x_6485 & x_6486;
assign x_37777 = x_37775 & x_37776;
assign x_37778 = x_37774 & x_37777;
assign x_37779 = x_6487 & x_6488;
assign x_37780 = x_6489 & x_6490;
assign x_37781 = x_37779 & x_37780;
assign x_37782 = x_6491 & x_6492;
assign x_37783 = x_6493 & x_6494;
assign x_37784 = x_37782 & x_37783;
assign x_37785 = x_37781 & x_37784;
assign x_37786 = x_37778 & x_37785;
assign x_37787 = x_6496 & x_6497;
assign x_37788 = x_6495 & x_37787;
assign x_37789 = x_6498 & x_6499;
assign x_37790 = x_6500 & x_6501;
assign x_37791 = x_37789 & x_37790;
assign x_37792 = x_37788 & x_37791;
assign x_37793 = x_6502 & x_6503;
assign x_37794 = x_6504 & x_6505;
assign x_37795 = x_37793 & x_37794;
assign x_37796 = x_6506 & x_6507;
assign x_37797 = x_6508 & x_6509;
assign x_37798 = x_37796 & x_37797;
assign x_37799 = x_37795 & x_37798;
assign x_37800 = x_37792 & x_37799;
assign x_37801 = x_37786 & x_37800;
assign x_37802 = x_6511 & x_6512;
assign x_37803 = x_6510 & x_37802;
assign x_37804 = x_6513 & x_6514;
assign x_37805 = x_6515 & x_6516;
assign x_37806 = x_37804 & x_37805;
assign x_37807 = x_37803 & x_37806;
assign x_37808 = x_6517 & x_6518;
assign x_37809 = x_6519 & x_6520;
assign x_37810 = x_37808 & x_37809;
assign x_37811 = x_6521 & x_6522;
assign x_37812 = x_6523 & x_6524;
assign x_37813 = x_37811 & x_37812;
assign x_37814 = x_37810 & x_37813;
assign x_37815 = x_37807 & x_37814;
assign x_37816 = x_6525 & x_6526;
assign x_37817 = x_6527 & x_6528;
assign x_37818 = x_37816 & x_37817;
assign x_37819 = x_6529 & x_6530;
assign x_37820 = x_6531 & x_6532;
assign x_37821 = x_37819 & x_37820;
assign x_37822 = x_37818 & x_37821;
assign x_37823 = x_6533 & x_6534;
assign x_37824 = x_6535 & x_6536;
assign x_37825 = x_37823 & x_37824;
assign x_37826 = x_6537 & x_6538;
assign x_37827 = x_6539 & x_6540;
assign x_37828 = x_37826 & x_37827;
assign x_37829 = x_37825 & x_37828;
assign x_37830 = x_37822 & x_37829;
assign x_37831 = x_37815 & x_37830;
assign x_37832 = x_37801 & x_37831;
assign x_37833 = x_6542 & x_6543;
assign x_37834 = x_6541 & x_37833;
assign x_37835 = x_6544 & x_6545;
assign x_37836 = x_6546 & x_6547;
assign x_37837 = x_37835 & x_37836;
assign x_37838 = x_37834 & x_37837;
assign x_37839 = x_6548 & x_6549;
assign x_37840 = x_6550 & x_6551;
assign x_37841 = x_37839 & x_37840;
assign x_37842 = x_6552 & x_6553;
assign x_37843 = x_6554 & x_6555;
assign x_37844 = x_37842 & x_37843;
assign x_37845 = x_37841 & x_37844;
assign x_37846 = x_37838 & x_37845;
assign x_37847 = x_6557 & x_6558;
assign x_37848 = x_6556 & x_37847;
assign x_37849 = x_6559 & x_6560;
assign x_37850 = x_6561 & x_6562;
assign x_37851 = x_37849 & x_37850;
assign x_37852 = x_37848 & x_37851;
assign x_37853 = x_6563 & x_6564;
assign x_37854 = x_6565 & x_6566;
assign x_37855 = x_37853 & x_37854;
assign x_37856 = x_6567 & x_6568;
assign x_37857 = x_6569 & x_6570;
assign x_37858 = x_37856 & x_37857;
assign x_37859 = x_37855 & x_37858;
assign x_37860 = x_37852 & x_37859;
assign x_37861 = x_37846 & x_37860;
assign x_37862 = x_6572 & x_6573;
assign x_37863 = x_6571 & x_37862;
assign x_37864 = x_6574 & x_6575;
assign x_37865 = x_6576 & x_6577;
assign x_37866 = x_37864 & x_37865;
assign x_37867 = x_37863 & x_37866;
assign x_37868 = x_6578 & x_6579;
assign x_37869 = x_6580 & x_6581;
assign x_37870 = x_37868 & x_37869;
assign x_37871 = x_6582 & x_6583;
assign x_37872 = x_6584 & x_6585;
assign x_37873 = x_37871 & x_37872;
assign x_37874 = x_37870 & x_37873;
assign x_37875 = x_37867 & x_37874;
assign x_37876 = x_6586 & x_6587;
assign x_37877 = x_6588 & x_6589;
assign x_37878 = x_37876 & x_37877;
assign x_37879 = x_6590 & x_6591;
assign x_37880 = x_6592 & x_6593;
assign x_37881 = x_37879 & x_37880;
assign x_37882 = x_37878 & x_37881;
assign x_37883 = x_6594 & x_6595;
assign x_37884 = x_6596 & x_6597;
assign x_37885 = x_37883 & x_37884;
assign x_37886 = x_6598 & x_6599;
assign x_37887 = x_6600 & x_6601;
assign x_37888 = x_37886 & x_37887;
assign x_37889 = x_37885 & x_37888;
assign x_37890 = x_37882 & x_37889;
assign x_37891 = x_37875 & x_37890;
assign x_37892 = x_37861 & x_37891;
assign x_37893 = x_37832 & x_37892;
assign x_37894 = x_37772 & x_37893;
assign x_37895 = x_6603 & x_6604;
assign x_37896 = x_6602 & x_37895;
assign x_37897 = x_6605 & x_6606;
assign x_37898 = x_6607 & x_6608;
assign x_37899 = x_37897 & x_37898;
assign x_37900 = x_37896 & x_37899;
assign x_37901 = x_6609 & x_6610;
assign x_37902 = x_6611 & x_6612;
assign x_37903 = x_37901 & x_37902;
assign x_37904 = x_6613 & x_6614;
assign x_37905 = x_6615 & x_6616;
assign x_37906 = x_37904 & x_37905;
assign x_37907 = x_37903 & x_37906;
assign x_37908 = x_37900 & x_37907;
assign x_37909 = x_6618 & x_6619;
assign x_37910 = x_6617 & x_37909;
assign x_37911 = x_6620 & x_6621;
assign x_37912 = x_6622 & x_6623;
assign x_37913 = x_37911 & x_37912;
assign x_37914 = x_37910 & x_37913;
assign x_37915 = x_6624 & x_6625;
assign x_37916 = x_6626 & x_6627;
assign x_37917 = x_37915 & x_37916;
assign x_37918 = x_6628 & x_6629;
assign x_37919 = x_6630 & x_6631;
assign x_37920 = x_37918 & x_37919;
assign x_37921 = x_37917 & x_37920;
assign x_37922 = x_37914 & x_37921;
assign x_37923 = x_37908 & x_37922;
assign x_37924 = x_6633 & x_6634;
assign x_37925 = x_6632 & x_37924;
assign x_37926 = x_6635 & x_6636;
assign x_37927 = x_6637 & x_6638;
assign x_37928 = x_37926 & x_37927;
assign x_37929 = x_37925 & x_37928;
assign x_37930 = x_6639 & x_6640;
assign x_37931 = x_6641 & x_6642;
assign x_37932 = x_37930 & x_37931;
assign x_37933 = x_6643 & x_6644;
assign x_37934 = x_6645 & x_6646;
assign x_37935 = x_37933 & x_37934;
assign x_37936 = x_37932 & x_37935;
assign x_37937 = x_37929 & x_37936;
assign x_37938 = x_6647 & x_6648;
assign x_37939 = x_6649 & x_6650;
assign x_37940 = x_37938 & x_37939;
assign x_37941 = x_6651 & x_6652;
assign x_37942 = x_6653 & x_6654;
assign x_37943 = x_37941 & x_37942;
assign x_37944 = x_37940 & x_37943;
assign x_37945 = x_6655 & x_6656;
assign x_37946 = x_6657 & x_6658;
assign x_37947 = x_37945 & x_37946;
assign x_37948 = x_6659 & x_6660;
assign x_37949 = x_6661 & x_6662;
assign x_37950 = x_37948 & x_37949;
assign x_37951 = x_37947 & x_37950;
assign x_37952 = x_37944 & x_37951;
assign x_37953 = x_37937 & x_37952;
assign x_37954 = x_37923 & x_37953;
assign x_37955 = x_6664 & x_6665;
assign x_37956 = x_6663 & x_37955;
assign x_37957 = x_6666 & x_6667;
assign x_37958 = x_6668 & x_6669;
assign x_37959 = x_37957 & x_37958;
assign x_37960 = x_37956 & x_37959;
assign x_37961 = x_6670 & x_6671;
assign x_37962 = x_6672 & x_6673;
assign x_37963 = x_37961 & x_37962;
assign x_37964 = x_6674 & x_6675;
assign x_37965 = x_6676 & x_6677;
assign x_37966 = x_37964 & x_37965;
assign x_37967 = x_37963 & x_37966;
assign x_37968 = x_37960 & x_37967;
assign x_37969 = x_6679 & x_6680;
assign x_37970 = x_6678 & x_37969;
assign x_37971 = x_6681 & x_6682;
assign x_37972 = x_6683 & x_6684;
assign x_37973 = x_37971 & x_37972;
assign x_37974 = x_37970 & x_37973;
assign x_37975 = x_6685 & x_6686;
assign x_37976 = x_6687 & x_6688;
assign x_37977 = x_37975 & x_37976;
assign x_37978 = x_6689 & x_6690;
assign x_37979 = x_6691 & x_6692;
assign x_37980 = x_37978 & x_37979;
assign x_37981 = x_37977 & x_37980;
assign x_37982 = x_37974 & x_37981;
assign x_37983 = x_37968 & x_37982;
assign x_37984 = x_6694 & x_6695;
assign x_37985 = x_6693 & x_37984;
assign x_37986 = x_6696 & x_6697;
assign x_37987 = x_6698 & x_6699;
assign x_37988 = x_37986 & x_37987;
assign x_37989 = x_37985 & x_37988;
assign x_37990 = x_6700 & x_6701;
assign x_37991 = x_6702 & x_6703;
assign x_37992 = x_37990 & x_37991;
assign x_37993 = x_6704 & x_6705;
assign x_37994 = x_6706 & x_6707;
assign x_37995 = x_37993 & x_37994;
assign x_37996 = x_37992 & x_37995;
assign x_37997 = x_37989 & x_37996;
assign x_37998 = x_6708 & x_6709;
assign x_37999 = x_6710 & x_6711;
assign x_38000 = x_37998 & x_37999;
assign x_38001 = x_6712 & x_6713;
assign x_38002 = x_6714 & x_6715;
assign x_38003 = x_38001 & x_38002;
assign x_38004 = x_38000 & x_38003;
assign x_38005 = x_6716 & x_6717;
assign x_38006 = x_6718 & x_6719;
assign x_38007 = x_38005 & x_38006;
assign x_38008 = x_6720 & x_6721;
assign x_38009 = x_6722 & x_6723;
assign x_38010 = x_38008 & x_38009;
assign x_38011 = x_38007 & x_38010;
assign x_38012 = x_38004 & x_38011;
assign x_38013 = x_37997 & x_38012;
assign x_38014 = x_37983 & x_38013;
assign x_38015 = x_37954 & x_38014;
assign x_38016 = x_6725 & x_6726;
assign x_38017 = x_6724 & x_38016;
assign x_38018 = x_6727 & x_6728;
assign x_38019 = x_6729 & x_6730;
assign x_38020 = x_38018 & x_38019;
assign x_38021 = x_38017 & x_38020;
assign x_38022 = x_6731 & x_6732;
assign x_38023 = x_6733 & x_6734;
assign x_38024 = x_38022 & x_38023;
assign x_38025 = x_6735 & x_6736;
assign x_38026 = x_6737 & x_6738;
assign x_38027 = x_38025 & x_38026;
assign x_38028 = x_38024 & x_38027;
assign x_38029 = x_38021 & x_38028;
assign x_38030 = x_6740 & x_6741;
assign x_38031 = x_6739 & x_38030;
assign x_38032 = x_6742 & x_6743;
assign x_38033 = x_6744 & x_6745;
assign x_38034 = x_38032 & x_38033;
assign x_38035 = x_38031 & x_38034;
assign x_38036 = x_6746 & x_6747;
assign x_38037 = x_6748 & x_6749;
assign x_38038 = x_38036 & x_38037;
assign x_38039 = x_6750 & x_6751;
assign x_38040 = x_6752 & x_6753;
assign x_38041 = x_38039 & x_38040;
assign x_38042 = x_38038 & x_38041;
assign x_38043 = x_38035 & x_38042;
assign x_38044 = x_38029 & x_38043;
assign x_38045 = x_6755 & x_6756;
assign x_38046 = x_6754 & x_38045;
assign x_38047 = x_6757 & x_6758;
assign x_38048 = x_6759 & x_6760;
assign x_38049 = x_38047 & x_38048;
assign x_38050 = x_38046 & x_38049;
assign x_38051 = x_6761 & x_6762;
assign x_38052 = x_6763 & x_6764;
assign x_38053 = x_38051 & x_38052;
assign x_38054 = x_6765 & x_6766;
assign x_38055 = x_6767 & x_6768;
assign x_38056 = x_38054 & x_38055;
assign x_38057 = x_38053 & x_38056;
assign x_38058 = x_38050 & x_38057;
assign x_38059 = x_6769 & x_6770;
assign x_38060 = x_6771 & x_6772;
assign x_38061 = x_38059 & x_38060;
assign x_38062 = x_6773 & x_6774;
assign x_38063 = x_6775 & x_6776;
assign x_38064 = x_38062 & x_38063;
assign x_38065 = x_38061 & x_38064;
assign x_38066 = x_6777 & x_6778;
assign x_38067 = x_6779 & x_6780;
assign x_38068 = x_38066 & x_38067;
assign x_38069 = x_6781 & x_6782;
assign x_38070 = x_6783 & x_6784;
assign x_38071 = x_38069 & x_38070;
assign x_38072 = x_38068 & x_38071;
assign x_38073 = x_38065 & x_38072;
assign x_38074 = x_38058 & x_38073;
assign x_38075 = x_38044 & x_38074;
assign x_38076 = x_6786 & x_6787;
assign x_38077 = x_6785 & x_38076;
assign x_38078 = x_6788 & x_6789;
assign x_38079 = x_6790 & x_6791;
assign x_38080 = x_38078 & x_38079;
assign x_38081 = x_38077 & x_38080;
assign x_38082 = x_6792 & x_6793;
assign x_38083 = x_6794 & x_6795;
assign x_38084 = x_38082 & x_38083;
assign x_38085 = x_6796 & x_6797;
assign x_38086 = x_6798 & x_6799;
assign x_38087 = x_38085 & x_38086;
assign x_38088 = x_38084 & x_38087;
assign x_38089 = x_38081 & x_38088;
assign x_38090 = x_6800 & x_6801;
assign x_38091 = x_6802 & x_6803;
assign x_38092 = x_38090 & x_38091;
assign x_38093 = x_6804 & x_6805;
assign x_38094 = x_6806 & x_6807;
assign x_38095 = x_38093 & x_38094;
assign x_38096 = x_38092 & x_38095;
assign x_38097 = x_6808 & x_6809;
assign x_38098 = x_6810 & x_6811;
assign x_38099 = x_38097 & x_38098;
assign x_38100 = x_6812 & x_6813;
assign x_38101 = x_6814 & x_6815;
assign x_38102 = x_38100 & x_38101;
assign x_38103 = x_38099 & x_38102;
assign x_38104 = x_38096 & x_38103;
assign x_38105 = x_38089 & x_38104;
assign x_38106 = x_6817 & x_6818;
assign x_38107 = x_6816 & x_38106;
assign x_38108 = x_6819 & x_6820;
assign x_38109 = x_6821 & x_6822;
assign x_38110 = x_38108 & x_38109;
assign x_38111 = x_38107 & x_38110;
assign x_38112 = x_6823 & x_6824;
assign x_38113 = x_6825 & x_6826;
assign x_38114 = x_38112 & x_38113;
assign x_38115 = x_6827 & x_6828;
assign x_38116 = x_6829 & x_6830;
assign x_38117 = x_38115 & x_38116;
assign x_38118 = x_38114 & x_38117;
assign x_38119 = x_38111 & x_38118;
assign x_38120 = x_6831 & x_6832;
assign x_38121 = x_6833 & x_6834;
assign x_38122 = x_38120 & x_38121;
assign x_38123 = x_6835 & x_6836;
assign x_38124 = x_6837 & x_6838;
assign x_38125 = x_38123 & x_38124;
assign x_38126 = x_38122 & x_38125;
assign x_38127 = x_6839 & x_6840;
assign x_38128 = x_6841 & x_6842;
assign x_38129 = x_38127 & x_38128;
assign x_38130 = x_6843 & x_6844;
assign x_38131 = x_6845 & x_6846;
assign x_38132 = x_38130 & x_38131;
assign x_38133 = x_38129 & x_38132;
assign x_38134 = x_38126 & x_38133;
assign x_38135 = x_38119 & x_38134;
assign x_38136 = x_38105 & x_38135;
assign x_38137 = x_38075 & x_38136;
assign x_38138 = x_38015 & x_38137;
assign x_38139 = x_37894 & x_38138;
assign x_38140 = x_37651 & x_38139;
assign x_38141 = x_6848 & x_6849;
assign x_38142 = x_6847 & x_38141;
assign x_38143 = x_6850 & x_6851;
assign x_38144 = x_6852 & x_6853;
assign x_38145 = x_38143 & x_38144;
assign x_38146 = x_38142 & x_38145;
assign x_38147 = x_6854 & x_6855;
assign x_38148 = x_6856 & x_6857;
assign x_38149 = x_38147 & x_38148;
assign x_38150 = x_6858 & x_6859;
assign x_38151 = x_6860 & x_6861;
assign x_38152 = x_38150 & x_38151;
assign x_38153 = x_38149 & x_38152;
assign x_38154 = x_38146 & x_38153;
assign x_38155 = x_6863 & x_6864;
assign x_38156 = x_6862 & x_38155;
assign x_38157 = x_6865 & x_6866;
assign x_38158 = x_6867 & x_6868;
assign x_38159 = x_38157 & x_38158;
assign x_38160 = x_38156 & x_38159;
assign x_38161 = x_6869 & x_6870;
assign x_38162 = x_6871 & x_6872;
assign x_38163 = x_38161 & x_38162;
assign x_38164 = x_6873 & x_6874;
assign x_38165 = x_6875 & x_6876;
assign x_38166 = x_38164 & x_38165;
assign x_38167 = x_38163 & x_38166;
assign x_38168 = x_38160 & x_38167;
assign x_38169 = x_38154 & x_38168;
assign x_38170 = x_6878 & x_6879;
assign x_38171 = x_6877 & x_38170;
assign x_38172 = x_6880 & x_6881;
assign x_38173 = x_6882 & x_6883;
assign x_38174 = x_38172 & x_38173;
assign x_38175 = x_38171 & x_38174;
assign x_38176 = x_6884 & x_6885;
assign x_38177 = x_6886 & x_6887;
assign x_38178 = x_38176 & x_38177;
assign x_38179 = x_6888 & x_6889;
assign x_38180 = x_6890 & x_6891;
assign x_38181 = x_38179 & x_38180;
assign x_38182 = x_38178 & x_38181;
assign x_38183 = x_38175 & x_38182;
assign x_38184 = x_6892 & x_6893;
assign x_38185 = x_6894 & x_6895;
assign x_38186 = x_38184 & x_38185;
assign x_38187 = x_6896 & x_6897;
assign x_38188 = x_6898 & x_6899;
assign x_38189 = x_38187 & x_38188;
assign x_38190 = x_38186 & x_38189;
assign x_38191 = x_6900 & x_6901;
assign x_38192 = x_6902 & x_6903;
assign x_38193 = x_38191 & x_38192;
assign x_38194 = x_6904 & x_6905;
assign x_38195 = x_6906 & x_6907;
assign x_38196 = x_38194 & x_38195;
assign x_38197 = x_38193 & x_38196;
assign x_38198 = x_38190 & x_38197;
assign x_38199 = x_38183 & x_38198;
assign x_38200 = x_38169 & x_38199;
assign x_38201 = x_6909 & x_6910;
assign x_38202 = x_6908 & x_38201;
assign x_38203 = x_6911 & x_6912;
assign x_38204 = x_6913 & x_6914;
assign x_38205 = x_38203 & x_38204;
assign x_38206 = x_38202 & x_38205;
assign x_38207 = x_6915 & x_6916;
assign x_38208 = x_6917 & x_6918;
assign x_38209 = x_38207 & x_38208;
assign x_38210 = x_6919 & x_6920;
assign x_38211 = x_6921 & x_6922;
assign x_38212 = x_38210 & x_38211;
assign x_38213 = x_38209 & x_38212;
assign x_38214 = x_38206 & x_38213;
assign x_38215 = x_6924 & x_6925;
assign x_38216 = x_6923 & x_38215;
assign x_38217 = x_6926 & x_6927;
assign x_38218 = x_6928 & x_6929;
assign x_38219 = x_38217 & x_38218;
assign x_38220 = x_38216 & x_38219;
assign x_38221 = x_6930 & x_6931;
assign x_38222 = x_6932 & x_6933;
assign x_38223 = x_38221 & x_38222;
assign x_38224 = x_6934 & x_6935;
assign x_38225 = x_6936 & x_6937;
assign x_38226 = x_38224 & x_38225;
assign x_38227 = x_38223 & x_38226;
assign x_38228 = x_38220 & x_38227;
assign x_38229 = x_38214 & x_38228;
assign x_38230 = x_6939 & x_6940;
assign x_38231 = x_6938 & x_38230;
assign x_38232 = x_6941 & x_6942;
assign x_38233 = x_6943 & x_6944;
assign x_38234 = x_38232 & x_38233;
assign x_38235 = x_38231 & x_38234;
assign x_38236 = x_6945 & x_6946;
assign x_38237 = x_6947 & x_6948;
assign x_38238 = x_38236 & x_38237;
assign x_38239 = x_6949 & x_6950;
assign x_38240 = x_6951 & x_6952;
assign x_38241 = x_38239 & x_38240;
assign x_38242 = x_38238 & x_38241;
assign x_38243 = x_38235 & x_38242;
assign x_38244 = x_6953 & x_6954;
assign x_38245 = x_6955 & x_6956;
assign x_38246 = x_38244 & x_38245;
assign x_38247 = x_6957 & x_6958;
assign x_38248 = x_6959 & x_6960;
assign x_38249 = x_38247 & x_38248;
assign x_38250 = x_38246 & x_38249;
assign x_38251 = x_6961 & x_6962;
assign x_38252 = x_6963 & x_6964;
assign x_38253 = x_38251 & x_38252;
assign x_38254 = x_6965 & x_6966;
assign x_38255 = x_6967 & x_6968;
assign x_38256 = x_38254 & x_38255;
assign x_38257 = x_38253 & x_38256;
assign x_38258 = x_38250 & x_38257;
assign x_38259 = x_38243 & x_38258;
assign x_38260 = x_38229 & x_38259;
assign x_38261 = x_38200 & x_38260;
assign x_38262 = x_6970 & x_6971;
assign x_38263 = x_6969 & x_38262;
assign x_38264 = x_6972 & x_6973;
assign x_38265 = x_6974 & x_6975;
assign x_38266 = x_38264 & x_38265;
assign x_38267 = x_38263 & x_38266;
assign x_38268 = x_6976 & x_6977;
assign x_38269 = x_6978 & x_6979;
assign x_38270 = x_38268 & x_38269;
assign x_38271 = x_6980 & x_6981;
assign x_38272 = x_6982 & x_6983;
assign x_38273 = x_38271 & x_38272;
assign x_38274 = x_38270 & x_38273;
assign x_38275 = x_38267 & x_38274;
assign x_38276 = x_6985 & x_6986;
assign x_38277 = x_6984 & x_38276;
assign x_38278 = x_6987 & x_6988;
assign x_38279 = x_6989 & x_6990;
assign x_38280 = x_38278 & x_38279;
assign x_38281 = x_38277 & x_38280;
assign x_38282 = x_6991 & x_6992;
assign x_38283 = x_6993 & x_6994;
assign x_38284 = x_38282 & x_38283;
assign x_38285 = x_6995 & x_6996;
assign x_38286 = x_6997 & x_6998;
assign x_38287 = x_38285 & x_38286;
assign x_38288 = x_38284 & x_38287;
assign x_38289 = x_38281 & x_38288;
assign x_38290 = x_38275 & x_38289;
assign x_38291 = x_7000 & x_7001;
assign x_38292 = x_6999 & x_38291;
assign x_38293 = x_7002 & x_7003;
assign x_38294 = x_7004 & x_7005;
assign x_38295 = x_38293 & x_38294;
assign x_38296 = x_38292 & x_38295;
assign x_38297 = x_7006 & x_7007;
assign x_38298 = x_7008 & x_7009;
assign x_38299 = x_38297 & x_38298;
assign x_38300 = x_7010 & x_7011;
assign x_38301 = x_7012 & x_7013;
assign x_38302 = x_38300 & x_38301;
assign x_38303 = x_38299 & x_38302;
assign x_38304 = x_38296 & x_38303;
assign x_38305 = x_7014 & x_7015;
assign x_38306 = x_7016 & x_7017;
assign x_38307 = x_38305 & x_38306;
assign x_38308 = x_7018 & x_7019;
assign x_38309 = x_7020 & x_7021;
assign x_38310 = x_38308 & x_38309;
assign x_38311 = x_38307 & x_38310;
assign x_38312 = x_7022 & x_7023;
assign x_38313 = x_7024 & x_7025;
assign x_38314 = x_38312 & x_38313;
assign x_38315 = x_7026 & x_7027;
assign x_38316 = x_7028 & x_7029;
assign x_38317 = x_38315 & x_38316;
assign x_38318 = x_38314 & x_38317;
assign x_38319 = x_38311 & x_38318;
assign x_38320 = x_38304 & x_38319;
assign x_38321 = x_38290 & x_38320;
assign x_38322 = x_7031 & x_7032;
assign x_38323 = x_7030 & x_38322;
assign x_38324 = x_7033 & x_7034;
assign x_38325 = x_7035 & x_7036;
assign x_38326 = x_38324 & x_38325;
assign x_38327 = x_38323 & x_38326;
assign x_38328 = x_7037 & x_7038;
assign x_38329 = x_7039 & x_7040;
assign x_38330 = x_38328 & x_38329;
assign x_38331 = x_7041 & x_7042;
assign x_38332 = x_7043 & x_7044;
assign x_38333 = x_38331 & x_38332;
assign x_38334 = x_38330 & x_38333;
assign x_38335 = x_38327 & x_38334;
assign x_38336 = x_7046 & x_7047;
assign x_38337 = x_7045 & x_38336;
assign x_38338 = x_7048 & x_7049;
assign x_38339 = x_7050 & x_7051;
assign x_38340 = x_38338 & x_38339;
assign x_38341 = x_38337 & x_38340;
assign x_38342 = x_7052 & x_7053;
assign x_38343 = x_7054 & x_7055;
assign x_38344 = x_38342 & x_38343;
assign x_38345 = x_7056 & x_7057;
assign x_38346 = x_7058 & x_7059;
assign x_38347 = x_38345 & x_38346;
assign x_38348 = x_38344 & x_38347;
assign x_38349 = x_38341 & x_38348;
assign x_38350 = x_38335 & x_38349;
assign x_38351 = x_7061 & x_7062;
assign x_38352 = x_7060 & x_38351;
assign x_38353 = x_7063 & x_7064;
assign x_38354 = x_7065 & x_7066;
assign x_38355 = x_38353 & x_38354;
assign x_38356 = x_38352 & x_38355;
assign x_38357 = x_7067 & x_7068;
assign x_38358 = x_7069 & x_7070;
assign x_38359 = x_38357 & x_38358;
assign x_38360 = x_7071 & x_7072;
assign x_38361 = x_7073 & x_7074;
assign x_38362 = x_38360 & x_38361;
assign x_38363 = x_38359 & x_38362;
assign x_38364 = x_38356 & x_38363;
assign x_38365 = x_7075 & x_7076;
assign x_38366 = x_7077 & x_7078;
assign x_38367 = x_38365 & x_38366;
assign x_38368 = x_7079 & x_7080;
assign x_38369 = x_7081 & x_7082;
assign x_38370 = x_38368 & x_38369;
assign x_38371 = x_38367 & x_38370;
assign x_38372 = x_7083 & x_7084;
assign x_38373 = x_7085 & x_7086;
assign x_38374 = x_38372 & x_38373;
assign x_38375 = x_7087 & x_7088;
assign x_38376 = x_7089 & x_7090;
assign x_38377 = x_38375 & x_38376;
assign x_38378 = x_38374 & x_38377;
assign x_38379 = x_38371 & x_38378;
assign x_38380 = x_38364 & x_38379;
assign x_38381 = x_38350 & x_38380;
assign x_38382 = x_38321 & x_38381;
assign x_38383 = x_38261 & x_38382;
assign x_38384 = x_7092 & x_7093;
assign x_38385 = x_7091 & x_38384;
assign x_38386 = x_7094 & x_7095;
assign x_38387 = x_7096 & x_7097;
assign x_38388 = x_38386 & x_38387;
assign x_38389 = x_38385 & x_38388;
assign x_38390 = x_7098 & x_7099;
assign x_38391 = x_7100 & x_7101;
assign x_38392 = x_38390 & x_38391;
assign x_38393 = x_7102 & x_7103;
assign x_38394 = x_7104 & x_7105;
assign x_38395 = x_38393 & x_38394;
assign x_38396 = x_38392 & x_38395;
assign x_38397 = x_38389 & x_38396;
assign x_38398 = x_7107 & x_7108;
assign x_38399 = x_7106 & x_38398;
assign x_38400 = x_7109 & x_7110;
assign x_38401 = x_7111 & x_7112;
assign x_38402 = x_38400 & x_38401;
assign x_38403 = x_38399 & x_38402;
assign x_38404 = x_7113 & x_7114;
assign x_38405 = x_7115 & x_7116;
assign x_38406 = x_38404 & x_38405;
assign x_38407 = x_7117 & x_7118;
assign x_38408 = x_7119 & x_7120;
assign x_38409 = x_38407 & x_38408;
assign x_38410 = x_38406 & x_38409;
assign x_38411 = x_38403 & x_38410;
assign x_38412 = x_38397 & x_38411;
assign x_38413 = x_7122 & x_7123;
assign x_38414 = x_7121 & x_38413;
assign x_38415 = x_7124 & x_7125;
assign x_38416 = x_7126 & x_7127;
assign x_38417 = x_38415 & x_38416;
assign x_38418 = x_38414 & x_38417;
assign x_38419 = x_7128 & x_7129;
assign x_38420 = x_7130 & x_7131;
assign x_38421 = x_38419 & x_38420;
assign x_38422 = x_7132 & x_7133;
assign x_38423 = x_7134 & x_7135;
assign x_38424 = x_38422 & x_38423;
assign x_38425 = x_38421 & x_38424;
assign x_38426 = x_38418 & x_38425;
assign x_38427 = x_7136 & x_7137;
assign x_38428 = x_7138 & x_7139;
assign x_38429 = x_38427 & x_38428;
assign x_38430 = x_7140 & x_7141;
assign x_38431 = x_7142 & x_7143;
assign x_38432 = x_38430 & x_38431;
assign x_38433 = x_38429 & x_38432;
assign x_38434 = x_7144 & x_7145;
assign x_38435 = x_7146 & x_7147;
assign x_38436 = x_38434 & x_38435;
assign x_38437 = x_7148 & x_7149;
assign x_38438 = x_7150 & x_7151;
assign x_38439 = x_38437 & x_38438;
assign x_38440 = x_38436 & x_38439;
assign x_38441 = x_38433 & x_38440;
assign x_38442 = x_38426 & x_38441;
assign x_38443 = x_38412 & x_38442;
assign x_38444 = x_7153 & x_7154;
assign x_38445 = x_7152 & x_38444;
assign x_38446 = x_7155 & x_7156;
assign x_38447 = x_7157 & x_7158;
assign x_38448 = x_38446 & x_38447;
assign x_38449 = x_38445 & x_38448;
assign x_38450 = x_7159 & x_7160;
assign x_38451 = x_7161 & x_7162;
assign x_38452 = x_38450 & x_38451;
assign x_38453 = x_7163 & x_7164;
assign x_38454 = x_7165 & x_7166;
assign x_38455 = x_38453 & x_38454;
assign x_38456 = x_38452 & x_38455;
assign x_38457 = x_38449 & x_38456;
assign x_38458 = x_7168 & x_7169;
assign x_38459 = x_7167 & x_38458;
assign x_38460 = x_7170 & x_7171;
assign x_38461 = x_7172 & x_7173;
assign x_38462 = x_38460 & x_38461;
assign x_38463 = x_38459 & x_38462;
assign x_38464 = x_7174 & x_7175;
assign x_38465 = x_7176 & x_7177;
assign x_38466 = x_38464 & x_38465;
assign x_38467 = x_7178 & x_7179;
assign x_38468 = x_7180 & x_7181;
assign x_38469 = x_38467 & x_38468;
assign x_38470 = x_38466 & x_38469;
assign x_38471 = x_38463 & x_38470;
assign x_38472 = x_38457 & x_38471;
assign x_38473 = x_7183 & x_7184;
assign x_38474 = x_7182 & x_38473;
assign x_38475 = x_7185 & x_7186;
assign x_38476 = x_7187 & x_7188;
assign x_38477 = x_38475 & x_38476;
assign x_38478 = x_38474 & x_38477;
assign x_38479 = x_7189 & x_7190;
assign x_38480 = x_7191 & x_7192;
assign x_38481 = x_38479 & x_38480;
assign x_38482 = x_7193 & x_7194;
assign x_38483 = x_7195 & x_7196;
assign x_38484 = x_38482 & x_38483;
assign x_38485 = x_38481 & x_38484;
assign x_38486 = x_38478 & x_38485;
assign x_38487 = x_7197 & x_7198;
assign x_38488 = x_7199 & x_7200;
assign x_38489 = x_38487 & x_38488;
assign x_38490 = x_7201 & x_7202;
assign x_38491 = x_7203 & x_7204;
assign x_38492 = x_38490 & x_38491;
assign x_38493 = x_38489 & x_38492;
assign x_38494 = x_7205 & x_7206;
assign x_38495 = x_7207 & x_7208;
assign x_38496 = x_38494 & x_38495;
assign x_38497 = x_7209 & x_7210;
assign x_38498 = x_7211 & x_7212;
assign x_38499 = x_38497 & x_38498;
assign x_38500 = x_38496 & x_38499;
assign x_38501 = x_38493 & x_38500;
assign x_38502 = x_38486 & x_38501;
assign x_38503 = x_38472 & x_38502;
assign x_38504 = x_38443 & x_38503;
assign x_38505 = x_7214 & x_7215;
assign x_38506 = x_7213 & x_38505;
assign x_38507 = x_7216 & x_7217;
assign x_38508 = x_7218 & x_7219;
assign x_38509 = x_38507 & x_38508;
assign x_38510 = x_38506 & x_38509;
assign x_38511 = x_7220 & x_7221;
assign x_38512 = x_7222 & x_7223;
assign x_38513 = x_38511 & x_38512;
assign x_38514 = x_7224 & x_7225;
assign x_38515 = x_7226 & x_7227;
assign x_38516 = x_38514 & x_38515;
assign x_38517 = x_38513 & x_38516;
assign x_38518 = x_38510 & x_38517;
assign x_38519 = x_7229 & x_7230;
assign x_38520 = x_7228 & x_38519;
assign x_38521 = x_7231 & x_7232;
assign x_38522 = x_7233 & x_7234;
assign x_38523 = x_38521 & x_38522;
assign x_38524 = x_38520 & x_38523;
assign x_38525 = x_7235 & x_7236;
assign x_38526 = x_7237 & x_7238;
assign x_38527 = x_38525 & x_38526;
assign x_38528 = x_7239 & x_7240;
assign x_38529 = x_7241 & x_7242;
assign x_38530 = x_38528 & x_38529;
assign x_38531 = x_38527 & x_38530;
assign x_38532 = x_38524 & x_38531;
assign x_38533 = x_38518 & x_38532;
assign x_38534 = x_7244 & x_7245;
assign x_38535 = x_7243 & x_38534;
assign x_38536 = x_7246 & x_7247;
assign x_38537 = x_7248 & x_7249;
assign x_38538 = x_38536 & x_38537;
assign x_38539 = x_38535 & x_38538;
assign x_38540 = x_7250 & x_7251;
assign x_38541 = x_7252 & x_7253;
assign x_38542 = x_38540 & x_38541;
assign x_38543 = x_7254 & x_7255;
assign x_38544 = x_7256 & x_7257;
assign x_38545 = x_38543 & x_38544;
assign x_38546 = x_38542 & x_38545;
assign x_38547 = x_38539 & x_38546;
assign x_38548 = x_7258 & x_7259;
assign x_38549 = x_7260 & x_7261;
assign x_38550 = x_38548 & x_38549;
assign x_38551 = x_7262 & x_7263;
assign x_38552 = x_7264 & x_7265;
assign x_38553 = x_38551 & x_38552;
assign x_38554 = x_38550 & x_38553;
assign x_38555 = x_7266 & x_7267;
assign x_38556 = x_7268 & x_7269;
assign x_38557 = x_38555 & x_38556;
assign x_38558 = x_7270 & x_7271;
assign x_38559 = x_7272 & x_7273;
assign x_38560 = x_38558 & x_38559;
assign x_38561 = x_38557 & x_38560;
assign x_38562 = x_38554 & x_38561;
assign x_38563 = x_38547 & x_38562;
assign x_38564 = x_38533 & x_38563;
assign x_38565 = x_7275 & x_7276;
assign x_38566 = x_7274 & x_38565;
assign x_38567 = x_7277 & x_7278;
assign x_38568 = x_7279 & x_7280;
assign x_38569 = x_38567 & x_38568;
assign x_38570 = x_38566 & x_38569;
assign x_38571 = x_7281 & x_7282;
assign x_38572 = x_7283 & x_7284;
assign x_38573 = x_38571 & x_38572;
assign x_38574 = x_7285 & x_7286;
assign x_38575 = x_7287 & x_7288;
assign x_38576 = x_38574 & x_38575;
assign x_38577 = x_38573 & x_38576;
assign x_38578 = x_38570 & x_38577;
assign x_38579 = x_7289 & x_7290;
assign x_38580 = x_7291 & x_7292;
assign x_38581 = x_38579 & x_38580;
assign x_38582 = x_7293 & x_7294;
assign x_38583 = x_7295 & x_7296;
assign x_38584 = x_38582 & x_38583;
assign x_38585 = x_38581 & x_38584;
assign x_38586 = x_7297 & x_7298;
assign x_38587 = x_7299 & x_7300;
assign x_38588 = x_38586 & x_38587;
assign x_38589 = x_7301 & x_7302;
assign x_38590 = x_7303 & x_7304;
assign x_38591 = x_38589 & x_38590;
assign x_38592 = x_38588 & x_38591;
assign x_38593 = x_38585 & x_38592;
assign x_38594 = x_38578 & x_38593;
assign x_38595 = x_7306 & x_7307;
assign x_38596 = x_7305 & x_38595;
assign x_38597 = x_7308 & x_7309;
assign x_38598 = x_7310 & x_7311;
assign x_38599 = x_38597 & x_38598;
assign x_38600 = x_38596 & x_38599;
assign x_38601 = x_7312 & x_7313;
assign x_38602 = x_7314 & x_7315;
assign x_38603 = x_38601 & x_38602;
assign x_38604 = x_7316 & x_7317;
assign x_38605 = x_7318 & x_7319;
assign x_38606 = x_38604 & x_38605;
assign x_38607 = x_38603 & x_38606;
assign x_38608 = x_38600 & x_38607;
assign x_38609 = x_7320 & x_7321;
assign x_38610 = x_7322 & x_7323;
assign x_38611 = x_38609 & x_38610;
assign x_38612 = x_7324 & x_7325;
assign x_38613 = x_7326 & x_7327;
assign x_38614 = x_38612 & x_38613;
assign x_38615 = x_38611 & x_38614;
assign x_38616 = x_7328 & x_7329;
assign x_38617 = x_7330 & x_7331;
assign x_38618 = x_38616 & x_38617;
assign x_38619 = x_7332 & x_7333;
assign x_38620 = x_7334 & x_7335;
assign x_38621 = x_38619 & x_38620;
assign x_38622 = x_38618 & x_38621;
assign x_38623 = x_38615 & x_38622;
assign x_38624 = x_38608 & x_38623;
assign x_38625 = x_38594 & x_38624;
assign x_38626 = x_38564 & x_38625;
assign x_38627 = x_38504 & x_38626;
assign x_38628 = x_38383 & x_38627;
assign x_38629 = x_7337 & x_7338;
assign x_38630 = x_7336 & x_38629;
assign x_38631 = x_7339 & x_7340;
assign x_38632 = x_7341 & x_7342;
assign x_38633 = x_38631 & x_38632;
assign x_38634 = x_38630 & x_38633;
assign x_38635 = x_7343 & x_7344;
assign x_38636 = x_7345 & x_7346;
assign x_38637 = x_38635 & x_38636;
assign x_38638 = x_7347 & x_7348;
assign x_38639 = x_7349 & x_7350;
assign x_38640 = x_38638 & x_38639;
assign x_38641 = x_38637 & x_38640;
assign x_38642 = x_38634 & x_38641;
assign x_38643 = x_7352 & x_7353;
assign x_38644 = x_7351 & x_38643;
assign x_38645 = x_7354 & x_7355;
assign x_38646 = x_7356 & x_7357;
assign x_38647 = x_38645 & x_38646;
assign x_38648 = x_38644 & x_38647;
assign x_38649 = x_7358 & x_7359;
assign x_38650 = x_7360 & x_7361;
assign x_38651 = x_38649 & x_38650;
assign x_38652 = x_7362 & x_7363;
assign x_38653 = x_7364 & x_7365;
assign x_38654 = x_38652 & x_38653;
assign x_38655 = x_38651 & x_38654;
assign x_38656 = x_38648 & x_38655;
assign x_38657 = x_38642 & x_38656;
assign x_38658 = x_7367 & x_7368;
assign x_38659 = x_7366 & x_38658;
assign x_38660 = x_7369 & x_7370;
assign x_38661 = x_7371 & x_7372;
assign x_38662 = x_38660 & x_38661;
assign x_38663 = x_38659 & x_38662;
assign x_38664 = x_7373 & x_7374;
assign x_38665 = x_7375 & x_7376;
assign x_38666 = x_38664 & x_38665;
assign x_38667 = x_7377 & x_7378;
assign x_38668 = x_7379 & x_7380;
assign x_38669 = x_38667 & x_38668;
assign x_38670 = x_38666 & x_38669;
assign x_38671 = x_38663 & x_38670;
assign x_38672 = x_7381 & x_7382;
assign x_38673 = x_7383 & x_7384;
assign x_38674 = x_38672 & x_38673;
assign x_38675 = x_7385 & x_7386;
assign x_38676 = x_7387 & x_7388;
assign x_38677 = x_38675 & x_38676;
assign x_38678 = x_38674 & x_38677;
assign x_38679 = x_7389 & x_7390;
assign x_38680 = x_7391 & x_7392;
assign x_38681 = x_38679 & x_38680;
assign x_38682 = x_7393 & x_7394;
assign x_38683 = x_7395 & x_7396;
assign x_38684 = x_38682 & x_38683;
assign x_38685 = x_38681 & x_38684;
assign x_38686 = x_38678 & x_38685;
assign x_38687 = x_38671 & x_38686;
assign x_38688 = x_38657 & x_38687;
assign x_38689 = x_7398 & x_7399;
assign x_38690 = x_7397 & x_38689;
assign x_38691 = x_7400 & x_7401;
assign x_38692 = x_7402 & x_7403;
assign x_38693 = x_38691 & x_38692;
assign x_38694 = x_38690 & x_38693;
assign x_38695 = x_7404 & x_7405;
assign x_38696 = x_7406 & x_7407;
assign x_38697 = x_38695 & x_38696;
assign x_38698 = x_7408 & x_7409;
assign x_38699 = x_7410 & x_7411;
assign x_38700 = x_38698 & x_38699;
assign x_38701 = x_38697 & x_38700;
assign x_38702 = x_38694 & x_38701;
assign x_38703 = x_7413 & x_7414;
assign x_38704 = x_7412 & x_38703;
assign x_38705 = x_7415 & x_7416;
assign x_38706 = x_7417 & x_7418;
assign x_38707 = x_38705 & x_38706;
assign x_38708 = x_38704 & x_38707;
assign x_38709 = x_7419 & x_7420;
assign x_38710 = x_7421 & x_7422;
assign x_38711 = x_38709 & x_38710;
assign x_38712 = x_7423 & x_7424;
assign x_38713 = x_7425 & x_7426;
assign x_38714 = x_38712 & x_38713;
assign x_38715 = x_38711 & x_38714;
assign x_38716 = x_38708 & x_38715;
assign x_38717 = x_38702 & x_38716;
assign x_38718 = x_7428 & x_7429;
assign x_38719 = x_7427 & x_38718;
assign x_38720 = x_7430 & x_7431;
assign x_38721 = x_7432 & x_7433;
assign x_38722 = x_38720 & x_38721;
assign x_38723 = x_38719 & x_38722;
assign x_38724 = x_7434 & x_7435;
assign x_38725 = x_7436 & x_7437;
assign x_38726 = x_38724 & x_38725;
assign x_38727 = x_7438 & x_7439;
assign x_38728 = x_7440 & x_7441;
assign x_38729 = x_38727 & x_38728;
assign x_38730 = x_38726 & x_38729;
assign x_38731 = x_38723 & x_38730;
assign x_38732 = x_7442 & x_7443;
assign x_38733 = x_7444 & x_7445;
assign x_38734 = x_38732 & x_38733;
assign x_38735 = x_7446 & x_7447;
assign x_38736 = x_7448 & x_7449;
assign x_38737 = x_38735 & x_38736;
assign x_38738 = x_38734 & x_38737;
assign x_38739 = x_7450 & x_7451;
assign x_38740 = x_7452 & x_7453;
assign x_38741 = x_38739 & x_38740;
assign x_38742 = x_7454 & x_7455;
assign x_38743 = x_7456 & x_7457;
assign x_38744 = x_38742 & x_38743;
assign x_38745 = x_38741 & x_38744;
assign x_38746 = x_38738 & x_38745;
assign x_38747 = x_38731 & x_38746;
assign x_38748 = x_38717 & x_38747;
assign x_38749 = x_38688 & x_38748;
assign x_38750 = x_7459 & x_7460;
assign x_38751 = x_7458 & x_38750;
assign x_38752 = x_7461 & x_7462;
assign x_38753 = x_7463 & x_7464;
assign x_38754 = x_38752 & x_38753;
assign x_38755 = x_38751 & x_38754;
assign x_38756 = x_7465 & x_7466;
assign x_38757 = x_7467 & x_7468;
assign x_38758 = x_38756 & x_38757;
assign x_38759 = x_7469 & x_7470;
assign x_38760 = x_7471 & x_7472;
assign x_38761 = x_38759 & x_38760;
assign x_38762 = x_38758 & x_38761;
assign x_38763 = x_38755 & x_38762;
assign x_38764 = x_7474 & x_7475;
assign x_38765 = x_7473 & x_38764;
assign x_38766 = x_7476 & x_7477;
assign x_38767 = x_7478 & x_7479;
assign x_38768 = x_38766 & x_38767;
assign x_38769 = x_38765 & x_38768;
assign x_38770 = x_7480 & x_7481;
assign x_38771 = x_7482 & x_7483;
assign x_38772 = x_38770 & x_38771;
assign x_38773 = x_7484 & x_7485;
assign x_38774 = x_7486 & x_7487;
assign x_38775 = x_38773 & x_38774;
assign x_38776 = x_38772 & x_38775;
assign x_38777 = x_38769 & x_38776;
assign x_38778 = x_38763 & x_38777;
assign x_38779 = x_7489 & x_7490;
assign x_38780 = x_7488 & x_38779;
assign x_38781 = x_7491 & x_7492;
assign x_38782 = x_7493 & x_7494;
assign x_38783 = x_38781 & x_38782;
assign x_38784 = x_38780 & x_38783;
assign x_38785 = x_7495 & x_7496;
assign x_38786 = x_7497 & x_7498;
assign x_38787 = x_38785 & x_38786;
assign x_38788 = x_7499 & x_7500;
assign x_38789 = x_7501 & x_7502;
assign x_38790 = x_38788 & x_38789;
assign x_38791 = x_38787 & x_38790;
assign x_38792 = x_38784 & x_38791;
assign x_38793 = x_7503 & x_7504;
assign x_38794 = x_7505 & x_7506;
assign x_38795 = x_38793 & x_38794;
assign x_38796 = x_7507 & x_7508;
assign x_38797 = x_7509 & x_7510;
assign x_38798 = x_38796 & x_38797;
assign x_38799 = x_38795 & x_38798;
assign x_38800 = x_7511 & x_7512;
assign x_38801 = x_7513 & x_7514;
assign x_38802 = x_38800 & x_38801;
assign x_38803 = x_7515 & x_7516;
assign x_38804 = x_7517 & x_7518;
assign x_38805 = x_38803 & x_38804;
assign x_38806 = x_38802 & x_38805;
assign x_38807 = x_38799 & x_38806;
assign x_38808 = x_38792 & x_38807;
assign x_38809 = x_38778 & x_38808;
assign x_38810 = x_7520 & x_7521;
assign x_38811 = x_7519 & x_38810;
assign x_38812 = x_7522 & x_7523;
assign x_38813 = x_7524 & x_7525;
assign x_38814 = x_38812 & x_38813;
assign x_38815 = x_38811 & x_38814;
assign x_38816 = x_7526 & x_7527;
assign x_38817 = x_7528 & x_7529;
assign x_38818 = x_38816 & x_38817;
assign x_38819 = x_7530 & x_7531;
assign x_38820 = x_7532 & x_7533;
assign x_38821 = x_38819 & x_38820;
assign x_38822 = x_38818 & x_38821;
assign x_38823 = x_38815 & x_38822;
assign x_38824 = x_7535 & x_7536;
assign x_38825 = x_7534 & x_38824;
assign x_38826 = x_7537 & x_7538;
assign x_38827 = x_7539 & x_7540;
assign x_38828 = x_38826 & x_38827;
assign x_38829 = x_38825 & x_38828;
assign x_38830 = x_7541 & x_7542;
assign x_38831 = x_7543 & x_7544;
assign x_38832 = x_38830 & x_38831;
assign x_38833 = x_7545 & x_7546;
assign x_38834 = x_7547 & x_7548;
assign x_38835 = x_38833 & x_38834;
assign x_38836 = x_38832 & x_38835;
assign x_38837 = x_38829 & x_38836;
assign x_38838 = x_38823 & x_38837;
assign x_38839 = x_7550 & x_7551;
assign x_38840 = x_7549 & x_38839;
assign x_38841 = x_7552 & x_7553;
assign x_38842 = x_7554 & x_7555;
assign x_38843 = x_38841 & x_38842;
assign x_38844 = x_38840 & x_38843;
assign x_38845 = x_7556 & x_7557;
assign x_38846 = x_7558 & x_7559;
assign x_38847 = x_38845 & x_38846;
assign x_38848 = x_7560 & x_7561;
assign x_38849 = x_7562 & x_7563;
assign x_38850 = x_38848 & x_38849;
assign x_38851 = x_38847 & x_38850;
assign x_38852 = x_38844 & x_38851;
assign x_38853 = x_7564 & x_7565;
assign x_38854 = x_7566 & x_7567;
assign x_38855 = x_38853 & x_38854;
assign x_38856 = x_7568 & x_7569;
assign x_38857 = x_7570 & x_7571;
assign x_38858 = x_38856 & x_38857;
assign x_38859 = x_38855 & x_38858;
assign x_38860 = x_7572 & x_7573;
assign x_38861 = x_7574 & x_7575;
assign x_38862 = x_38860 & x_38861;
assign x_38863 = x_7576 & x_7577;
assign x_38864 = x_7578 & x_7579;
assign x_38865 = x_38863 & x_38864;
assign x_38866 = x_38862 & x_38865;
assign x_38867 = x_38859 & x_38866;
assign x_38868 = x_38852 & x_38867;
assign x_38869 = x_38838 & x_38868;
assign x_38870 = x_38809 & x_38869;
assign x_38871 = x_38749 & x_38870;
assign x_38872 = x_7581 & x_7582;
assign x_38873 = x_7580 & x_38872;
assign x_38874 = x_7583 & x_7584;
assign x_38875 = x_7585 & x_7586;
assign x_38876 = x_38874 & x_38875;
assign x_38877 = x_38873 & x_38876;
assign x_38878 = x_7587 & x_7588;
assign x_38879 = x_7589 & x_7590;
assign x_38880 = x_38878 & x_38879;
assign x_38881 = x_7591 & x_7592;
assign x_38882 = x_7593 & x_7594;
assign x_38883 = x_38881 & x_38882;
assign x_38884 = x_38880 & x_38883;
assign x_38885 = x_38877 & x_38884;
assign x_38886 = x_7596 & x_7597;
assign x_38887 = x_7595 & x_38886;
assign x_38888 = x_7598 & x_7599;
assign x_38889 = x_7600 & x_7601;
assign x_38890 = x_38888 & x_38889;
assign x_38891 = x_38887 & x_38890;
assign x_38892 = x_7602 & x_7603;
assign x_38893 = x_7604 & x_7605;
assign x_38894 = x_38892 & x_38893;
assign x_38895 = x_7606 & x_7607;
assign x_38896 = x_7608 & x_7609;
assign x_38897 = x_38895 & x_38896;
assign x_38898 = x_38894 & x_38897;
assign x_38899 = x_38891 & x_38898;
assign x_38900 = x_38885 & x_38899;
assign x_38901 = x_7611 & x_7612;
assign x_38902 = x_7610 & x_38901;
assign x_38903 = x_7613 & x_7614;
assign x_38904 = x_7615 & x_7616;
assign x_38905 = x_38903 & x_38904;
assign x_38906 = x_38902 & x_38905;
assign x_38907 = x_7617 & x_7618;
assign x_38908 = x_7619 & x_7620;
assign x_38909 = x_38907 & x_38908;
assign x_38910 = x_7621 & x_7622;
assign x_38911 = x_7623 & x_7624;
assign x_38912 = x_38910 & x_38911;
assign x_38913 = x_38909 & x_38912;
assign x_38914 = x_38906 & x_38913;
assign x_38915 = x_7625 & x_7626;
assign x_38916 = x_7627 & x_7628;
assign x_38917 = x_38915 & x_38916;
assign x_38918 = x_7629 & x_7630;
assign x_38919 = x_7631 & x_7632;
assign x_38920 = x_38918 & x_38919;
assign x_38921 = x_38917 & x_38920;
assign x_38922 = x_7633 & x_7634;
assign x_38923 = x_7635 & x_7636;
assign x_38924 = x_38922 & x_38923;
assign x_38925 = x_7637 & x_7638;
assign x_38926 = x_7639 & x_7640;
assign x_38927 = x_38925 & x_38926;
assign x_38928 = x_38924 & x_38927;
assign x_38929 = x_38921 & x_38928;
assign x_38930 = x_38914 & x_38929;
assign x_38931 = x_38900 & x_38930;
assign x_38932 = x_7642 & x_7643;
assign x_38933 = x_7641 & x_38932;
assign x_38934 = x_7644 & x_7645;
assign x_38935 = x_7646 & x_7647;
assign x_38936 = x_38934 & x_38935;
assign x_38937 = x_38933 & x_38936;
assign x_38938 = x_7648 & x_7649;
assign x_38939 = x_7650 & x_7651;
assign x_38940 = x_38938 & x_38939;
assign x_38941 = x_7652 & x_7653;
assign x_38942 = x_7654 & x_7655;
assign x_38943 = x_38941 & x_38942;
assign x_38944 = x_38940 & x_38943;
assign x_38945 = x_38937 & x_38944;
assign x_38946 = x_7657 & x_7658;
assign x_38947 = x_7656 & x_38946;
assign x_38948 = x_7659 & x_7660;
assign x_38949 = x_7661 & x_7662;
assign x_38950 = x_38948 & x_38949;
assign x_38951 = x_38947 & x_38950;
assign x_38952 = x_7663 & x_7664;
assign x_38953 = x_7665 & x_7666;
assign x_38954 = x_38952 & x_38953;
assign x_38955 = x_7667 & x_7668;
assign x_38956 = x_7669 & x_7670;
assign x_38957 = x_38955 & x_38956;
assign x_38958 = x_38954 & x_38957;
assign x_38959 = x_38951 & x_38958;
assign x_38960 = x_38945 & x_38959;
assign x_38961 = x_7672 & x_7673;
assign x_38962 = x_7671 & x_38961;
assign x_38963 = x_7674 & x_7675;
assign x_38964 = x_7676 & x_7677;
assign x_38965 = x_38963 & x_38964;
assign x_38966 = x_38962 & x_38965;
assign x_38967 = x_7678 & x_7679;
assign x_38968 = x_7680 & x_7681;
assign x_38969 = x_38967 & x_38968;
assign x_38970 = x_7682 & x_7683;
assign x_38971 = x_7684 & x_7685;
assign x_38972 = x_38970 & x_38971;
assign x_38973 = x_38969 & x_38972;
assign x_38974 = x_38966 & x_38973;
assign x_38975 = x_7686 & x_7687;
assign x_38976 = x_7688 & x_7689;
assign x_38977 = x_38975 & x_38976;
assign x_38978 = x_7690 & x_7691;
assign x_38979 = x_7692 & x_7693;
assign x_38980 = x_38978 & x_38979;
assign x_38981 = x_38977 & x_38980;
assign x_38982 = x_7694 & x_7695;
assign x_38983 = x_7696 & x_7697;
assign x_38984 = x_38982 & x_38983;
assign x_38985 = x_7698 & x_7699;
assign x_38986 = x_7700 & x_7701;
assign x_38987 = x_38985 & x_38986;
assign x_38988 = x_38984 & x_38987;
assign x_38989 = x_38981 & x_38988;
assign x_38990 = x_38974 & x_38989;
assign x_38991 = x_38960 & x_38990;
assign x_38992 = x_38931 & x_38991;
assign x_38993 = x_7703 & x_7704;
assign x_38994 = x_7702 & x_38993;
assign x_38995 = x_7705 & x_7706;
assign x_38996 = x_7707 & x_7708;
assign x_38997 = x_38995 & x_38996;
assign x_38998 = x_38994 & x_38997;
assign x_38999 = x_7709 & x_7710;
assign x_39000 = x_7711 & x_7712;
assign x_39001 = x_38999 & x_39000;
assign x_39002 = x_7713 & x_7714;
assign x_39003 = x_7715 & x_7716;
assign x_39004 = x_39002 & x_39003;
assign x_39005 = x_39001 & x_39004;
assign x_39006 = x_38998 & x_39005;
assign x_39007 = x_7718 & x_7719;
assign x_39008 = x_7717 & x_39007;
assign x_39009 = x_7720 & x_7721;
assign x_39010 = x_7722 & x_7723;
assign x_39011 = x_39009 & x_39010;
assign x_39012 = x_39008 & x_39011;
assign x_39013 = x_7724 & x_7725;
assign x_39014 = x_7726 & x_7727;
assign x_39015 = x_39013 & x_39014;
assign x_39016 = x_7728 & x_7729;
assign x_39017 = x_7730 & x_7731;
assign x_39018 = x_39016 & x_39017;
assign x_39019 = x_39015 & x_39018;
assign x_39020 = x_39012 & x_39019;
assign x_39021 = x_39006 & x_39020;
assign x_39022 = x_7733 & x_7734;
assign x_39023 = x_7732 & x_39022;
assign x_39024 = x_7735 & x_7736;
assign x_39025 = x_7737 & x_7738;
assign x_39026 = x_39024 & x_39025;
assign x_39027 = x_39023 & x_39026;
assign x_39028 = x_7739 & x_7740;
assign x_39029 = x_7741 & x_7742;
assign x_39030 = x_39028 & x_39029;
assign x_39031 = x_7743 & x_7744;
assign x_39032 = x_7745 & x_7746;
assign x_39033 = x_39031 & x_39032;
assign x_39034 = x_39030 & x_39033;
assign x_39035 = x_39027 & x_39034;
assign x_39036 = x_7747 & x_7748;
assign x_39037 = x_7749 & x_7750;
assign x_39038 = x_39036 & x_39037;
assign x_39039 = x_7751 & x_7752;
assign x_39040 = x_7753 & x_7754;
assign x_39041 = x_39039 & x_39040;
assign x_39042 = x_39038 & x_39041;
assign x_39043 = x_7755 & x_7756;
assign x_39044 = x_7757 & x_7758;
assign x_39045 = x_39043 & x_39044;
assign x_39046 = x_7759 & x_7760;
assign x_39047 = x_7761 & x_7762;
assign x_39048 = x_39046 & x_39047;
assign x_39049 = x_39045 & x_39048;
assign x_39050 = x_39042 & x_39049;
assign x_39051 = x_39035 & x_39050;
assign x_39052 = x_39021 & x_39051;
assign x_39053 = x_7764 & x_7765;
assign x_39054 = x_7763 & x_39053;
assign x_39055 = x_7766 & x_7767;
assign x_39056 = x_7768 & x_7769;
assign x_39057 = x_39055 & x_39056;
assign x_39058 = x_39054 & x_39057;
assign x_39059 = x_7770 & x_7771;
assign x_39060 = x_7772 & x_7773;
assign x_39061 = x_39059 & x_39060;
assign x_39062 = x_7774 & x_7775;
assign x_39063 = x_7776 & x_7777;
assign x_39064 = x_39062 & x_39063;
assign x_39065 = x_39061 & x_39064;
assign x_39066 = x_39058 & x_39065;
assign x_39067 = x_7778 & x_7779;
assign x_39068 = x_7780 & x_7781;
assign x_39069 = x_39067 & x_39068;
assign x_39070 = x_7782 & x_7783;
assign x_39071 = x_7784 & x_7785;
assign x_39072 = x_39070 & x_39071;
assign x_39073 = x_39069 & x_39072;
assign x_39074 = x_7786 & x_7787;
assign x_39075 = x_7788 & x_7789;
assign x_39076 = x_39074 & x_39075;
assign x_39077 = x_7790 & x_7791;
assign x_39078 = x_7792 & x_7793;
assign x_39079 = x_39077 & x_39078;
assign x_39080 = x_39076 & x_39079;
assign x_39081 = x_39073 & x_39080;
assign x_39082 = x_39066 & x_39081;
assign x_39083 = x_7795 & x_7796;
assign x_39084 = x_7794 & x_39083;
assign x_39085 = x_7797 & x_7798;
assign x_39086 = x_7799 & x_7800;
assign x_39087 = x_39085 & x_39086;
assign x_39088 = x_39084 & x_39087;
assign x_39089 = x_7801 & x_7802;
assign x_39090 = x_7803 & x_7804;
assign x_39091 = x_39089 & x_39090;
assign x_39092 = x_7805 & x_7806;
assign x_39093 = x_7807 & x_7808;
assign x_39094 = x_39092 & x_39093;
assign x_39095 = x_39091 & x_39094;
assign x_39096 = x_39088 & x_39095;
assign x_39097 = x_7809 & x_7810;
assign x_39098 = x_7811 & x_7812;
assign x_39099 = x_39097 & x_39098;
assign x_39100 = x_7813 & x_7814;
assign x_39101 = x_7815 & x_7816;
assign x_39102 = x_39100 & x_39101;
assign x_39103 = x_39099 & x_39102;
assign x_39104 = x_7817 & x_7818;
assign x_39105 = x_7819 & x_7820;
assign x_39106 = x_39104 & x_39105;
assign x_39107 = x_7821 & x_7822;
assign x_39108 = x_7823 & x_7824;
assign x_39109 = x_39107 & x_39108;
assign x_39110 = x_39106 & x_39109;
assign x_39111 = x_39103 & x_39110;
assign x_39112 = x_39096 & x_39111;
assign x_39113 = x_39082 & x_39112;
assign x_39114 = x_39052 & x_39113;
assign x_39115 = x_38992 & x_39114;
assign x_39116 = x_38871 & x_39115;
assign x_39117 = x_38628 & x_39116;
assign x_39118 = x_38140 & x_39117;
assign x_39119 = x_37163 & x_39118;
assign x_39120 = x_35208 & x_39119;
assign x_39121 = x_7826 & x_7827;
assign x_39122 = x_7825 & x_39121;
assign x_39123 = x_7828 & x_7829;
assign x_39124 = x_7830 & x_7831;
assign x_39125 = x_39123 & x_39124;
assign x_39126 = x_39122 & x_39125;
assign x_39127 = x_7832 & x_7833;
assign x_39128 = x_7834 & x_7835;
assign x_39129 = x_39127 & x_39128;
assign x_39130 = x_7836 & x_7837;
assign x_39131 = x_7838 & x_7839;
assign x_39132 = x_39130 & x_39131;
assign x_39133 = x_39129 & x_39132;
assign x_39134 = x_39126 & x_39133;
assign x_39135 = x_7841 & x_7842;
assign x_39136 = x_7840 & x_39135;
assign x_39137 = x_7843 & x_7844;
assign x_39138 = x_7845 & x_7846;
assign x_39139 = x_39137 & x_39138;
assign x_39140 = x_39136 & x_39139;
assign x_39141 = x_7847 & x_7848;
assign x_39142 = x_7849 & x_7850;
assign x_39143 = x_39141 & x_39142;
assign x_39144 = x_7851 & x_7852;
assign x_39145 = x_7853 & x_7854;
assign x_39146 = x_39144 & x_39145;
assign x_39147 = x_39143 & x_39146;
assign x_39148 = x_39140 & x_39147;
assign x_39149 = x_39134 & x_39148;
assign x_39150 = x_7856 & x_7857;
assign x_39151 = x_7855 & x_39150;
assign x_39152 = x_7858 & x_7859;
assign x_39153 = x_7860 & x_7861;
assign x_39154 = x_39152 & x_39153;
assign x_39155 = x_39151 & x_39154;
assign x_39156 = x_7862 & x_7863;
assign x_39157 = x_7864 & x_7865;
assign x_39158 = x_39156 & x_39157;
assign x_39159 = x_7866 & x_7867;
assign x_39160 = x_7868 & x_7869;
assign x_39161 = x_39159 & x_39160;
assign x_39162 = x_39158 & x_39161;
assign x_39163 = x_39155 & x_39162;
assign x_39164 = x_7870 & x_7871;
assign x_39165 = x_7872 & x_7873;
assign x_39166 = x_39164 & x_39165;
assign x_39167 = x_7874 & x_7875;
assign x_39168 = x_7876 & x_7877;
assign x_39169 = x_39167 & x_39168;
assign x_39170 = x_39166 & x_39169;
assign x_39171 = x_7878 & x_7879;
assign x_39172 = x_7880 & x_7881;
assign x_39173 = x_39171 & x_39172;
assign x_39174 = x_7882 & x_7883;
assign x_39175 = x_7884 & x_7885;
assign x_39176 = x_39174 & x_39175;
assign x_39177 = x_39173 & x_39176;
assign x_39178 = x_39170 & x_39177;
assign x_39179 = x_39163 & x_39178;
assign x_39180 = x_39149 & x_39179;
assign x_39181 = x_7887 & x_7888;
assign x_39182 = x_7886 & x_39181;
assign x_39183 = x_7889 & x_7890;
assign x_39184 = x_7891 & x_7892;
assign x_39185 = x_39183 & x_39184;
assign x_39186 = x_39182 & x_39185;
assign x_39187 = x_7893 & x_7894;
assign x_39188 = x_7895 & x_7896;
assign x_39189 = x_39187 & x_39188;
assign x_39190 = x_7897 & x_7898;
assign x_39191 = x_7899 & x_7900;
assign x_39192 = x_39190 & x_39191;
assign x_39193 = x_39189 & x_39192;
assign x_39194 = x_39186 & x_39193;
assign x_39195 = x_7902 & x_7903;
assign x_39196 = x_7901 & x_39195;
assign x_39197 = x_7904 & x_7905;
assign x_39198 = x_7906 & x_7907;
assign x_39199 = x_39197 & x_39198;
assign x_39200 = x_39196 & x_39199;
assign x_39201 = x_7908 & x_7909;
assign x_39202 = x_7910 & x_7911;
assign x_39203 = x_39201 & x_39202;
assign x_39204 = x_7912 & x_7913;
assign x_39205 = x_7914 & x_7915;
assign x_39206 = x_39204 & x_39205;
assign x_39207 = x_39203 & x_39206;
assign x_39208 = x_39200 & x_39207;
assign x_39209 = x_39194 & x_39208;
assign x_39210 = x_7917 & x_7918;
assign x_39211 = x_7916 & x_39210;
assign x_39212 = x_7919 & x_7920;
assign x_39213 = x_7921 & x_7922;
assign x_39214 = x_39212 & x_39213;
assign x_39215 = x_39211 & x_39214;
assign x_39216 = x_7923 & x_7924;
assign x_39217 = x_7925 & x_7926;
assign x_39218 = x_39216 & x_39217;
assign x_39219 = x_7927 & x_7928;
assign x_39220 = x_7929 & x_7930;
assign x_39221 = x_39219 & x_39220;
assign x_39222 = x_39218 & x_39221;
assign x_39223 = x_39215 & x_39222;
assign x_39224 = x_7931 & x_7932;
assign x_39225 = x_7933 & x_7934;
assign x_39226 = x_39224 & x_39225;
assign x_39227 = x_7935 & x_7936;
assign x_39228 = x_7937 & x_7938;
assign x_39229 = x_39227 & x_39228;
assign x_39230 = x_39226 & x_39229;
assign x_39231 = x_7939 & x_7940;
assign x_39232 = x_7941 & x_7942;
assign x_39233 = x_39231 & x_39232;
assign x_39234 = x_7943 & x_7944;
assign x_39235 = x_7945 & x_7946;
assign x_39236 = x_39234 & x_39235;
assign x_39237 = x_39233 & x_39236;
assign x_39238 = x_39230 & x_39237;
assign x_39239 = x_39223 & x_39238;
assign x_39240 = x_39209 & x_39239;
assign x_39241 = x_39180 & x_39240;
assign x_39242 = x_7948 & x_7949;
assign x_39243 = x_7947 & x_39242;
assign x_39244 = x_7950 & x_7951;
assign x_39245 = x_7952 & x_7953;
assign x_39246 = x_39244 & x_39245;
assign x_39247 = x_39243 & x_39246;
assign x_39248 = x_7954 & x_7955;
assign x_39249 = x_7956 & x_7957;
assign x_39250 = x_39248 & x_39249;
assign x_39251 = x_7958 & x_7959;
assign x_39252 = x_7960 & x_7961;
assign x_39253 = x_39251 & x_39252;
assign x_39254 = x_39250 & x_39253;
assign x_39255 = x_39247 & x_39254;
assign x_39256 = x_7963 & x_7964;
assign x_39257 = x_7962 & x_39256;
assign x_39258 = x_7965 & x_7966;
assign x_39259 = x_7967 & x_7968;
assign x_39260 = x_39258 & x_39259;
assign x_39261 = x_39257 & x_39260;
assign x_39262 = x_7969 & x_7970;
assign x_39263 = x_7971 & x_7972;
assign x_39264 = x_39262 & x_39263;
assign x_39265 = x_7973 & x_7974;
assign x_39266 = x_7975 & x_7976;
assign x_39267 = x_39265 & x_39266;
assign x_39268 = x_39264 & x_39267;
assign x_39269 = x_39261 & x_39268;
assign x_39270 = x_39255 & x_39269;
assign x_39271 = x_7978 & x_7979;
assign x_39272 = x_7977 & x_39271;
assign x_39273 = x_7980 & x_7981;
assign x_39274 = x_7982 & x_7983;
assign x_39275 = x_39273 & x_39274;
assign x_39276 = x_39272 & x_39275;
assign x_39277 = x_7984 & x_7985;
assign x_39278 = x_7986 & x_7987;
assign x_39279 = x_39277 & x_39278;
assign x_39280 = x_7988 & x_7989;
assign x_39281 = x_7990 & x_7991;
assign x_39282 = x_39280 & x_39281;
assign x_39283 = x_39279 & x_39282;
assign x_39284 = x_39276 & x_39283;
assign x_39285 = x_7992 & x_7993;
assign x_39286 = x_7994 & x_7995;
assign x_39287 = x_39285 & x_39286;
assign x_39288 = x_7996 & x_7997;
assign x_39289 = x_7998 & x_7999;
assign x_39290 = x_39288 & x_39289;
assign x_39291 = x_39287 & x_39290;
assign x_39292 = x_8000 & x_8001;
assign x_39293 = x_8002 & x_8003;
assign x_39294 = x_39292 & x_39293;
assign x_39295 = x_8004 & x_8005;
assign x_39296 = x_8006 & x_8007;
assign x_39297 = x_39295 & x_39296;
assign x_39298 = x_39294 & x_39297;
assign x_39299 = x_39291 & x_39298;
assign x_39300 = x_39284 & x_39299;
assign x_39301 = x_39270 & x_39300;
assign x_39302 = x_8009 & x_8010;
assign x_39303 = x_8008 & x_39302;
assign x_39304 = x_8011 & x_8012;
assign x_39305 = x_8013 & x_8014;
assign x_39306 = x_39304 & x_39305;
assign x_39307 = x_39303 & x_39306;
assign x_39308 = x_8015 & x_8016;
assign x_39309 = x_8017 & x_8018;
assign x_39310 = x_39308 & x_39309;
assign x_39311 = x_8019 & x_8020;
assign x_39312 = x_8021 & x_8022;
assign x_39313 = x_39311 & x_39312;
assign x_39314 = x_39310 & x_39313;
assign x_39315 = x_39307 & x_39314;
assign x_39316 = x_8024 & x_8025;
assign x_39317 = x_8023 & x_39316;
assign x_39318 = x_8026 & x_8027;
assign x_39319 = x_8028 & x_8029;
assign x_39320 = x_39318 & x_39319;
assign x_39321 = x_39317 & x_39320;
assign x_39322 = x_8030 & x_8031;
assign x_39323 = x_8032 & x_8033;
assign x_39324 = x_39322 & x_39323;
assign x_39325 = x_8034 & x_8035;
assign x_39326 = x_8036 & x_8037;
assign x_39327 = x_39325 & x_39326;
assign x_39328 = x_39324 & x_39327;
assign x_39329 = x_39321 & x_39328;
assign x_39330 = x_39315 & x_39329;
assign x_39331 = x_8039 & x_8040;
assign x_39332 = x_8038 & x_39331;
assign x_39333 = x_8041 & x_8042;
assign x_39334 = x_8043 & x_8044;
assign x_39335 = x_39333 & x_39334;
assign x_39336 = x_39332 & x_39335;
assign x_39337 = x_8045 & x_8046;
assign x_39338 = x_8047 & x_8048;
assign x_39339 = x_39337 & x_39338;
assign x_39340 = x_8049 & x_8050;
assign x_39341 = x_8051 & x_8052;
assign x_39342 = x_39340 & x_39341;
assign x_39343 = x_39339 & x_39342;
assign x_39344 = x_39336 & x_39343;
assign x_39345 = x_8053 & x_8054;
assign x_39346 = x_8055 & x_8056;
assign x_39347 = x_39345 & x_39346;
assign x_39348 = x_8057 & x_8058;
assign x_39349 = x_8059 & x_8060;
assign x_39350 = x_39348 & x_39349;
assign x_39351 = x_39347 & x_39350;
assign x_39352 = x_8061 & x_8062;
assign x_39353 = x_8063 & x_8064;
assign x_39354 = x_39352 & x_39353;
assign x_39355 = x_8065 & x_8066;
assign x_39356 = x_8067 & x_8068;
assign x_39357 = x_39355 & x_39356;
assign x_39358 = x_39354 & x_39357;
assign x_39359 = x_39351 & x_39358;
assign x_39360 = x_39344 & x_39359;
assign x_39361 = x_39330 & x_39360;
assign x_39362 = x_39301 & x_39361;
assign x_39363 = x_39241 & x_39362;
assign x_39364 = x_8070 & x_8071;
assign x_39365 = x_8069 & x_39364;
assign x_39366 = x_8072 & x_8073;
assign x_39367 = x_8074 & x_8075;
assign x_39368 = x_39366 & x_39367;
assign x_39369 = x_39365 & x_39368;
assign x_39370 = x_8076 & x_8077;
assign x_39371 = x_8078 & x_8079;
assign x_39372 = x_39370 & x_39371;
assign x_39373 = x_8080 & x_8081;
assign x_39374 = x_8082 & x_8083;
assign x_39375 = x_39373 & x_39374;
assign x_39376 = x_39372 & x_39375;
assign x_39377 = x_39369 & x_39376;
assign x_39378 = x_8085 & x_8086;
assign x_39379 = x_8084 & x_39378;
assign x_39380 = x_8087 & x_8088;
assign x_39381 = x_8089 & x_8090;
assign x_39382 = x_39380 & x_39381;
assign x_39383 = x_39379 & x_39382;
assign x_39384 = x_8091 & x_8092;
assign x_39385 = x_8093 & x_8094;
assign x_39386 = x_39384 & x_39385;
assign x_39387 = x_8095 & x_8096;
assign x_39388 = x_8097 & x_8098;
assign x_39389 = x_39387 & x_39388;
assign x_39390 = x_39386 & x_39389;
assign x_39391 = x_39383 & x_39390;
assign x_39392 = x_39377 & x_39391;
assign x_39393 = x_8100 & x_8101;
assign x_39394 = x_8099 & x_39393;
assign x_39395 = x_8102 & x_8103;
assign x_39396 = x_8104 & x_8105;
assign x_39397 = x_39395 & x_39396;
assign x_39398 = x_39394 & x_39397;
assign x_39399 = x_8106 & x_8107;
assign x_39400 = x_8108 & x_8109;
assign x_39401 = x_39399 & x_39400;
assign x_39402 = x_8110 & x_8111;
assign x_39403 = x_8112 & x_8113;
assign x_39404 = x_39402 & x_39403;
assign x_39405 = x_39401 & x_39404;
assign x_39406 = x_39398 & x_39405;
assign x_39407 = x_8114 & x_8115;
assign x_39408 = x_8116 & x_8117;
assign x_39409 = x_39407 & x_39408;
assign x_39410 = x_8118 & x_8119;
assign x_39411 = x_8120 & x_8121;
assign x_39412 = x_39410 & x_39411;
assign x_39413 = x_39409 & x_39412;
assign x_39414 = x_8122 & x_8123;
assign x_39415 = x_8124 & x_8125;
assign x_39416 = x_39414 & x_39415;
assign x_39417 = x_8126 & x_8127;
assign x_39418 = x_8128 & x_8129;
assign x_39419 = x_39417 & x_39418;
assign x_39420 = x_39416 & x_39419;
assign x_39421 = x_39413 & x_39420;
assign x_39422 = x_39406 & x_39421;
assign x_39423 = x_39392 & x_39422;
assign x_39424 = x_8131 & x_8132;
assign x_39425 = x_8130 & x_39424;
assign x_39426 = x_8133 & x_8134;
assign x_39427 = x_8135 & x_8136;
assign x_39428 = x_39426 & x_39427;
assign x_39429 = x_39425 & x_39428;
assign x_39430 = x_8137 & x_8138;
assign x_39431 = x_8139 & x_8140;
assign x_39432 = x_39430 & x_39431;
assign x_39433 = x_8141 & x_8142;
assign x_39434 = x_8143 & x_8144;
assign x_39435 = x_39433 & x_39434;
assign x_39436 = x_39432 & x_39435;
assign x_39437 = x_39429 & x_39436;
assign x_39438 = x_8146 & x_8147;
assign x_39439 = x_8145 & x_39438;
assign x_39440 = x_8148 & x_8149;
assign x_39441 = x_8150 & x_8151;
assign x_39442 = x_39440 & x_39441;
assign x_39443 = x_39439 & x_39442;
assign x_39444 = x_8152 & x_8153;
assign x_39445 = x_8154 & x_8155;
assign x_39446 = x_39444 & x_39445;
assign x_39447 = x_8156 & x_8157;
assign x_39448 = x_8158 & x_8159;
assign x_39449 = x_39447 & x_39448;
assign x_39450 = x_39446 & x_39449;
assign x_39451 = x_39443 & x_39450;
assign x_39452 = x_39437 & x_39451;
assign x_39453 = x_8161 & x_8162;
assign x_39454 = x_8160 & x_39453;
assign x_39455 = x_8163 & x_8164;
assign x_39456 = x_8165 & x_8166;
assign x_39457 = x_39455 & x_39456;
assign x_39458 = x_39454 & x_39457;
assign x_39459 = x_8167 & x_8168;
assign x_39460 = x_8169 & x_8170;
assign x_39461 = x_39459 & x_39460;
assign x_39462 = x_8171 & x_8172;
assign x_39463 = x_8173 & x_8174;
assign x_39464 = x_39462 & x_39463;
assign x_39465 = x_39461 & x_39464;
assign x_39466 = x_39458 & x_39465;
assign x_39467 = x_8175 & x_8176;
assign x_39468 = x_8177 & x_8178;
assign x_39469 = x_39467 & x_39468;
assign x_39470 = x_8179 & x_8180;
assign x_39471 = x_8181 & x_8182;
assign x_39472 = x_39470 & x_39471;
assign x_39473 = x_39469 & x_39472;
assign x_39474 = x_8183 & x_8184;
assign x_39475 = x_8185 & x_8186;
assign x_39476 = x_39474 & x_39475;
assign x_39477 = x_8187 & x_8188;
assign x_39478 = x_8189 & x_8190;
assign x_39479 = x_39477 & x_39478;
assign x_39480 = x_39476 & x_39479;
assign x_39481 = x_39473 & x_39480;
assign x_39482 = x_39466 & x_39481;
assign x_39483 = x_39452 & x_39482;
assign x_39484 = x_39423 & x_39483;
assign x_39485 = x_8192 & x_8193;
assign x_39486 = x_8191 & x_39485;
assign x_39487 = x_8194 & x_8195;
assign x_39488 = x_8196 & x_8197;
assign x_39489 = x_39487 & x_39488;
assign x_39490 = x_39486 & x_39489;
assign x_39491 = x_8198 & x_8199;
assign x_39492 = x_8200 & x_8201;
assign x_39493 = x_39491 & x_39492;
assign x_39494 = x_8202 & x_8203;
assign x_39495 = x_8204 & x_8205;
assign x_39496 = x_39494 & x_39495;
assign x_39497 = x_39493 & x_39496;
assign x_39498 = x_39490 & x_39497;
assign x_39499 = x_8207 & x_8208;
assign x_39500 = x_8206 & x_39499;
assign x_39501 = x_8209 & x_8210;
assign x_39502 = x_8211 & x_8212;
assign x_39503 = x_39501 & x_39502;
assign x_39504 = x_39500 & x_39503;
assign x_39505 = x_8213 & x_8214;
assign x_39506 = x_8215 & x_8216;
assign x_39507 = x_39505 & x_39506;
assign x_39508 = x_8217 & x_8218;
assign x_39509 = x_8219 & x_8220;
assign x_39510 = x_39508 & x_39509;
assign x_39511 = x_39507 & x_39510;
assign x_39512 = x_39504 & x_39511;
assign x_39513 = x_39498 & x_39512;
assign x_39514 = x_8222 & x_8223;
assign x_39515 = x_8221 & x_39514;
assign x_39516 = x_8224 & x_8225;
assign x_39517 = x_8226 & x_8227;
assign x_39518 = x_39516 & x_39517;
assign x_39519 = x_39515 & x_39518;
assign x_39520 = x_8228 & x_8229;
assign x_39521 = x_8230 & x_8231;
assign x_39522 = x_39520 & x_39521;
assign x_39523 = x_8232 & x_8233;
assign x_39524 = x_8234 & x_8235;
assign x_39525 = x_39523 & x_39524;
assign x_39526 = x_39522 & x_39525;
assign x_39527 = x_39519 & x_39526;
assign x_39528 = x_8236 & x_8237;
assign x_39529 = x_8238 & x_8239;
assign x_39530 = x_39528 & x_39529;
assign x_39531 = x_8240 & x_8241;
assign x_39532 = x_8242 & x_8243;
assign x_39533 = x_39531 & x_39532;
assign x_39534 = x_39530 & x_39533;
assign x_39535 = x_8244 & x_8245;
assign x_39536 = x_8246 & x_8247;
assign x_39537 = x_39535 & x_39536;
assign x_39538 = x_8248 & x_8249;
assign x_39539 = x_8250 & x_8251;
assign x_39540 = x_39538 & x_39539;
assign x_39541 = x_39537 & x_39540;
assign x_39542 = x_39534 & x_39541;
assign x_39543 = x_39527 & x_39542;
assign x_39544 = x_39513 & x_39543;
assign x_39545 = x_8253 & x_8254;
assign x_39546 = x_8252 & x_39545;
assign x_39547 = x_8255 & x_8256;
assign x_39548 = x_8257 & x_8258;
assign x_39549 = x_39547 & x_39548;
assign x_39550 = x_39546 & x_39549;
assign x_39551 = x_8259 & x_8260;
assign x_39552 = x_8261 & x_8262;
assign x_39553 = x_39551 & x_39552;
assign x_39554 = x_8263 & x_8264;
assign x_39555 = x_8265 & x_8266;
assign x_39556 = x_39554 & x_39555;
assign x_39557 = x_39553 & x_39556;
assign x_39558 = x_39550 & x_39557;
assign x_39559 = x_8267 & x_8268;
assign x_39560 = x_8269 & x_8270;
assign x_39561 = x_39559 & x_39560;
assign x_39562 = x_8271 & x_8272;
assign x_39563 = x_8273 & x_8274;
assign x_39564 = x_39562 & x_39563;
assign x_39565 = x_39561 & x_39564;
assign x_39566 = x_8275 & x_8276;
assign x_39567 = x_8277 & x_8278;
assign x_39568 = x_39566 & x_39567;
assign x_39569 = x_8279 & x_8280;
assign x_39570 = x_8281 & x_8282;
assign x_39571 = x_39569 & x_39570;
assign x_39572 = x_39568 & x_39571;
assign x_39573 = x_39565 & x_39572;
assign x_39574 = x_39558 & x_39573;
assign x_39575 = x_8284 & x_8285;
assign x_39576 = x_8283 & x_39575;
assign x_39577 = x_8286 & x_8287;
assign x_39578 = x_8288 & x_8289;
assign x_39579 = x_39577 & x_39578;
assign x_39580 = x_39576 & x_39579;
assign x_39581 = x_8290 & x_8291;
assign x_39582 = x_8292 & x_8293;
assign x_39583 = x_39581 & x_39582;
assign x_39584 = x_8294 & x_8295;
assign x_39585 = x_8296 & x_8297;
assign x_39586 = x_39584 & x_39585;
assign x_39587 = x_39583 & x_39586;
assign x_39588 = x_39580 & x_39587;
assign x_39589 = x_8298 & x_8299;
assign x_39590 = x_8300 & x_8301;
assign x_39591 = x_39589 & x_39590;
assign x_39592 = x_8302 & x_8303;
assign x_39593 = x_8304 & x_8305;
assign x_39594 = x_39592 & x_39593;
assign x_39595 = x_39591 & x_39594;
assign x_39596 = x_8306 & x_8307;
assign x_39597 = x_8308 & x_8309;
assign x_39598 = x_39596 & x_39597;
assign x_39599 = x_8310 & x_8311;
assign x_39600 = x_8312 & x_8313;
assign x_39601 = x_39599 & x_39600;
assign x_39602 = x_39598 & x_39601;
assign x_39603 = x_39595 & x_39602;
assign x_39604 = x_39588 & x_39603;
assign x_39605 = x_39574 & x_39604;
assign x_39606 = x_39544 & x_39605;
assign x_39607 = x_39484 & x_39606;
assign x_39608 = x_39363 & x_39607;
assign x_39609 = x_8315 & x_8316;
assign x_39610 = x_8314 & x_39609;
assign x_39611 = x_8317 & x_8318;
assign x_39612 = x_8319 & x_8320;
assign x_39613 = x_39611 & x_39612;
assign x_39614 = x_39610 & x_39613;
assign x_39615 = x_8321 & x_8322;
assign x_39616 = x_8323 & x_8324;
assign x_39617 = x_39615 & x_39616;
assign x_39618 = x_8325 & x_8326;
assign x_39619 = x_8327 & x_8328;
assign x_39620 = x_39618 & x_39619;
assign x_39621 = x_39617 & x_39620;
assign x_39622 = x_39614 & x_39621;
assign x_39623 = x_8330 & x_8331;
assign x_39624 = x_8329 & x_39623;
assign x_39625 = x_8332 & x_8333;
assign x_39626 = x_8334 & x_8335;
assign x_39627 = x_39625 & x_39626;
assign x_39628 = x_39624 & x_39627;
assign x_39629 = x_8336 & x_8337;
assign x_39630 = x_8338 & x_8339;
assign x_39631 = x_39629 & x_39630;
assign x_39632 = x_8340 & x_8341;
assign x_39633 = x_8342 & x_8343;
assign x_39634 = x_39632 & x_39633;
assign x_39635 = x_39631 & x_39634;
assign x_39636 = x_39628 & x_39635;
assign x_39637 = x_39622 & x_39636;
assign x_39638 = x_8345 & x_8346;
assign x_39639 = x_8344 & x_39638;
assign x_39640 = x_8347 & x_8348;
assign x_39641 = x_8349 & x_8350;
assign x_39642 = x_39640 & x_39641;
assign x_39643 = x_39639 & x_39642;
assign x_39644 = x_8351 & x_8352;
assign x_39645 = x_8353 & x_8354;
assign x_39646 = x_39644 & x_39645;
assign x_39647 = x_8355 & x_8356;
assign x_39648 = x_8357 & x_8358;
assign x_39649 = x_39647 & x_39648;
assign x_39650 = x_39646 & x_39649;
assign x_39651 = x_39643 & x_39650;
assign x_39652 = x_8359 & x_8360;
assign x_39653 = x_8361 & x_8362;
assign x_39654 = x_39652 & x_39653;
assign x_39655 = x_8363 & x_8364;
assign x_39656 = x_8365 & x_8366;
assign x_39657 = x_39655 & x_39656;
assign x_39658 = x_39654 & x_39657;
assign x_39659 = x_8367 & x_8368;
assign x_39660 = x_8369 & x_8370;
assign x_39661 = x_39659 & x_39660;
assign x_39662 = x_8371 & x_8372;
assign x_39663 = x_8373 & x_8374;
assign x_39664 = x_39662 & x_39663;
assign x_39665 = x_39661 & x_39664;
assign x_39666 = x_39658 & x_39665;
assign x_39667 = x_39651 & x_39666;
assign x_39668 = x_39637 & x_39667;
assign x_39669 = x_8376 & x_8377;
assign x_39670 = x_8375 & x_39669;
assign x_39671 = x_8378 & x_8379;
assign x_39672 = x_8380 & x_8381;
assign x_39673 = x_39671 & x_39672;
assign x_39674 = x_39670 & x_39673;
assign x_39675 = x_8382 & x_8383;
assign x_39676 = x_8384 & x_8385;
assign x_39677 = x_39675 & x_39676;
assign x_39678 = x_8386 & x_8387;
assign x_39679 = x_8388 & x_8389;
assign x_39680 = x_39678 & x_39679;
assign x_39681 = x_39677 & x_39680;
assign x_39682 = x_39674 & x_39681;
assign x_39683 = x_8391 & x_8392;
assign x_39684 = x_8390 & x_39683;
assign x_39685 = x_8393 & x_8394;
assign x_39686 = x_8395 & x_8396;
assign x_39687 = x_39685 & x_39686;
assign x_39688 = x_39684 & x_39687;
assign x_39689 = x_8397 & x_8398;
assign x_39690 = x_8399 & x_8400;
assign x_39691 = x_39689 & x_39690;
assign x_39692 = x_8401 & x_8402;
assign x_39693 = x_8403 & x_8404;
assign x_39694 = x_39692 & x_39693;
assign x_39695 = x_39691 & x_39694;
assign x_39696 = x_39688 & x_39695;
assign x_39697 = x_39682 & x_39696;
assign x_39698 = x_8406 & x_8407;
assign x_39699 = x_8405 & x_39698;
assign x_39700 = x_8408 & x_8409;
assign x_39701 = x_8410 & x_8411;
assign x_39702 = x_39700 & x_39701;
assign x_39703 = x_39699 & x_39702;
assign x_39704 = x_8412 & x_8413;
assign x_39705 = x_8414 & x_8415;
assign x_39706 = x_39704 & x_39705;
assign x_39707 = x_8416 & x_8417;
assign x_39708 = x_8418 & x_8419;
assign x_39709 = x_39707 & x_39708;
assign x_39710 = x_39706 & x_39709;
assign x_39711 = x_39703 & x_39710;
assign x_39712 = x_8420 & x_8421;
assign x_39713 = x_8422 & x_8423;
assign x_39714 = x_39712 & x_39713;
assign x_39715 = x_8424 & x_8425;
assign x_39716 = x_8426 & x_8427;
assign x_39717 = x_39715 & x_39716;
assign x_39718 = x_39714 & x_39717;
assign x_39719 = x_8428 & x_8429;
assign x_39720 = x_8430 & x_8431;
assign x_39721 = x_39719 & x_39720;
assign x_39722 = x_8432 & x_8433;
assign x_39723 = x_8434 & x_8435;
assign x_39724 = x_39722 & x_39723;
assign x_39725 = x_39721 & x_39724;
assign x_39726 = x_39718 & x_39725;
assign x_39727 = x_39711 & x_39726;
assign x_39728 = x_39697 & x_39727;
assign x_39729 = x_39668 & x_39728;
assign x_39730 = x_8437 & x_8438;
assign x_39731 = x_8436 & x_39730;
assign x_39732 = x_8439 & x_8440;
assign x_39733 = x_8441 & x_8442;
assign x_39734 = x_39732 & x_39733;
assign x_39735 = x_39731 & x_39734;
assign x_39736 = x_8443 & x_8444;
assign x_39737 = x_8445 & x_8446;
assign x_39738 = x_39736 & x_39737;
assign x_39739 = x_8447 & x_8448;
assign x_39740 = x_8449 & x_8450;
assign x_39741 = x_39739 & x_39740;
assign x_39742 = x_39738 & x_39741;
assign x_39743 = x_39735 & x_39742;
assign x_39744 = x_8452 & x_8453;
assign x_39745 = x_8451 & x_39744;
assign x_39746 = x_8454 & x_8455;
assign x_39747 = x_8456 & x_8457;
assign x_39748 = x_39746 & x_39747;
assign x_39749 = x_39745 & x_39748;
assign x_39750 = x_8458 & x_8459;
assign x_39751 = x_8460 & x_8461;
assign x_39752 = x_39750 & x_39751;
assign x_39753 = x_8462 & x_8463;
assign x_39754 = x_8464 & x_8465;
assign x_39755 = x_39753 & x_39754;
assign x_39756 = x_39752 & x_39755;
assign x_39757 = x_39749 & x_39756;
assign x_39758 = x_39743 & x_39757;
assign x_39759 = x_8467 & x_8468;
assign x_39760 = x_8466 & x_39759;
assign x_39761 = x_8469 & x_8470;
assign x_39762 = x_8471 & x_8472;
assign x_39763 = x_39761 & x_39762;
assign x_39764 = x_39760 & x_39763;
assign x_39765 = x_8473 & x_8474;
assign x_39766 = x_8475 & x_8476;
assign x_39767 = x_39765 & x_39766;
assign x_39768 = x_8477 & x_8478;
assign x_39769 = x_8479 & x_8480;
assign x_39770 = x_39768 & x_39769;
assign x_39771 = x_39767 & x_39770;
assign x_39772 = x_39764 & x_39771;
assign x_39773 = x_8481 & x_8482;
assign x_39774 = x_8483 & x_8484;
assign x_39775 = x_39773 & x_39774;
assign x_39776 = x_8485 & x_8486;
assign x_39777 = x_8487 & x_8488;
assign x_39778 = x_39776 & x_39777;
assign x_39779 = x_39775 & x_39778;
assign x_39780 = x_8489 & x_8490;
assign x_39781 = x_8491 & x_8492;
assign x_39782 = x_39780 & x_39781;
assign x_39783 = x_8493 & x_8494;
assign x_39784 = x_8495 & x_8496;
assign x_39785 = x_39783 & x_39784;
assign x_39786 = x_39782 & x_39785;
assign x_39787 = x_39779 & x_39786;
assign x_39788 = x_39772 & x_39787;
assign x_39789 = x_39758 & x_39788;
assign x_39790 = x_8498 & x_8499;
assign x_39791 = x_8497 & x_39790;
assign x_39792 = x_8500 & x_8501;
assign x_39793 = x_8502 & x_8503;
assign x_39794 = x_39792 & x_39793;
assign x_39795 = x_39791 & x_39794;
assign x_39796 = x_8504 & x_8505;
assign x_39797 = x_8506 & x_8507;
assign x_39798 = x_39796 & x_39797;
assign x_39799 = x_8508 & x_8509;
assign x_39800 = x_8510 & x_8511;
assign x_39801 = x_39799 & x_39800;
assign x_39802 = x_39798 & x_39801;
assign x_39803 = x_39795 & x_39802;
assign x_39804 = x_8513 & x_8514;
assign x_39805 = x_8512 & x_39804;
assign x_39806 = x_8515 & x_8516;
assign x_39807 = x_8517 & x_8518;
assign x_39808 = x_39806 & x_39807;
assign x_39809 = x_39805 & x_39808;
assign x_39810 = x_8519 & x_8520;
assign x_39811 = x_8521 & x_8522;
assign x_39812 = x_39810 & x_39811;
assign x_39813 = x_8523 & x_8524;
assign x_39814 = x_8525 & x_8526;
assign x_39815 = x_39813 & x_39814;
assign x_39816 = x_39812 & x_39815;
assign x_39817 = x_39809 & x_39816;
assign x_39818 = x_39803 & x_39817;
assign x_39819 = x_8528 & x_8529;
assign x_39820 = x_8527 & x_39819;
assign x_39821 = x_8530 & x_8531;
assign x_39822 = x_8532 & x_8533;
assign x_39823 = x_39821 & x_39822;
assign x_39824 = x_39820 & x_39823;
assign x_39825 = x_8534 & x_8535;
assign x_39826 = x_8536 & x_8537;
assign x_39827 = x_39825 & x_39826;
assign x_39828 = x_8538 & x_8539;
assign x_39829 = x_8540 & x_8541;
assign x_39830 = x_39828 & x_39829;
assign x_39831 = x_39827 & x_39830;
assign x_39832 = x_39824 & x_39831;
assign x_39833 = x_8542 & x_8543;
assign x_39834 = x_8544 & x_8545;
assign x_39835 = x_39833 & x_39834;
assign x_39836 = x_8546 & x_8547;
assign x_39837 = x_8548 & x_8549;
assign x_39838 = x_39836 & x_39837;
assign x_39839 = x_39835 & x_39838;
assign x_39840 = x_8550 & x_8551;
assign x_39841 = x_8552 & x_8553;
assign x_39842 = x_39840 & x_39841;
assign x_39843 = x_8554 & x_8555;
assign x_39844 = x_8556 & x_8557;
assign x_39845 = x_39843 & x_39844;
assign x_39846 = x_39842 & x_39845;
assign x_39847 = x_39839 & x_39846;
assign x_39848 = x_39832 & x_39847;
assign x_39849 = x_39818 & x_39848;
assign x_39850 = x_39789 & x_39849;
assign x_39851 = x_39729 & x_39850;
assign x_39852 = x_8559 & x_8560;
assign x_39853 = x_8558 & x_39852;
assign x_39854 = x_8561 & x_8562;
assign x_39855 = x_8563 & x_8564;
assign x_39856 = x_39854 & x_39855;
assign x_39857 = x_39853 & x_39856;
assign x_39858 = x_8565 & x_8566;
assign x_39859 = x_8567 & x_8568;
assign x_39860 = x_39858 & x_39859;
assign x_39861 = x_8569 & x_8570;
assign x_39862 = x_8571 & x_8572;
assign x_39863 = x_39861 & x_39862;
assign x_39864 = x_39860 & x_39863;
assign x_39865 = x_39857 & x_39864;
assign x_39866 = x_8574 & x_8575;
assign x_39867 = x_8573 & x_39866;
assign x_39868 = x_8576 & x_8577;
assign x_39869 = x_8578 & x_8579;
assign x_39870 = x_39868 & x_39869;
assign x_39871 = x_39867 & x_39870;
assign x_39872 = x_8580 & x_8581;
assign x_39873 = x_8582 & x_8583;
assign x_39874 = x_39872 & x_39873;
assign x_39875 = x_8584 & x_8585;
assign x_39876 = x_8586 & x_8587;
assign x_39877 = x_39875 & x_39876;
assign x_39878 = x_39874 & x_39877;
assign x_39879 = x_39871 & x_39878;
assign x_39880 = x_39865 & x_39879;
assign x_39881 = x_8589 & x_8590;
assign x_39882 = x_8588 & x_39881;
assign x_39883 = x_8591 & x_8592;
assign x_39884 = x_8593 & x_8594;
assign x_39885 = x_39883 & x_39884;
assign x_39886 = x_39882 & x_39885;
assign x_39887 = x_8595 & x_8596;
assign x_39888 = x_8597 & x_8598;
assign x_39889 = x_39887 & x_39888;
assign x_39890 = x_8599 & x_8600;
assign x_39891 = x_8601 & x_8602;
assign x_39892 = x_39890 & x_39891;
assign x_39893 = x_39889 & x_39892;
assign x_39894 = x_39886 & x_39893;
assign x_39895 = x_8603 & x_8604;
assign x_39896 = x_8605 & x_8606;
assign x_39897 = x_39895 & x_39896;
assign x_39898 = x_8607 & x_8608;
assign x_39899 = x_8609 & x_8610;
assign x_39900 = x_39898 & x_39899;
assign x_39901 = x_39897 & x_39900;
assign x_39902 = x_8611 & x_8612;
assign x_39903 = x_8613 & x_8614;
assign x_39904 = x_39902 & x_39903;
assign x_39905 = x_8615 & x_8616;
assign x_39906 = x_8617 & x_8618;
assign x_39907 = x_39905 & x_39906;
assign x_39908 = x_39904 & x_39907;
assign x_39909 = x_39901 & x_39908;
assign x_39910 = x_39894 & x_39909;
assign x_39911 = x_39880 & x_39910;
assign x_39912 = x_8620 & x_8621;
assign x_39913 = x_8619 & x_39912;
assign x_39914 = x_8622 & x_8623;
assign x_39915 = x_8624 & x_8625;
assign x_39916 = x_39914 & x_39915;
assign x_39917 = x_39913 & x_39916;
assign x_39918 = x_8626 & x_8627;
assign x_39919 = x_8628 & x_8629;
assign x_39920 = x_39918 & x_39919;
assign x_39921 = x_8630 & x_8631;
assign x_39922 = x_8632 & x_8633;
assign x_39923 = x_39921 & x_39922;
assign x_39924 = x_39920 & x_39923;
assign x_39925 = x_39917 & x_39924;
assign x_39926 = x_8635 & x_8636;
assign x_39927 = x_8634 & x_39926;
assign x_39928 = x_8637 & x_8638;
assign x_39929 = x_8639 & x_8640;
assign x_39930 = x_39928 & x_39929;
assign x_39931 = x_39927 & x_39930;
assign x_39932 = x_8641 & x_8642;
assign x_39933 = x_8643 & x_8644;
assign x_39934 = x_39932 & x_39933;
assign x_39935 = x_8645 & x_8646;
assign x_39936 = x_8647 & x_8648;
assign x_39937 = x_39935 & x_39936;
assign x_39938 = x_39934 & x_39937;
assign x_39939 = x_39931 & x_39938;
assign x_39940 = x_39925 & x_39939;
assign x_39941 = x_8650 & x_8651;
assign x_39942 = x_8649 & x_39941;
assign x_39943 = x_8652 & x_8653;
assign x_39944 = x_8654 & x_8655;
assign x_39945 = x_39943 & x_39944;
assign x_39946 = x_39942 & x_39945;
assign x_39947 = x_8656 & x_8657;
assign x_39948 = x_8658 & x_8659;
assign x_39949 = x_39947 & x_39948;
assign x_39950 = x_8660 & x_8661;
assign x_39951 = x_8662 & x_8663;
assign x_39952 = x_39950 & x_39951;
assign x_39953 = x_39949 & x_39952;
assign x_39954 = x_39946 & x_39953;
assign x_39955 = x_8664 & x_8665;
assign x_39956 = x_8666 & x_8667;
assign x_39957 = x_39955 & x_39956;
assign x_39958 = x_8668 & x_8669;
assign x_39959 = x_8670 & x_8671;
assign x_39960 = x_39958 & x_39959;
assign x_39961 = x_39957 & x_39960;
assign x_39962 = x_8672 & x_8673;
assign x_39963 = x_8674 & x_8675;
assign x_39964 = x_39962 & x_39963;
assign x_39965 = x_8676 & x_8677;
assign x_39966 = x_8678 & x_8679;
assign x_39967 = x_39965 & x_39966;
assign x_39968 = x_39964 & x_39967;
assign x_39969 = x_39961 & x_39968;
assign x_39970 = x_39954 & x_39969;
assign x_39971 = x_39940 & x_39970;
assign x_39972 = x_39911 & x_39971;
assign x_39973 = x_8681 & x_8682;
assign x_39974 = x_8680 & x_39973;
assign x_39975 = x_8683 & x_8684;
assign x_39976 = x_8685 & x_8686;
assign x_39977 = x_39975 & x_39976;
assign x_39978 = x_39974 & x_39977;
assign x_39979 = x_8687 & x_8688;
assign x_39980 = x_8689 & x_8690;
assign x_39981 = x_39979 & x_39980;
assign x_39982 = x_8691 & x_8692;
assign x_39983 = x_8693 & x_8694;
assign x_39984 = x_39982 & x_39983;
assign x_39985 = x_39981 & x_39984;
assign x_39986 = x_39978 & x_39985;
assign x_39987 = x_8696 & x_8697;
assign x_39988 = x_8695 & x_39987;
assign x_39989 = x_8698 & x_8699;
assign x_39990 = x_8700 & x_8701;
assign x_39991 = x_39989 & x_39990;
assign x_39992 = x_39988 & x_39991;
assign x_39993 = x_8702 & x_8703;
assign x_39994 = x_8704 & x_8705;
assign x_39995 = x_39993 & x_39994;
assign x_39996 = x_8706 & x_8707;
assign x_39997 = x_8708 & x_8709;
assign x_39998 = x_39996 & x_39997;
assign x_39999 = x_39995 & x_39998;
assign x_40000 = x_39992 & x_39999;
assign x_40001 = x_39986 & x_40000;
assign x_40002 = x_8711 & x_8712;
assign x_40003 = x_8710 & x_40002;
assign x_40004 = x_8713 & x_8714;
assign x_40005 = x_8715 & x_8716;
assign x_40006 = x_40004 & x_40005;
assign x_40007 = x_40003 & x_40006;
assign x_40008 = x_8717 & x_8718;
assign x_40009 = x_8719 & x_8720;
assign x_40010 = x_40008 & x_40009;
assign x_40011 = x_8721 & x_8722;
assign x_40012 = x_8723 & x_8724;
assign x_40013 = x_40011 & x_40012;
assign x_40014 = x_40010 & x_40013;
assign x_40015 = x_40007 & x_40014;
assign x_40016 = x_8725 & x_8726;
assign x_40017 = x_8727 & x_8728;
assign x_40018 = x_40016 & x_40017;
assign x_40019 = x_8729 & x_8730;
assign x_40020 = x_8731 & x_8732;
assign x_40021 = x_40019 & x_40020;
assign x_40022 = x_40018 & x_40021;
assign x_40023 = x_8733 & x_8734;
assign x_40024 = x_8735 & x_8736;
assign x_40025 = x_40023 & x_40024;
assign x_40026 = x_8737 & x_8738;
assign x_40027 = x_8739 & x_8740;
assign x_40028 = x_40026 & x_40027;
assign x_40029 = x_40025 & x_40028;
assign x_40030 = x_40022 & x_40029;
assign x_40031 = x_40015 & x_40030;
assign x_40032 = x_40001 & x_40031;
assign x_40033 = x_8742 & x_8743;
assign x_40034 = x_8741 & x_40033;
assign x_40035 = x_8744 & x_8745;
assign x_40036 = x_8746 & x_8747;
assign x_40037 = x_40035 & x_40036;
assign x_40038 = x_40034 & x_40037;
assign x_40039 = x_8748 & x_8749;
assign x_40040 = x_8750 & x_8751;
assign x_40041 = x_40039 & x_40040;
assign x_40042 = x_8752 & x_8753;
assign x_40043 = x_8754 & x_8755;
assign x_40044 = x_40042 & x_40043;
assign x_40045 = x_40041 & x_40044;
assign x_40046 = x_40038 & x_40045;
assign x_40047 = x_8756 & x_8757;
assign x_40048 = x_8758 & x_8759;
assign x_40049 = x_40047 & x_40048;
assign x_40050 = x_8760 & x_8761;
assign x_40051 = x_8762 & x_8763;
assign x_40052 = x_40050 & x_40051;
assign x_40053 = x_40049 & x_40052;
assign x_40054 = x_8764 & x_8765;
assign x_40055 = x_8766 & x_8767;
assign x_40056 = x_40054 & x_40055;
assign x_40057 = x_8768 & x_8769;
assign x_40058 = x_8770 & x_8771;
assign x_40059 = x_40057 & x_40058;
assign x_40060 = x_40056 & x_40059;
assign x_40061 = x_40053 & x_40060;
assign x_40062 = x_40046 & x_40061;
assign x_40063 = x_8773 & x_8774;
assign x_40064 = x_8772 & x_40063;
assign x_40065 = x_8775 & x_8776;
assign x_40066 = x_8777 & x_8778;
assign x_40067 = x_40065 & x_40066;
assign x_40068 = x_40064 & x_40067;
assign x_40069 = x_8779 & x_8780;
assign x_40070 = x_8781 & x_8782;
assign x_40071 = x_40069 & x_40070;
assign x_40072 = x_8783 & x_8784;
assign x_40073 = x_8785 & x_8786;
assign x_40074 = x_40072 & x_40073;
assign x_40075 = x_40071 & x_40074;
assign x_40076 = x_40068 & x_40075;
assign x_40077 = x_8787 & x_8788;
assign x_40078 = x_8789 & x_8790;
assign x_40079 = x_40077 & x_40078;
assign x_40080 = x_8791 & x_8792;
assign x_40081 = x_8793 & x_8794;
assign x_40082 = x_40080 & x_40081;
assign x_40083 = x_40079 & x_40082;
assign x_40084 = x_8795 & x_8796;
assign x_40085 = x_8797 & x_8798;
assign x_40086 = x_40084 & x_40085;
assign x_40087 = x_8799 & x_8800;
assign x_40088 = x_8801 & x_8802;
assign x_40089 = x_40087 & x_40088;
assign x_40090 = x_40086 & x_40089;
assign x_40091 = x_40083 & x_40090;
assign x_40092 = x_40076 & x_40091;
assign x_40093 = x_40062 & x_40092;
assign x_40094 = x_40032 & x_40093;
assign x_40095 = x_39972 & x_40094;
assign x_40096 = x_39851 & x_40095;
assign x_40097 = x_39608 & x_40096;
assign x_40098 = x_8804 & x_8805;
assign x_40099 = x_8803 & x_40098;
assign x_40100 = x_8806 & x_8807;
assign x_40101 = x_8808 & x_8809;
assign x_40102 = x_40100 & x_40101;
assign x_40103 = x_40099 & x_40102;
assign x_40104 = x_8810 & x_8811;
assign x_40105 = x_8812 & x_8813;
assign x_40106 = x_40104 & x_40105;
assign x_40107 = x_8814 & x_8815;
assign x_40108 = x_8816 & x_8817;
assign x_40109 = x_40107 & x_40108;
assign x_40110 = x_40106 & x_40109;
assign x_40111 = x_40103 & x_40110;
assign x_40112 = x_8819 & x_8820;
assign x_40113 = x_8818 & x_40112;
assign x_40114 = x_8821 & x_8822;
assign x_40115 = x_8823 & x_8824;
assign x_40116 = x_40114 & x_40115;
assign x_40117 = x_40113 & x_40116;
assign x_40118 = x_8825 & x_8826;
assign x_40119 = x_8827 & x_8828;
assign x_40120 = x_40118 & x_40119;
assign x_40121 = x_8829 & x_8830;
assign x_40122 = x_8831 & x_8832;
assign x_40123 = x_40121 & x_40122;
assign x_40124 = x_40120 & x_40123;
assign x_40125 = x_40117 & x_40124;
assign x_40126 = x_40111 & x_40125;
assign x_40127 = x_8834 & x_8835;
assign x_40128 = x_8833 & x_40127;
assign x_40129 = x_8836 & x_8837;
assign x_40130 = x_8838 & x_8839;
assign x_40131 = x_40129 & x_40130;
assign x_40132 = x_40128 & x_40131;
assign x_40133 = x_8840 & x_8841;
assign x_40134 = x_8842 & x_8843;
assign x_40135 = x_40133 & x_40134;
assign x_40136 = x_8844 & x_8845;
assign x_40137 = x_8846 & x_8847;
assign x_40138 = x_40136 & x_40137;
assign x_40139 = x_40135 & x_40138;
assign x_40140 = x_40132 & x_40139;
assign x_40141 = x_8848 & x_8849;
assign x_40142 = x_8850 & x_8851;
assign x_40143 = x_40141 & x_40142;
assign x_40144 = x_8852 & x_8853;
assign x_40145 = x_8854 & x_8855;
assign x_40146 = x_40144 & x_40145;
assign x_40147 = x_40143 & x_40146;
assign x_40148 = x_8856 & x_8857;
assign x_40149 = x_8858 & x_8859;
assign x_40150 = x_40148 & x_40149;
assign x_40151 = x_8860 & x_8861;
assign x_40152 = x_8862 & x_8863;
assign x_40153 = x_40151 & x_40152;
assign x_40154 = x_40150 & x_40153;
assign x_40155 = x_40147 & x_40154;
assign x_40156 = x_40140 & x_40155;
assign x_40157 = x_40126 & x_40156;
assign x_40158 = x_8865 & x_8866;
assign x_40159 = x_8864 & x_40158;
assign x_40160 = x_8867 & x_8868;
assign x_40161 = x_8869 & x_8870;
assign x_40162 = x_40160 & x_40161;
assign x_40163 = x_40159 & x_40162;
assign x_40164 = x_8871 & x_8872;
assign x_40165 = x_8873 & x_8874;
assign x_40166 = x_40164 & x_40165;
assign x_40167 = x_8875 & x_8876;
assign x_40168 = x_8877 & x_8878;
assign x_40169 = x_40167 & x_40168;
assign x_40170 = x_40166 & x_40169;
assign x_40171 = x_40163 & x_40170;
assign x_40172 = x_8880 & x_8881;
assign x_40173 = x_8879 & x_40172;
assign x_40174 = x_8882 & x_8883;
assign x_40175 = x_8884 & x_8885;
assign x_40176 = x_40174 & x_40175;
assign x_40177 = x_40173 & x_40176;
assign x_40178 = x_8886 & x_8887;
assign x_40179 = x_8888 & x_8889;
assign x_40180 = x_40178 & x_40179;
assign x_40181 = x_8890 & x_8891;
assign x_40182 = x_8892 & x_8893;
assign x_40183 = x_40181 & x_40182;
assign x_40184 = x_40180 & x_40183;
assign x_40185 = x_40177 & x_40184;
assign x_40186 = x_40171 & x_40185;
assign x_40187 = x_8895 & x_8896;
assign x_40188 = x_8894 & x_40187;
assign x_40189 = x_8897 & x_8898;
assign x_40190 = x_8899 & x_8900;
assign x_40191 = x_40189 & x_40190;
assign x_40192 = x_40188 & x_40191;
assign x_40193 = x_8901 & x_8902;
assign x_40194 = x_8903 & x_8904;
assign x_40195 = x_40193 & x_40194;
assign x_40196 = x_8905 & x_8906;
assign x_40197 = x_8907 & x_8908;
assign x_40198 = x_40196 & x_40197;
assign x_40199 = x_40195 & x_40198;
assign x_40200 = x_40192 & x_40199;
assign x_40201 = x_8909 & x_8910;
assign x_40202 = x_8911 & x_8912;
assign x_40203 = x_40201 & x_40202;
assign x_40204 = x_8913 & x_8914;
assign x_40205 = x_8915 & x_8916;
assign x_40206 = x_40204 & x_40205;
assign x_40207 = x_40203 & x_40206;
assign x_40208 = x_8917 & x_8918;
assign x_40209 = x_8919 & x_8920;
assign x_40210 = x_40208 & x_40209;
assign x_40211 = x_8921 & x_8922;
assign x_40212 = x_8923 & x_8924;
assign x_40213 = x_40211 & x_40212;
assign x_40214 = x_40210 & x_40213;
assign x_40215 = x_40207 & x_40214;
assign x_40216 = x_40200 & x_40215;
assign x_40217 = x_40186 & x_40216;
assign x_40218 = x_40157 & x_40217;
assign x_40219 = x_8926 & x_8927;
assign x_40220 = x_8925 & x_40219;
assign x_40221 = x_8928 & x_8929;
assign x_40222 = x_8930 & x_8931;
assign x_40223 = x_40221 & x_40222;
assign x_40224 = x_40220 & x_40223;
assign x_40225 = x_8932 & x_8933;
assign x_40226 = x_8934 & x_8935;
assign x_40227 = x_40225 & x_40226;
assign x_40228 = x_8936 & x_8937;
assign x_40229 = x_8938 & x_8939;
assign x_40230 = x_40228 & x_40229;
assign x_40231 = x_40227 & x_40230;
assign x_40232 = x_40224 & x_40231;
assign x_40233 = x_8941 & x_8942;
assign x_40234 = x_8940 & x_40233;
assign x_40235 = x_8943 & x_8944;
assign x_40236 = x_8945 & x_8946;
assign x_40237 = x_40235 & x_40236;
assign x_40238 = x_40234 & x_40237;
assign x_40239 = x_8947 & x_8948;
assign x_40240 = x_8949 & x_8950;
assign x_40241 = x_40239 & x_40240;
assign x_40242 = x_8951 & x_8952;
assign x_40243 = x_8953 & x_8954;
assign x_40244 = x_40242 & x_40243;
assign x_40245 = x_40241 & x_40244;
assign x_40246 = x_40238 & x_40245;
assign x_40247 = x_40232 & x_40246;
assign x_40248 = x_8956 & x_8957;
assign x_40249 = x_8955 & x_40248;
assign x_40250 = x_8958 & x_8959;
assign x_40251 = x_8960 & x_8961;
assign x_40252 = x_40250 & x_40251;
assign x_40253 = x_40249 & x_40252;
assign x_40254 = x_8962 & x_8963;
assign x_40255 = x_8964 & x_8965;
assign x_40256 = x_40254 & x_40255;
assign x_40257 = x_8966 & x_8967;
assign x_40258 = x_8968 & x_8969;
assign x_40259 = x_40257 & x_40258;
assign x_40260 = x_40256 & x_40259;
assign x_40261 = x_40253 & x_40260;
assign x_40262 = x_8970 & x_8971;
assign x_40263 = x_8972 & x_8973;
assign x_40264 = x_40262 & x_40263;
assign x_40265 = x_8974 & x_8975;
assign x_40266 = x_8976 & x_8977;
assign x_40267 = x_40265 & x_40266;
assign x_40268 = x_40264 & x_40267;
assign x_40269 = x_8978 & x_8979;
assign x_40270 = x_8980 & x_8981;
assign x_40271 = x_40269 & x_40270;
assign x_40272 = x_8982 & x_8983;
assign x_40273 = x_8984 & x_8985;
assign x_40274 = x_40272 & x_40273;
assign x_40275 = x_40271 & x_40274;
assign x_40276 = x_40268 & x_40275;
assign x_40277 = x_40261 & x_40276;
assign x_40278 = x_40247 & x_40277;
assign x_40279 = x_8987 & x_8988;
assign x_40280 = x_8986 & x_40279;
assign x_40281 = x_8989 & x_8990;
assign x_40282 = x_8991 & x_8992;
assign x_40283 = x_40281 & x_40282;
assign x_40284 = x_40280 & x_40283;
assign x_40285 = x_8993 & x_8994;
assign x_40286 = x_8995 & x_8996;
assign x_40287 = x_40285 & x_40286;
assign x_40288 = x_8997 & x_8998;
assign x_40289 = x_8999 & x_9000;
assign x_40290 = x_40288 & x_40289;
assign x_40291 = x_40287 & x_40290;
assign x_40292 = x_40284 & x_40291;
assign x_40293 = x_9002 & x_9003;
assign x_40294 = x_9001 & x_40293;
assign x_40295 = x_9004 & x_9005;
assign x_40296 = x_9006 & x_9007;
assign x_40297 = x_40295 & x_40296;
assign x_40298 = x_40294 & x_40297;
assign x_40299 = x_9008 & x_9009;
assign x_40300 = x_9010 & x_9011;
assign x_40301 = x_40299 & x_40300;
assign x_40302 = x_9012 & x_9013;
assign x_40303 = x_9014 & x_9015;
assign x_40304 = x_40302 & x_40303;
assign x_40305 = x_40301 & x_40304;
assign x_40306 = x_40298 & x_40305;
assign x_40307 = x_40292 & x_40306;
assign x_40308 = x_9017 & x_9018;
assign x_40309 = x_9016 & x_40308;
assign x_40310 = x_9019 & x_9020;
assign x_40311 = x_9021 & x_9022;
assign x_40312 = x_40310 & x_40311;
assign x_40313 = x_40309 & x_40312;
assign x_40314 = x_9023 & x_9024;
assign x_40315 = x_9025 & x_9026;
assign x_40316 = x_40314 & x_40315;
assign x_40317 = x_9027 & x_9028;
assign x_40318 = x_9029 & x_9030;
assign x_40319 = x_40317 & x_40318;
assign x_40320 = x_40316 & x_40319;
assign x_40321 = x_40313 & x_40320;
assign x_40322 = x_9031 & x_9032;
assign x_40323 = x_9033 & x_9034;
assign x_40324 = x_40322 & x_40323;
assign x_40325 = x_9035 & x_9036;
assign x_40326 = x_9037 & x_9038;
assign x_40327 = x_40325 & x_40326;
assign x_40328 = x_40324 & x_40327;
assign x_40329 = x_9039 & x_9040;
assign x_40330 = x_9041 & x_9042;
assign x_40331 = x_40329 & x_40330;
assign x_40332 = x_9043 & x_9044;
assign x_40333 = x_9045 & x_9046;
assign x_40334 = x_40332 & x_40333;
assign x_40335 = x_40331 & x_40334;
assign x_40336 = x_40328 & x_40335;
assign x_40337 = x_40321 & x_40336;
assign x_40338 = x_40307 & x_40337;
assign x_40339 = x_40278 & x_40338;
assign x_40340 = x_40218 & x_40339;
assign x_40341 = x_9048 & x_9049;
assign x_40342 = x_9047 & x_40341;
assign x_40343 = x_9050 & x_9051;
assign x_40344 = x_9052 & x_9053;
assign x_40345 = x_40343 & x_40344;
assign x_40346 = x_40342 & x_40345;
assign x_40347 = x_9054 & x_9055;
assign x_40348 = x_9056 & x_9057;
assign x_40349 = x_40347 & x_40348;
assign x_40350 = x_9058 & x_9059;
assign x_40351 = x_9060 & x_9061;
assign x_40352 = x_40350 & x_40351;
assign x_40353 = x_40349 & x_40352;
assign x_40354 = x_40346 & x_40353;
assign x_40355 = x_9063 & x_9064;
assign x_40356 = x_9062 & x_40355;
assign x_40357 = x_9065 & x_9066;
assign x_40358 = x_9067 & x_9068;
assign x_40359 = x_40357 & x_40358;
assign x_40360 = x_40356 & x_40359;
assign x_40361 = x_9069 & x_9070;
assign x_40362 = x_9071 & x_9072;
assign x_40363 = x_40361 & x_40362;
assign x_40364 = x_9073 & x_9074;
assign x_40365 = x_9075 & x_9076;
assign x_40366 = x_40364 & x_40365;
assign x_40367 = x_40363 & x_40366;
assign x_40368 = x_40360 & x_40367;
assign x_40369 = x_40354 & x_40368;
assign x_40370 = x_9078 & x_9079;
assign x_40371 = x_9077 & x_40370;
assign x_40372 = x_9080 & x_9081;
assign x_40373 = x_9082 & x_9083;
assign x_40374 = x_40372 & x_40373;
assign x_40375 = x_40371 & x_40374;
assign x_40376 = x_9084 & x_9085;
assign x_40377 = x_9086 & x_9087;
assign x_40378 = x_40376 & x_40377;
assign x_40379 = x_9088 & x_9089;
assign x_40380 = x_9090 & x_9091;
assign x_40381 = x_40379 & x_40380;
assign x_40382 = x_40378 & x_40381;
assign x_40383 = x_40375 & x_40382;
assign x_40384 = x_9092 & x_9093;
assign x_40385 = x_9094 & x_9095;
assign x_40386 = x_40384 & x_40385;
assign x_40387 = x_9096 & x_9097;
assign x_40388 = x_9098 & x_9099;
assign x_40389 = x_40387 & x_40388;
assign x_40390 = x_40386 & x_40389;
assign x_40391 = x_9100 & x_9101;
assign x_40392 = x_9102 & x_9103;
assign x_40393 = x_40391 & x_40392;
assign x_40394 = x_9104 & x_9105;
assign x_40395 = x_9106 & x_9107;
assign x_40396 = x_40394 & x_40395;
assign x_40397 = x_40393 & x_40396;
assign x_40398 = x_40390 & x_40397;
assign x_40399 = x_40383 & x_40398;
assign x_40400 = x_40369 & x_40399;
assign x_40401 = x_9109 & x_9110;
assign x_40402 = x_9108 & x_40401;
assign x_40403 = x_9111 & x_9112;
assign x_40404 = x_9113 & x_9114;
assign x_40405 = x_40403 & x_40404;
assign x_40406 = x_40402 & x_40405;
assign x_40407 = x_9115 & x_9116;
assign x_40408 = x_9117 & x_9118;
assign x_40409 = x_40407 & x_40408;
assign x_40410 = x_9119 & x_9120;
assign x_40411 = x_9121 & x_9122;
assign x_40412 = x_40410 & x_40411;
assign x_40413 = x_40409 & x_40412;
assign x_40414 = x_40406 & x_40413;
assign x_40415 = x_9124 & x_9125;
assign x_40416 = x_9123 & x_40415;
assign x_40417 = x_9126 & x_9127;
assign x_40418 = x_9128 & x_9129;
assign x_40419 = x_40417 & x_40418;
assign x_40420 = x_40416 & x_40419;
assign x_40421 = x_9130 & x_9131;
assign x_40422 = x_9132 & x_9133;
assign x_40423 = x_40421 & x_40422;
assign x_40424 = x_9134 & x_9135;
assign x_40425 = x_9136 & x_9137;
assign x_40426 = x_40424 & x_40425;
assign x_40427 = x_40423 & x_40426;
assign x_40428 = x_40420 & x_40427;
assign x_40429 = x_40414 & x_40428;
assign x_40430 = x_9139 & x_9140;
assign x_40431 = x_9138 & x_40430;
assign x_40432 = x_9141 & x_9142;
assign x_40433 = x_9143 & x_9144;
assign x_40434 = x_40432 & x_40433;
assign x_40435 = x_40431 & x_40434;
assign x_40436 = x_9145 & x_9146;
assign x_40437 = x_9147 & x_9148;
assign x_40438 = x_40436 & x_40437;
assign x_40439 = x_9149 & x_9150;
assign x_40440 = x_9151 & x_9152;
assign x_40441 = x_40439 & x_40440;
assign x_40442 = x_40438 & x_40441;
assign x_40443 = x_40435 & x_40442;
assign x_40444 = x_9153 & x_9154;
assign x_40445 = x_9155 & x_9156;
assign x_40446 = x_40444 & x_40445;
assign x_40447 = x_9157 & x_9158;
assign x_40448 = x_9159 & x_9160;
assign x_40449 = x_40447 & x_40448;
assign x_40450 = x_40446 & x_40449;
assign x_40451 = x_9161 & x_9162;
assign x_40452 = x_9163 & x_9164;
assign x_40453 = x_40451 & x_40452;
assign x_40454 = x_9165 & x_9166;
assign x_40455 = x_9167 & x_9168;
assign x_40456 = x_40454 & x_40455;
assign x_40457 = x_40453 & x_40456;
assign x_40458 = x_40450 & x_40457;
assign x_40459 = x_40443 & x_40458;
assign x_40460 = x_40429 & x_40459;
assign x_40461 = x_40400 & x_40460;
assign x_40462 = x_9170 & x_9171;
assign x_40463 = x_9169 & x_40462;
assign x_40464 = x_9172 & x_9173;
assign x_40465 = x_9174 & x_9175;
assign x_40466 = x_40464 & x_40465;
assign x_40467 = x_40463 & x_40466;
assign x_40468 = x_9176 & x_9177;
assign x_40469 = x_9178 & x_9179;
assign x_40470 = x_40468 & x_40469;
assign x_40471 = x_9180 & x_9181;
assign x_40472 = x_9182 & x_9183;
assign x_40473 = x_40471 & x_40472;
assign x_40474 = x_40470 & x_40473;
assign x_40475 = x_40467 & x_40474;
assign x_40476 = x_9185 & x_9186;
assign x_40477 = x_9184 & x_40476;
assign x_40478 = x_9187 & x_9188;
assign x_40479 = x_9189 & x_9190;
assign x_40480 = x_40478 & x_40479;
assign x_40481 = x_40477 & x_40480;
assign x_40482 = x_9191 & x_9192;
assign x_40483 = x_9193 & x_9194;
assign x_40484 = x_40482 & x_40483;
assign x_40485 = x_9195 & x_9196;
assign x_40486 = x_9197 & x_9198;
assign x_40487 = x_40485 & x_40486;
assign x_40488 = x_40484 & x_40487;
assign x_40489 = x_40481 & x_40488;
assign x_40490 = x_40475 & x_40489;
assign x_40491 = x_9200 & x_9201;
assign x_40492 = x_9199 & x_40491;
assign x_40493 = x_9202 & x_9203;
assign x_40494 = x_9204 & x_9205;
assign x_40495 = x_40493 & x_40494;
assign x_40496 = x_40492 & x_40495;
assign x_40497 = x_9206 & x_9207;
assign x_40498 = x_9208 & x_9209;
assign x_40499 = x_40497 & x_40498;
assign x_40500 = x_9210 & x_9211;
assign x_40501 = x_9212 & x_9213;
assign x_40502 = x_40500 & x_40501;
assign x_40503 = x_40499 & x_40502;
assign x_40504 = x_40496 & x_40503;
assign x_40505 = x_9214 & x_9215;
assign x_40506 = x_9216 & x_9217;
assign x_40507 = x_40505 & x_40506;
assign x_40508 = x_9218 & x_9219;
assign x_40509 = x_9220 & x_9221;
assign x_40510 = x_40508 & x_40509;
assign x_40511 = x_40507 & x_40510;
assign x_40512 = x_9222 & x_9223;
assign x_40513 = x_9224 & x_9225;
assign x_40514 = x_40512 & x_40513;
assign x_40515 = x_9226 & x_9227;
assign x_40516 = x_9228 & x_9229;
assign x_40517 = x_40515 & x_40516;
assign x_40518 = x_40514 & x_40517;
assign x_40519 = x_40511 & x_40518;
assign x_40520 = x_40504 & x_40519;
assign x_40521 = x_40490 & x_40520;
assign x_40522 = x_9231 & x_9232;
assign x_40523 = x_9230 & x_40522;
assign x_40524 = x_9233 & x_9234;
assign x_40525 = x_9235 & x_9236;
assign x_40526 = x_40524 & x_40525;
assign x_40527 = x_40523 & x_40526;
assign x_40528 = x_9237 & x_9238;
assign x_40529 = x_9239 & x_9240;
assign x_40530 = x_40528 & x_40529;
assign x_40531 = x_9241 & x_9242;
assign x_40532 = x_9243 & x_9244;
assign x_40533 = x_40531 & x_40532;
assign x_40534 = x_40530 & x_40533;
assign x_40535 = x_40527 & x_40534;
assign x_40536 = x_9245 & x_9246;
assign x_40537 = x_9247 & x_9248;
assign x_40538 = x_40536 & x_40537;
assign x_40539 = x_9249 & x_9250;
assign x_40540 = x_9251 & x_9252;
assign x_40541 = x_40539 & x_40540;
assign x_40542 = x_40538 & x_40541;
assign x_40543 = x_9253 & x_9254;
assign x_40544 = x_9255 & x_9256;
assign x_40545 = x_40543 & x_40544;
assign x_40546 = x_9257 & x_9258;
assign x_40547 = x_9259 & x_9260;
assign x_40548 = x_40546 & x_40547;
assign x_40549 = x_40545 & x_40548;
assign x_40550 = x_40542 & x_40549;
assign x_40551 = x_40535 & x_40550;
assign x_40552 = x_9262 & x_9263;
assign x_40553 = x_9261 & x_40552;
assign x_40554 = x_9264 & x_9265;
assign x_40555 = x_9266 & x_9267;
assign x_40556 = x_40554 & x_40555;
assign x_40557 = x_40553 & x_40556;
assign x_40558 = x_9268 & x_9269;
assign x_40559 = x_9270 & x_9271;
assign x_40560 = x_40558 & x_40559;
assign x_40561 = x_9272 & x_9273;
assign x_40562 = x_9274 & x_9275;
assign x_40563 = x_40561 & x_40562;
assign x_40564 = x_40560 & x_40563;
assign x_40565 = x_40557 & x_40564;
assign x_40566 = x_9276 & x_9277;
assign x_40567 = x_9278 & x_9279;
assign x_40568 = x_40566 & x_40567;
assign x_40569 = x_9280 & x_9281;
assign x_40570 = x_9282 & x_9283;
assign x_40571 = x_40569 & x_40570;
assign x_40572 = x_40568 & x_40571;
assign x_40573 = x_9284 & x_9285;
assign x_40574 = x_9286 & x_9287;
assign x_40575 = x_40573 & x_40574;
assign x_40576 = x_9288 & x_9289;
assign x_40577 = x_9290 & x_9291;
assign x_40578 = x_40576 & x_40577;
assign x_40579 = x_40575 & x_40578;
assign x_40580 = x_40572 & x_40579;
assign x_40581 = x_40565 & x_40580;
assign x_40582 = x_40551 & x_40581;
assign x_40583 = x_40521 & x_40582;
assign x_40584 = x_40461 & x_40583;
assign x_40585 = x_40340 & x_40584;
assign x_40586 = x_9293 & x_9294;
assign x_40587 = x_9292 & x_40586;
assign x_40588 = x_9295 & x_9296;
assign x_40589 = x_9297 & x_9298;
assign x_40590 = x_40588 & x_40589;
assign x_40591 = x_40587 & x_40590;
assign x_40592 = x_9299 & x_9300;
assign x_40593 = x_9301 & x_9302;
assign x_40594 = x_40592 & x_40593;
assign x_40595 = x_9303 & x_9304;
assign x_40596 = x_9305 & x_9306;
assign x_40597 = x_40595 & x_40596;
assign x_40598 = x_40594 & x_40597;
assign x_40599 = x_40591 & x_40598;
assign x_40600 = x_9308 & x_9309;
assign x_40601 = x_9307 & x_40600;
assign x_40602 = x_9310 & x_9311;
assign x_40603 = x_9312 & x_9313;
assign x_40604 = x_40602 & x_40603;
assign x_40605 = x_40601 & x_40604;
assign x_40606 = x_9314 & x_9315;
assign x_40607 = x_9316 & x_9317;
assign x_40608 = x_40606 & x_40607;
assign x_40609 = x_9318 & x_9319;
assign x_40610 = x_9320 & x_9321;
assign x_40611 = x_40609 & x_40610;
assign x_40612 = x_40608 & x_40611;
assign x_40613 = x_40605 & x_40612;
assign x_40614 = x_40599 & x_40613;
assign x_40615 = x_9323 & x_9324;
assign x_40616 = x_9322 & x_40615;
assign x_40617 = x_9325 & x_9326;
assign x_40618 = x_9327 & x_9328;
assign x_40619 = x_40617 & x_40618;
assign x_40620 = x_40616 & x_40619;
assign x_40621 = x_9329 & x_9330;
assign x_40622 = x_9331 & x_9332;
assign x_40623 = x_40621 & x_40622;
assign x_40624 = x_9333 & x_9334;
assign x_40625 = x_9335 & x_9336;
assign x_40626 = x_40624 & x_40625;
assign x_40627 = x_40623 & x_40626;
assign x_40628 = x_40620 & x_40627;
assign x_40629 = x_9337 & x_9338;
assign x_40630 = x_9339 & x_9340;
assign x_40631 = x_40629 & x_40630;
assign x_40632 = x_9341 & x_9342;
assign x_40633 = x_9343 & x_9344;
assign x_40634 = x_40632 & x_40633;
assign x_40635 = x_40631 & x_40634;
assign x_40636 = x_9345 & x_9346;
assign x_40637 = x_9347 & x_9348;
assign x_40638 = x_40636 & x_40637;
assign x_40639 = x_9349 & x_9350;
assign x_40640 = x_9351 & x_9352;
assign x_40641 = x_40639 & x_40640;
assign x_40642 = x_40638 & x_40641;
assign x_40643 = x_40635 & x_40642;
assign x_40644 = x_40628 & x_40643;
assign x_40645 = x_40614 & x_40644;
assign x_40646 = x_9354 & x_9355;
assign x_40647 = x_9353 & x_40646;
assign x_40648 = x_9356 & x_9357;
assign x_40649 = x_9358 & x_9359;
assign x_40650 = x_40648 & x_40649;
assign x_40651 = x_40647 & x_40650;
assign x_40652 = x_9360 & x_9361;
assign x_40653 = x_9362 & x_9363;
assign x_40654 = x_40652 & x_40653;
assign x_40655 = x_9364 & x_9365;
assign x_40656 = x_9366 & x_9367;
assign x_40657 = x_40655 & x_40656;
assign x_40658 = x_40654 & x_40657;
assign x_40659 = x_40651 & x_40658;
assign x_40660 = x_9369 & x_9370;
assign x_40661 = x_9368 & x_40660;
assign x_40662 = x_9371 & x_9372;
assign x_40663 = x_9373 & x_9374;
assign x_40664 = x_40662 & x_40663;
assign x_40665 = x_40661 & x_40664;
assign x_40666 = x_9375 & x_9376;
assign x_40667 = x_9377 & x_9378;
assign x_40668 = x_40666 & x_40667;
assign x_40669 = x_9379 & x_9380;
assign x_40670 = x_9381 & x_9382;
assign x_40671 = x_40669 & x_40670;
assign x_40672 = x_40668 & x_40671;
assign x_40673 = x_40665 & x_40672;
assign x_40674 = x_40659 & x_40673;
assign x_40675 = x_9384 & x_9385;
assign x_40676 = x_9383 & x_40675;
assign x_40677 = x_9386 & x_9387;
assign x_40678 = x_9388 & x_9389;
assign x_40679 = x_40677 & x_40678;
assign x_40680 = x_40676 & x_40679;
assign x_40681 = x_9390 & x_9391;
assign x_40682 = x_9392 & x_9393;
assign x_40683 = x_40681 & x_40682;
assign x_40684 = x_9394 & x_9395;
assign x_40685 = x_9396 & x_9397;
assign x_40686 = x_40684 & x_40685;
assign x_40687 = x_40683 & x_40686;
assign x_40688 = x_40680 & x_40687;
assign x_40689 = x_9398 & x_9399;
assign x_40690 = x_9400 & x_9401;
assign x_40691 = x_40689 & x_40690;
assign x_40692 = x_9402 & x_9403;
assign x_40693 = x_9404 & x_9405;
assign x_40694 = x_40692 & x_40693;
assign x_40695 = x_40691 & x_40694;
assign x_40696 = x_9406 & x_9407;
assign x_40697 = x_9408 & x_9409;
assign x_40698 = x_40696 & x_40697;
assign x_40699 = x_9410 & x_9411;
assign x_40700 = x_9412 & x_9413;
assign x_40701 = x_40699 & x_40700;
assign x_40702 = x_40698 & x_40701;
assign x_40703 = x_40695 & x_40702;
assign x_40704 = x_40688 & x_40703;
assign x_40705 = x_40674 & x_40704;
assign x_40706 = x_40645 & x_40705;
assign x_40707 = x_9415 & x_9416;
assign x_40708 = x_9414 & x_40707;
assign x_40709 = x_9417 & x_9418;
assign x_40710 = x_9419 & x_9420;
assign x_40711 = x_40709 & x_40710;
assign x_40712 = x_40708 & x_40711;
assign x_40713 = x_9421 & x_9422;
assign x_40714 = x_9423 & x_9424;
assign x_40715 = x_40713 & x_40714;
assign x_40716 = x_9425 & x_9426;
assign x_40717 = x_9427 & x_9428;
assign x_40718 = x_40716 & x_40717;
assign x_40719 = x_40715 & x_40718;
assign x_40720 = x_40712 & x_40719;
assign x_40721 = x_9430 & x_9431;
assign x_40722 = x_9429 & x_40721;
assign x_40723 = x_9432 & x_9433;
assign x_40724 = x_9434 & x_9435;
assign x_40725 = x_40723 & x_40724;
assign x_40726 = x_40722 & x_40725;
assign x_40727 = x_9436 & x_9437;
assign x_40728 = x_9438 & x_9439;
assign x_40729 = x_40727 & x_40728;
assign x_40730 = x_9440 & x_9441;
assign x_40731 = x_9442 & x_9443;
assign x_40732 = x_40730 & x_40731;
assign x_40733 = x_40729 & x_40732;
assign x_40734 = x_40726 & x_40733;
assign x_40735 = x_40720 & x_40734;
assign x_40736 = x_9445 & x_9446;
assign x_40737 = x_9444 & x_40736;
assign x_40738 = x_9447 & x_9448;
assign x_40739 = x_9449 & x_9450;
assign x_40740 = x_40738 & x_40739;
assign x_40741 = x_40737 & x_40740;
assign x_40742 = x_9451 & x_9452;
assign x_40743 = x_9453 & x_9454;
assign x_40744 = x_40742 & x_40743;
assign x_40745 = x_9455 & x_9456;
assign x_40746 = x_9457 & x_9458;
assign x_40747 = x_40745 & x_40746;
assign x_40748 = x_40744 & x_40747;
assign x_40749 = x_40741 & x_40748;
assign x_40750 = x_9459 & x_9460;
assign x_40751 = x_9461 & x_9462;
assign x_40752 = x_40750 & x_40751;
assign x_40753 = x_9463 & x_9464;
assign x_40754 = x_9465 & x_9466;
assign x_40755 = x_40753 & x_40754;
assign x_40756 = x_40752 & x_40755;
assign x_40757 = x_9467 & x_9468;
assign x_40758 = x_9469 & x_9470;
assign x_40759 = x_40757 & x_40758;
assign x_40760 = x_9471 & x_9472;
assign x_40761 = x_9473 & x_9474;
assign x_40762 = x_40760 & x_40761;
assign x_40763 = x_40759 & x_40762;
assign x_40764 = x_40756 & x_40763;
assign x_40765 = x_40749 & x_40764;
assign x_40766 = x_40735 & x_40765;
assign x_40767 = x_9476 & x_9477;
assign x_40768 = x_9475 & x_40767;
assign x_40769 = x_9478 & x_9479;
assign x_40770 = x_9480 & x_9481;
assign x_40771 = x_40769 & x_40770;
assign x_40772 = x_40768 & x_40771;
assign x_40773 = x_9482 & x_9483;
assign x_40774 = x_9484 & x_9485;
assign x_40775 = x_40773 & x_40774;
assign x_40776 = x_9486 & x_9487;
assign x_40777 = x_9488 & x_9489;
assign x_40778 = x_40776 & x_40777;
assign x_40779 = x_40775 & x_40778;
assign x_40780 = x_40772 & x_40779;
assign x_40781 = x_9491 & x_9492;
assign x_40782 = x_9490 & x_40781;
assign x_40783 = x_9493 & x_9494;
assign x_40784 = x_9495 & x_9496;
assign x_40785 = x_40783 & x_40784;
assign x_40786 = x_40782 & x_40785;
assign x_40787 = x_9497 & x_9498;
assign x_40788 = x_9499 & x_9500;
assign x_40789 = x_40787 & x_40788;
assign x_40790 = x_9501 & x_9502;
assign x_40791 = x_9503 & x_9504;
assign x_40792 = x_40790 & x_40791;
assign x_40793 = x_40789 & x_40792;
assign x_40794 = x_40786 & x_40793;
assign x_40795 = x_40780 & x_40794;
assign x_40796 = x_9506 & x_9507;
assign x_40797 = x_9505 & x_40796;
assign x_40798 = x_9508 & x_9509;
assign x_40799 = x_9510 & x_9511;
assign x_40800 = x_40798 & x_40799;
assign x_40801 = x_40797 & x_40800;
assign x_40802 = x_9512 & x_9513;
assign x_40803 = x_9514 & x_9515;
assign x_40804 = x_40802 & x_40803;
assign x_40805 = x_9516 & x_9517;
assign x_40806 = x_9518 & x_9519;
assign x_40807 = x_40805 & x_40806;
assign x_40808 = x_40804 & x_40807;
assign x_40809 = x_40801 & x_40808;
assign x_40810 = x_9520 & x_9521;
assign x_40811 = x_9522 & x_9523;
assign x_40812 = x_40810 & x_40811;
assign x_40813 = x_9524 & x_9525;
assign x_40814 = x_9526 & x_9527;
assign x_40815 = x_40813 & x_40814;
assign x_40816 = x_40812 & x_40815;
assign x_40817 = x_9528 & x_9529;
assign x_40818 = x_9530 & x_9531;
assign x_40819 = x_40817 & x_40818;
assign x_40820 = x_9532 & x_9533;
assign x_40821 = x_9534 & x_9535;
assign x_40822 = x_40820 & x_40821;
assign x_40823 = x_40819 & x_40822;
assign x_40824 = x_40816 & x_40823;
assign x_40825 = x_40809 & x_40824;
assign x_40826 = x_40795 & x_40825;
assign x_40827 = x_40766 & x_40826;
assign x_40828 = x_40706 & x_40827;
assign x_40829 = x_9537 & x_9538;
assign x_40830 = x_9536 & x_40829;
assign x_40831 = x_9539 & x_9540;
assign x_40832 = x_9541 & x_9542;
assign x_40833 = x_40831 & x_40832;
assign x_40834 = x_40830 & x_40833;
assign x_40835 = x_9543 & x_9544;
assign x_40836 = x_9545 & x_9546;
assign x_40837 = x_40835 & x_40836;
assign x_40838 = x_9547 & x_9548;
assign x_40839 = x_9549 & x_9550;
assign x_40840 = x_40838 & x_40839;
assign x_40841 = x_40837 & x_40840;
assign x_40842 = x_40834 & x_40841;
assign x_40843 = x_9552 & x_9553;
assign x_40844 = x_9551 & x_40843;
assign x_40845 = x_9554 & x_9555;
assign x_40846 = x_9556 & x_9557;
assign x_40847 = x_40845 & x_40846;
assign x_40848 = x_40844 & x_40847;
assign x_40849 = x_9558 & x_9559;
assign x_40850 = x_9560 & x_9561;
assign x_40851 = x_40849 & x_40850;
assign x_40852 = x_9562 & x_9563;
assign x_40853 = x_9564 & x_9565;
assign x_40854 = x_40852 & x_40853;
assign x_40855 = x_40851 & x_40854;
assign x_40856 = x_40848 & x_40855;
assign x_40857 = x_40842 & x_40856;
assign x_40858 = x_9567 & x_9568;
assign x_40859 = x_9566 & x_40858;
assign x_40860 = x_9569 & x_9570;
assign x_40861 = x_9571 & x_9572;
assign x_40862 = x_40860 & x_40861;
assign x_40863 = x_40859 & x_40862;
assign x_40864 = x_9573 & x_9574;
assign x_40865 = x_9575 & x_9576;
assign x_40866 = x_40864 & x_40865;
assign x_40867 = x_9577 & x_9578;
assign x_40868 = x_9579 & x_9580;
assign x_40869 = x_40867 & x_40868;
assign x_40870 = x_40866 & x_40869;
assign x_40871 = x_40863 & x_40870;
assign x_40872 = x_9581 & x_9582;
assign x_40873 = x_9583 & x_9584;
assign x_40874 = x_40872 & x_40873;
assign x_40875 = x_9585 & x_9586;
assign x_40876 = x_9587 & x_9588;
assign x_40877 = x_40875 & x_40876;
assign x_40878 = x_40874 & x_40877;
assign x_40879 = x_9589 & x_9590;
assign x_40880 = x_9591 & x_9592;
assign x_40881 = x_40879 & x_40880;
assign x_40882 = x_9593 & x_9594;
assign x_40883 = x_9595 & x_9596;
assign x_40884 = x_40882 & x_40883;
assign x_40885 = x_40881 & x_40884;
assign x_40886 = x_40878 & x_40885;
assign x_40887 = x_40871 & x_40886;
assign x_40888 = x_40857 & x_40887;
assign x_40889 = x_9598 & x_9599;
assign x_40890 = x_9597 & x_40889;
assign x_40891 = x_9600 & x_9601;
assign x_40892 = x_9602 & x_9603;
assign x_40893 = x_40891 & x_40892;
assign x_40894 = x_40890 & x_40893;
assign x_40895 = x_9604 & x_9605;
assign x_40896 = x_9606 & x_9607;
assign x_40897 = x_40895 & x_40896;
assign x_40898 = x_9608 & x_9609;
assign x_40899 = x_9610 & x_9611;
assign x_40900 = x_40898 & x_40899;
assign x_40901 = x_40897 & x_40900;
assign x_40902 = x_40894 & x_40901;
assign x_40903 = x_9613 & x_9614;
assign x_40904 = x_9612 & x_40903;
assign x_40905 = x_9615 & x_9616;
assign x_40906 = x_9617 & x_9618;
assign x_40907 = x_40905 & x_40906;
assign x_40908 = x_40904 & x_40907;
assign x_40909 = x_9619 & x_9620;
assign x_40910 = x_9621 & x_9622;
assign x_40911 = x_40909 & x_40910;
assign x_40912 = x_9623 & x_9624;
assign x_40913 = x_9625 & x_9626;
assign x_40914 = x_40912 & x_40913;
assign x_40915 = x_40911 & x_40914;
assign x_40916 = x_40908 & x_40915;
assign x_40917 = x_40902 & x_40916;
assign x_40918 = x_9628 & x_9629;
assign x_40919 = x_9627 & x_40918;
assign x_40920 = x_9630 & x_9631;
assign x_40921 = x_9632 & x_9633;
assign x_40922 = x_40920 & x_40921;
assign x_40923 = x_40919 & x_40922;
assign x_40924 = x_9634 & x_9635;
assign x_40925 = x_9636 & x_9637;
assign x_40926 = x_40924 & x_40925;
assign x_40927 = x_9638 & x_9639;
assign x_40928 = x_9640 & x_9641;
assign x_40929 = x_40927 & x_40928;
assign x_40930 = x_40926 & x_40929;
assign x_40931 = x_40923 & x_40930;
assign x_40932 = x_9642 & x_9643;
assign x_40933 = x_9644 & x_9645;
assign x_40934 = x_40932 & x_40933;
assign x_40935 = x_9646 & x_9647;
assign x_40936 = x_9648 & x_9649;
assign x_40937 = x_40935 & x_40936;
assign x_40938 = x_40934 & x_40937;
assign x_40939 = x_9650 & x_9651;
assign x_40940 = x_9652 & x_9653;
assign x_40941 = x_40939 & x_40940;
assign x_40942 = x_9654 & x_9655;
assign x_40943 = x_9656 & x_9657;
assign x_40944 = x_40942 & x_40943;
assign x_40945 = x_40941 & x_40944;
assign x_40946 = x_40938 & x_40945;
assign x_40947 = x_40931 & x_40946;
assign x_40948 = x_40917 & x_40947;
assign x_40949 = x_40888 & x_40948;
assign x_40950 = x_9659 & x_9660;
assign x_40951 = x_9658 & x_40950;
assign x_40952 = x_9661 & x_9662;
assign x_40953 = x_9663 & x_9664;
assign x_40954 = x_40952 & x_40953;
assign x_40955 = x_40951 & x_40954;
assign x_40956 = x_9665 & x_9666;
assign x_40957 = x_9667 & x_9668;
assign x_40958 = x_40956 & x_40957;
assign x_40959 = x_9669 & x_9670;
assign x_40960 = x_9671 & x_9672;
assign x_40961 = x_40959 & x_40960;
assign x_40962 = x_40958 & x_40961;
assign x_40963 = x_40955 & x_40962;
assign x_40964 = x_9674 & x_9675;
assign x_40965 = x_9673 & x_40964;
assign x_40966 = x_9676 & x_9677;
assign x_40967 = x_9678 & x_9679;
assign x_40968 = x_40966 & x_40967;
assign x_40969 = x_40965 & x_40968;
assign x_40970 = x_9680 & x_9681;
assign x_40971 = x_9682 & x_9683;
assign x_40972 = x_40970 & x_40971;
assign x_40973 = x_9684 & x_9685;
assign x_40974 = x_9686 & x_9687;
assign x_40975 = x_40973 & x_40974;
assign x_40976 = x_40972 & x_40975;
assign x_40977 = x_40969 & x_40976;
assign x_40978 = x_40963 & x_40977;
assign x_40979 = x_9689 & x_9690;
assign x_40980 = x_9688 & x_40979;
assign x_40981 = x_9691 & x_9692;
assign x_40982 = x_9693 & x_9694;
assign x_40983 = x_40981 & x_40982;
assign x_40984 = x_40980 & x_40983;
assign x_40985 = x_9695 & x_9696;
assign x_40986 = x_9697 & x_9698;
assign x_40987 = x_40985 & x_40986;
assign x_40988 = x_9699 & x_9700;
assign x_40989 = x_9701 & x_9702;
assign x_40990 = x_40988 & x_40989;
assign x_40991 = x_40987 & x_40990;
assign x_40992 = x_40984 & x_40991;
assign x_40993 = x_9703 & x_9704;
assign x_40994 = x_9705 & x_9706;
assign x_40995 = x_40993 & x_40994;
assign x_40996 = x_9707 & x_9708;
assign x_40997 = x_9709 & x_9710;
assign x_40998 = x_40996 & x_40997;
assign x_40999 = x_40995 & x_40998;
assign x_41000 = x_9711 & x_9712;
assign x_41001 = x_9713 & x_9714;
assign x_41002 = x_41000 & x_41001;
assign x_41003 = x_9715 & x_9716;
assign x_41004 = x_9717 & x_9718;
assign x_41005 = x_41003 & x_41004;
assign x_41006 = x_41002 & x_41005;
assign x_41007 = x_40999 & x_41006;
assign x_41008 = x_40992 & x_41007;
assign x_41009 = x_40978 & x_41008;
assign x_41010 = x_9720 & x_9721;
assign x_41011 = x_9719 & x_41010;
assign x_41012 = x_9722 & x_9723;
assign x_41013 = x_9724 & x_9725;
assign x_41014 = x_41012 & x_41013;
assign x_41015 = x_41011 & x_41014;
assign x_41016 = x_9726 & x_9727;
assign x_41017 = x_9728 & x_9729;
assign x_41018 = x_41016 & x_41017;
assign x_41019 = x_9730 & x_9731;
assign x_41020 = x_9732 & x_9733;
assign x_41021 = x_41019 & x_41020;
assign x_41022 = x_41018 & x_41021;
assign x_41023 = x_41015 & x_41022;
assign x_41024 = x_9734 & x_9735;
assign x_41025 = x_9736 & x_9737;
assign x_41026 = x_41024 & x_41025;
assign x_41027 = x_9738 & x_9739;
assign x_41028 = x_9740 & x_9741;
assign x_41029 = x_41027 & x_41028;
assign x_41030 = x_41026 & x_41029;
assign x_41031 = x_9742 & x_9743;
assign x_41032 = x_9744 & x_9745;
assign x_41033 = x_41031 & x_41032;
assign x_41034 = x_9746 & x_9747;
assign x_41035 = x_9748 & x_9749;
assign x_41036 = x_41034 & x_41035;
assign x_41037 = x_41033 & x_41036;
assign x_41038 = x_41030 & x_41037;
assign x_41039 = x_41023 & x_41038;
assign x_41040 = x_9751 & x_9752;
assign x_41041 = x_9750 & x_41040;
assign x_41042 = x_9753 & x_9754;
assign x_41043 = x_9755 & x_9756;
assign x_41044 = x_41042 & x_41043;
assign x_41045 = x_41041 & x_41044;
assign x_41046 = x_9757 & x_9758;
assign x_41047 = x_9759 & x_9760;
assign x_41048 = x_41046 & x_41047;
assign x_41049 = x_9761 & x_9762;
assign x_41050 = x_9763 & x_9764;
assign x_41051 = x_41049 & x_41050;
assign x_41052 = x_41048 & x_41051;
assign x_41053 = x_41045 & x_41052;
assign x_41054 = x_9765 & x_9766;
assign x_41055 = x_9767 & x_9768;
assign x_41056 = x_41054 & x_41055;
assign x_41057 = x_9769 & x_9770;
assign x_41058 = x_9771 & x_9772;
assign x_41059 = x_41057 & x_41058;
assign x_41060 = x_41056 & x_41059;
assign x_41061 = x_9773 & x_9774;
assign x_41062 = x_9775 & x_9776;
assign x_41063 = x_41061 & x_41062;
assign x_41064 = x_9777 & x_9778;
assign x_41065 = x_9779 & x_9780;
assign x_41066 = x_41064 & x_41065;
assign x_41067 = x_41063 & x_41066;
assign x_41068 = x_41060 & x_41067;
assign x_41069 = x_41053 & x_41068;
assign x_41070 = x_41039 & x_41069;
assign x_41071 = x_41009 & x_41070;
assign x_41072 = x_40949 & x_41071;
assign x_41073 = x_40828 & x_41072;
assign x_41074 = x_40585 & x_41073;
assign x_41075 = x_40097 & x_41074;
assign x_41076 = x_9782 & x_9783;
assign x_41077 = x_9781 & x_41076;
assign x_41078 = x_9784 & x_9785;
assign x_41079 = x_9786 & x_9787;
assign x_41080 = x_41078 & x_41079;
assign x_41081 = x_41077 & x_41080;
assign x_41082 = x_9788 & x_9789;
assign x_41083 = x_9790 & x_9791;
assign x_41084 = x_41082 & x_41083;
assign x_41085 = x_9792 & x_9793;
assign x_41086 = x_9794 & x_9795;
assign x_41087 = x_41085 & x_41086;
assign x_41088 = x_41084 & x_41087;
assign x_41089 = x_41081 & x_41088;
assign x_41090 = x_9797 & x_9798;
assign x_41091 = x_9796 & x_41090;
assign x_41092 = x_9799 & x_9800;
assign x_41093 = x_9801 & x_9802;
assign x_41094 = x_41092 & x_41093;
assign x_41095 = x_41091 & x_41094;
assign x_41096 = x_9803 & x_9804;
assign x_41097 = x_9805 & x_9806;
assign x_41098 = x_41096 & x_41097;
assign x_41099 = x_9807 & x_9808;
assign x_41100 = x_9809 & x_9810;
assign x_41101 = x_41099 & x_41100;
assign x_41102 = x_41098 & x_41101;
assign x_41103 = x_41095 & x_41102;
assign x_41104 = x_41089 & x_41103;
assign x_41105 = x_9812 & x_9813;
assign x_41106 = x_9811 & x_41105;
assign x_41107 = x_9814 & x_9815;
assign x_41108 = x_9816 & x_9817;
assign x_41109 = x_41107 & x_41108;
assign x_41110 = x_41106 & x_41109;
assign x_41111 = x_9818 & x_9819;
assign x_41112 = x_9820 & x_9821;
assign x_41113 = x_41111 & x_41112;
assign x_41114 = x_9822 & x_9823;
assign x_41115 = x_9824 & x_9825;
assign x_41116 = x_41114 & x_41115;
assign x_41117 = x_41113 & x_41116;
assign x_41118 = x_41110 & x_41117;
assign x_41119 = x_9826 & x_9827;
assign x_41120 = x_9828 & x_9829;
assign x_41121 = x_41119 & x_41120;
assign x_41122 = x_9830 & x_9831;
assign x_41123 = x_9832 & x_9833;
assign x_41124 = x_41122 & x_41123;
assign x_41125 = x_41121 & x_41124;
assign x_41126 = x_9834 & x_9835;
assign x_41127 = x_9836 & x_9837;
assign x_41128 = x_41126 & x_41127;
assign x_41129 = x_9838 & x_9839;
assign x_41130 = x_9840 & x_9841;
assign x_41131 = x_41129 & x_41130;
assign x_41132 = x_41128 & x_41131;
assign x_41133 = x_41125 & x_41132;
assign x_41134 = x_41118 & x_41133;
assign x_41135 = x_41104 & x_41134;
assign x_41136 = x_9843 & x_9844;
assign x_41137 = x_9842 & x_41136;
assign x_41138 = x_9845 & x_9846;
assign x_41139 = x_9847 & x_9848;
assign x_41140 = x_41138 & x_41139;
assign x_41141 = x_41137 & x_41140;
assign x_41142 = x_9849 & x_9850;
assign x_41143 = x_9851 & x_9852;
assign x_41144 = x_41142 & x_41143;
assign x_41145 = x_9853 & x_9854;
assign x_41146 = x_9855 & x_9856;
assign x_41147 = x_41145 & x_41146;
assign x_41148 = x_41144 & x_41147;
assign x_41149 = x_41141 & x_41148;
assign x_41150 = x_9858 & x_9859;
assign x_41151 = x_9857 & x_41150;
assign x_41152 = x_9860 & x_9861;
assign x_41153 = x_9862 & x_9863;
assign x_41154 = x_41152 & x_41153;
assign x_41155 = x_41151 & x_41154;
assign x_41156 = x_9864 & x_9865;
assign x_41157 = x_9866 & x_9867;
assign x_41158 = x_41156 & x_41157;
assign x_41159 = x_9868 & x_9869;
assign x_41160 = x_9870 & x_9871;
assign x_41161 = x_41159 & x_41160;
assign x_41162 = x_41158 & x_41161;
assign x_41163 = x_41155 & x_41162;
assign x_41164 = x_41149 & x_41163;
assign x_41165 = x_9873 & x_9874;
assign x_41166 = x_9872 & x_41165;
assign x_41167 = x_9875 & x_9876;
assign x_41168 = x_9877 & x_9878;
assign x_41169 = x_41167 & x_41168;
assign x_41170 = x_41166 & x_41169;
assign x_41171 = x_9879 & x_9880;
assign x_41172 = x_9881 & x_9882;
assign x_41173 = x_41171 & x_41172;
assign x_41174 = x_9883 & x_9884;
assign x_41175 = x_9885 & x_9886;
assign x_41176 = x_41174 & x_41175;
assign x_41177 = x_41173 & x_41176;
assign x_41178 = x_41170 & x_41177;
assign x_41179 = x_9887 & x_9888;
assign x_41180 = x_9889 & x_9890;
assign x_41181 = x_41179 & x_41180;
assign x_41182 = x_9891 & x_9892;
assign x_41183 = x_9893 & x_9894;
assign x_41184 = x_41182 & x_41183;
assign x_41185 = x_41181 & x_41184;
assign x_41186 = x_9895 & x_9896;
assign x_41187 = x_9897 & x_9898;
assign x_41188 = x_41186 & x_41187;
assign x_41189 = x_9899 & x_9900;
assign x_41190 = x_9901 & x_9902;
assign x_41191 = x_41189 & x_41190;
assign x_41192 = x_41188 & x_41191;
assign x_41193 = x_41185 & x_41192;
assign x_41194 = x_41178 & x_41193;
assign x_41195 = x_41164 & x_41194;
assign x_41196 = x_41135 & x_41195;
assign x_41197 = x_9904 & x_9905;
assign x_41198 = x_9903 & x_41197;
assign x_41199 = x_9906 & x_9907;
assign x_41200 = x_9908 & x_9909;
assign x_41201 = x_41199 & x_41200;
assign x_41202 = x_41198 & x_41201;
assign x_41203 = x_9910 & x_9911;
assign x_41204 = x_9912 & x_9913;
assign x_41205 = x_41203 & x_41204;
assign x_41206 = x_9914 & x_9915;
assign x_41207 = x_9916 & x_9917;
assign x_41208 = x_41206 & x_41207;
assign x_41209 = x_41205 & x_41208;
assign x_41210 = x_41202 & x_41209;
assign x_41211 = x_9919 & x_9920;
assign x_41212 = x_9918 & x_41211;
assign x_41213 = x_9921 & x_9922;
assign x_41214 = x_9923 & x_9924;
assign x_41215 = x_41213 & x_41214;
assign x_41216 = x_41212 & x_41215;
assign x_41217 = x_9925 & x_9926;
assign x_41218 = x_9927 & x_9928;
assign x_41219 = x_41217 & x_41218;
assign x_41220 = x_9929 & x_9930;
assign x_41221 = x_9931 & x_9932;
assign x_41222 = x_41220 & x_41221;
assign x_41223 = x_41219 & x_41222;
assign x_41224 = x_41216 & x_41223;
assign x_41225 = x_41210 & x_41224;
assign x_41226 = x_9934 & x_9935;
assign x_41227 = x_9933 & x_41226;
assign x_41228 = x_9936 & x_9937;
assign x_41229 = x_9938 & x_9939;
assign x_41230 = x_41228 & x_41229;
assign x_41231 = x_41227 & x_41230;
assign x_41232 = x_9940 & x_9941;
assign x_41233 = x_9942 & x_9943;
assign x_41234 = x_41232 & x_41233;
assign x_41235 = x_9944 & x_9945;
assign x_41236 = x_9946 & x_9947;
assign x_41237 = x_41235 & x_41236;
assign x_41238 = x_41234 & x_41237;
assign x_41239 = x_41231 & x_41238;
assign x_41240 = x_9948 & x_9949;
assign x_41241 = x_9950 & x_9951;
assign x_41242 = x_41240 & x_41241;
assign x_41243 = x_9952 & x_9953;
assign x_41244 = x_9954 & x_9955;
assign x_41245 = x_41243 & x_41244;
assign x_41246 = x_41242 & x_41245;
assign x_41247 = x_9956 & x_9957;
assign x_41248 = x_9958 & x_9959;
assign x_41249 = x_41247 & x_41248;
assign x_41250 = x_9960 & x_9961;
assign x_41251 = x_9962 & x_9963;
assign x_41252 = x_41250 & x_41251;
assign x_41253 = x_41249 & x_41252;
assign x_41254 = x_41246 & x_41253;
assign x_41255 = x_41239 & x_41254;
assign x_41256 = x_41225 & x_41255;
assign x_41257 = x_9965 & x_9966;
assign x_41258 = x_9964 & x_41257;
assign x_41259 = x_9967 & x_9968;
assign x_41260 = x_9969 & x_9970;
assign x_41261 = x_41259 & x_41260;
assign x_41262 = x_41258 & x_41261;
assign x_41263 = x_9971 & x_9972;
assign x_41264 = x_9973 & x_9974;
assign x_41265 = x_41263 & x_41264;
assign x_41266 = x_9975 & x_9976;
assign x_41267 = x_9977 & x_9978;
assign x_41268 = x_41266 & x_41267;
assign x_41269 = x_41265 & x_41268;
assign x_41270 = x_41262 & x_41269;
assign x_41271 = x_9980 & x_9981;
assign x_41272 = x_9979 & x_41271;
assign x_41273 = x_9982 & x_9983;
assign x_41274 = x_9984 & x_9985;
assign x_41275 = x_41273 & x_41274;
assign x_41276 = x_41272 & x_41275;
assign x_41277 = x_9986 & x_9987;
assign x_41278 = x_9988 & x_9989;
assign x_41279 = x_41277 & x_41278;
assign x_41280 = x_9990 & x_9991;
assign x_41281 = x_9992 & x_9993;
assign x_41282 = x_41280 & x_41281;
assign x_41283 = x_41279 & x_41282;
assign x_41284 = x_41276 & x_41283;
assign x_41285 = x_41270 & x_41284;
assign x_41286 = x_9995 & x_9996;
assign x_41287 = x_9994 & x_41286;
assign x_41288 = x_9997 & x_9998;
assign x_41289 = x_9999 & x_10000;
assign x_41290 = x_41288 & x_41289;
assign x_41291 = x_41287 & x_41290;
assign x_41292 = x_10001 & x_10002;
assign x_41293 = x_10003 & x_10004;
assign x_41294 = x_41292 & x_41293;
assign x_41295 = x_10005 & x_10006;
assign x_41296 = x_10007 & x_10008;
assign x_41297 = x_41295 & x_41296;
assign x_41298 = x_41294 & x_41297;
assign x_41299 = x_41291 & x_41298;
assign x_41300 = x_10009 & x_10010;
assign x_41301 = x_10011 & x_10012;
assign x_41302 = x_41300 & x_41301;
assign x_41303 = x_10013 & x_10014;
assign x_41304 = x_10015 & x_10016;
assign x_41305 = x_41303 & x_41304;
assign x_41306 = x_41302 & x_41305;
assign x_41307 = x_10017 & x_10018;
assign x_41308 = x_10019 & x_10020;
assign x_41309 = x_41307 & x_41308;
assign x_41310 = x_10021 & x_10022;
assign x_41311 = x_10023 & x_10024;
assign x_41312 = x_41310 & x_41311;
assign x_41313 = x_41309 & x_41312;
assign x_41314 = x_41306 & x_41313;
assign x_41315 = x_41299 & x_41314;
assign x_41316 = x_41285 & x_41315;
assign x_41317 = x_41256 & x_41316;
assign x_41318 = x_41196 & x_41317;
assign x_41319 = x_10026 & x_10027;
assign x_41320 = x_10025 & x_41319;
assign x_41321 = x_10028 & x_10029;
assign x_41322 = x_10030 & x_10031;
assign x_41323 = x_41321 & x_41322;
assign x_41324 = x_41320 & x_41323;
assign x_41325 = x_10032 & x_10033;
assign x_41326 = x_10034 & x_10035;
assign x_41327 = x_41325 & x_41326;
assign x_41328 = x_10036 & x_10037;
assign x_41329 = x_10038 & x_10039;
assign x_41330 = x_41328 & x_41329;
assign x_41331 = x_41327 & x_41330;
assign x_41332 = x_41324 & x_41331;
assign x_41333 = x_10041 & x_10042;
assign x_41334 = x_10040 & x_41333;
assign x_41335 = x_10043 & x_10044;
assign x_41336 = x_10045 & x_10046;
assign x_41337 = x_41335 & x_41336;
assign x_41338 = x_41334 & x_41337;
assign x_41339 = x_10047 & x_10048;
assign x_41340 = x_10049 & x_10050;
assign x_41341 = x_41339 & x_41340;
assign x_41342 = x_10051 & x_10052;
assign x_41343 = x_10053 & x_10054;
assign x_41344 = x_41342 & x_41343;
assign x_41345 = x_41341 & x_41344;
assign x_41346 = x_41338 & x_41345;
assign x_41347 = x_41332 & x_41346;
assign x_41348 = x_10056 & x_10057;
assign x_41349 = x_10055 & x_41348;
assign x_41350 = x_10058 & x_10059;
assign x_41351 = x_10060 & x_10061;
assign x_41352 = x_41350 & x_41351;
assign x_41353 = x_41349 & x_41352;
assign x_41354 = x_10062 & x_10063;
assign x_41355 = x_10064 & x_10065;
assign x_41356 = x_41354 & x_41355;
assign x_41357 = x_10066 & x_10067;
assign x_41358 = x_10068 & x_10069;
assign x_41359 = x_41357 & x_41358;
assign x_41360 = x_41356 & x_41359;
assign x_41361 = x_41353 & x_41360;
assign x_41362 = x_10070 & x_10071;
assign x_41363 = x_10072 & x_10073;
assign x_41364 = x_41362 & x_41363;
assign x_41365 = x_10074 & x_10075;
assign x_41366 = x_10076 & x_10077;
assign x_41367 = x_41365 & x_41366;
assign x_41368 = x_41364 & x_41367;
assign x_41369 = x_10078 & x_10079;
assign x_41370 = x_10080 & x_10081;
assign x_41371 = x_41369 & x_41370;
assign x_41372 = x_10082 & x_10083;
assign x_41373 = x_10084 & x_10085;
assign x_41374 = x_41372 & x_41373;
assign x_41375 = x_41371 & x_41374;
assign x_41376 = x_41368 & x_41375;
assign x_41377 = x_41361 & x_41376;
assign x_41378 = x_41347 & x_41377;
assign x_41379 = x_10087 & x_10088;
assign x_41380 = x_10086 & x_41379;
assign x_41381 = x_10089 & x_10090;
assign x_41382 = x_10091 & x_10092;
assign x_41383 = x_41381 & x_41382;
assign x_41384 = x_41380 & x_41383;
assign x_41385 = x_10093 & x_10094;
assign x_41386 = x_10095 & x_10096;
assign x_41387 = x_41385 & x_41386;
assign x_41388 = x_10097 & x_10098;
assign x_41389 = x_10099 & x_10100;
assign x_41390 = x_41388 & x_41389;
assign x_41391 = x_41387 & x_41390;
assign x_41392 = x_41384 & x_41391;
assign x_41393 = x_10102 & x_10103;
assign x_41394 = x_10101 & x_41393;
assign x_41395 = x_10104 & x_10105;
assign x_41396 = x_10106 & x_10107;
assign x_41397 = x_41395 & x_41396;
assign x_41398 = x_41394 & x_41397;
assign x_41399 = x_10108 & x_10109;
assign x_41400 = x_10110 & x_10111;
assign x_41401 = x_41399 & x_41400;
assign x_41402 = x_10112 & x_10113;
assign x_41403 = x_10114 & x_10115;
assign x_41404 = x_41402 & x_41403;
assign x_41405 = x_41401 & x_41404;
assign x_41406 = x_41398 & x_41405;
assign x_41407 = x_41392 & x_41406;
assign x_41408 = x_10117 & x_10118;
assign x_41409 = x_10116 & x_41408;
assign x_41410 = x_10119 & x_10120;
assign x_41411 = x_10121 & x_10122;
assign x_41412 = x_41410 & x_41411;
assign x_41413 = x_41409 & x_41412;
assign x_41414 = x_10123 & x_10124;
assign x_41415 = x_10125 & x_10126;
assign x_41416 = x_41414 & x_41415;
assign x_41417 = x_10127 & x_10128;
assign x_41418 = x_10129 & x_10130;
assign x_41419 = x_41417 & x_41418;
assign x_41420 = x_41416 & x_41419;
assign x_41421 = x_41413 & x_41420;
assign x_41422 = x_10131 & x_10132;
assign x_41423 = x_10133 & x_10134;
assign x_41424 = x_41422 & x_41423;
assign x_41425 = x_10135 & x_10136;
assign x_41426 = x_10137 & x_10138;
assign x_41427 = x_41425 & x_41426;
assign x_41428 = x_41424 & x_41427;
assign x_41429 = x_10139 & x_10140;
assign x_41430 = x_10141 & x_10142;
assign x_41431 = x_41429 & x_41430;
assign x_41432 = x_10143 & x_10144;
assign x_41433 = x_10145 & x_10146;
assign x_41434 = x_41432 & x_41433;
assign x_41435 = x_41431 & x_41434;
assign x_41436 = x_41428 & x_41435;
assign x_41437 = x_41421 & x_41436;
assign x_41438 = x_41407 & x_41437;
assign x_41439 = x_41378 & x_41438;
assign x_41440 = x_10148 & x_10149;
assign x_41441 = x_10147 & x_41440;
assign x_41442 = x_10150 & x_10151;
assign x_41443 = x_10152 & x_10153;
assign x_41444 = x_41442 & x_41443;
assign x_41445 = x_41441 & x_41444;
assign x_41446 = x_10154 & x_10155;
assign x_41447 = x_10156 & x_10157;
assign x_41448 = x_41446 & x_41447;
assign x_41449 = x_10158 & x_10159;
assign x_41450 = x_10160 & x_10161;
assign x_41451 = x_41449 & x_41450;
assign x_41452 = x_41448 & x_41451;
assign x_41453 = x_41445 & x_41452;
assign x_41454 = x_10163 & x_10164;
assign x_41455 = x_10162 & x_41454;
assign x_41456 = x_10165 & x_10166;
assign x_41457 = x_10167 & x_10168;
assign x_41458 = x_41456 & x_41457;
assign x_41459 = x_41455 & x_41458;
assign x_41460 = x_10169 & x_10170;
assign x_41461 = x_10171 & x_10172;
assign x_41462 = x_41460 & x_41461;
assign x_41463 = x_10173 & x_10174;
assign x_41464 = x_10175 & x_10176;
assign x_41465 = x_41463 & x_41464;
assign x_41466 = x_41462 & x_41465;
assign x_41467 = x_41459 & x_41466;
assign x_41468 = x_41453 & x_41467;
assign x_41469 = x_10178 & x_10179;
assign x_41470 = x_10177 & x_41469;
assign x_41471 = x_10180 & x_10181;
assign x_41472 = x_10182 & x_10183;
assign x_41473 = x_41471 & x_41472;
assign x_41474 = x_41470 & x_41473;
assign x_41475 = x_10184 & x_10185;
assign x_41476 = x_10186 & x_10187;
assign x_41477 = x_41475 & x_41476;
assign x_41478 = x_10188 & x_10189;
assign x_41479 = x_10190 & x_10191;
assign x_41480 = x_41478 & x_41479;
assign x_41481 = x_41477 & x_41480;
assign x_41482 = x_41474 & x_41481;
assign x_41483 = x_10192 & x_10193;
assign x_41484 = x_10194 & x_10195;
assign x_41485 = x_41483 & x_41484;
assign x_41486 = x_10196 & x_10197;
assign x_41487 = x_10198 & x_10199;
assign x_41488 = x_41486 & x_41487;
assign x_41489 = x_41485 & x_41488;
assign x_41490 = x_10200 & x_10201;
assign x_41491 = x_10202 & x_10203;
assign x_41492 = x_41490 & x_41491;
assign x_41493 = x_10204 & x_10205;
assign x_41494 = x_10206 & x_10207;
assign x_41495 = x_41493 & x_41494;
assign x_41496 = x_41492 & x_41495;
assign x_41497 = x_41489 & x_41496;
assign x_41498 = x_41482 & x_41497;
assign x_41499 = x_41468 & x_41498;
assign x_41500 = x_10209 & x_10210;
assign x_41501 = x_10208 & x_41500;
assign x_41502 = x_10211 & x_10212;
assign x_41503 = x_10213 & x_10214;
assign x_41504 = x_41502 & x_41503;
assign x_41505 = x_41501 & x_41504;
assign x_41506 = x_10215 & x_10216;
assign x_41507 = x_10217 & x_10218;
assign x_41508 = x_41506 & x_41507;
assign x_41509 = x_10219 & x_10220;
assign x_41510 = x_10221 & x_10222;
assign x_41511 = x_41509 & x_41510;
assign x_41512 = x_41508 & x_41511;
assign x_41513 = x_41505 & x_41512;
assign x_41514 = x_10223 & x_10224;
assign x_41515 = x_10225 & x_10226;
assign x_41516 = x_41514 & x_41515;
assign x_41517 = x_10227 & x_10228;
assign x_41518 = x_10229 & x_10230;
assign x_41519 = x_41517 & x_41518;
assign x_41520 = x_41516 & x_41519;
assign x_41521 = x_10231 & x_10232;
assign x_41522 = x_10233 & x_10234;
assign x_41523 = x_41521 & x_41522;
assign x_41524 = x_10235 & x_10236;
assign x_41525 = x_10237 & x_10238;
assign x_41526 = x_41524 & x_41525;
assign x_41527 = x_41523 & x_41526;
assign x_41528 = x_41520 & x_41527;
assign x_41529 = x_41513 & x_41528;
assign x_41530 = x_10240 & x_10241;
assign x_41531 = x_10239 & x_41530;
assign x_41532 = x_10242 & x_10243;
assign x_41533 = x_10244 & x_10245;
assign x_41534 = x_41532 & x_41533;
assign x_41535 = x_41531 & x_41534;
assign x_41536 = x_10246 & x_10247;
assign x_41537 = x_10248 & x_10249;
assign x_41538 = x_41536 & x_41537;
assign x_41539 = x_10250 & x_10251;
assign x_41540 = x_10252 & x_10253;
assign x_41541 = x_41539 & x_41540;
assign x_41542 = x_41538 & x_41541;
assign x_41543 = x_41535 & x_41542;
assign x_41544 = x_10254 & x_10255;
assign x_41545 = x_10256 & x_10257;
assign x_41546 = x_41544 & x_41545;
assign x_41547 = x_10258 & x_10259;
assign x_41548 = x_10260 & x_10261;
assign x_41549 = x_41547 & x_41548;
assign x_41550 = x_41546 & x_41549;
assign x_41551 = x_10262 & x_10263;
assign x_41552 = x_10264 & x_10265;
assign x_41553 = x_41551 & x_41552;
assign x_41554 = x_10266 & x_10267;
assign x_41555 = x_10268 & x_10269;
assign x_41556 = x_41554 & x_41555;
assign x_41557 = x_41553 & x_41556;
assign x_41558 = x_41550 & x_41557;
assign x_41559 = x_41543 & x_41558;
assign x_41560 = x_41529 & x_41559;
assign x_41561 = x_41499 & x_41560;
assign x_41562 = x_41439 & x_41561;
assign x_41563 = x_41318 & x_41562;
assign x_41564 = x_10271 & x_10272;
assign x_41565 = x_10270 & x_41564;
assign x_41566 = x_10273 & x_10274;
assign x_41567 = x_10275 & x_10276;
assign x_41568 = x_41566 & x_41567;
assign x_41569 = x_41565 & x_41568;
assign x_41570 = x_10277 & x_10278;
assign x_41571 = x_10279 & x_10280;
assign x_41572 = x_41570 & x_41571;
assign x_41573 = x_10281 & x_10282;
assign x_41574 = x_10283 & x_10284;
assign x_41575 = x_41573 & x_41574;
assign x_41576 = x_41572 & x_41575;
assign x_41577 = x_41569 & x_41576;
assign x_41578 = x_10286 & x_10287;
assign x_41579 = x_10285 & x_41578;
assign x_41580 = x_10288 & x_10289;
assign x_41581 = x_10290 & x_10291;
assign x_41582 = x_41580 & x_41581;
assign x_41583 = x_41579 & x_41582;
assign x_41584 = x_10292 & x_10293;
assign x_41585 = x_10294 & x_10295;
assign x_41586 = x_41584 & x_41585;
assign x_41587 = x_10296 & x_10297;
assign x_41588 = x_10298 & x_10299;
assign x_41589 = x_41587 & x_41588;
assign x_41590 = x_41586 & x_41589;
assign x_41591 = x_41583 & x_41590;
assign x_41592 = x_41577 & x_41591;
assign x_41593 = x_10301 & x_10302;
assign x_41594 = x_10300 & x_41593;
assign x_41595 = x_10303 & x_10304;
assign x_41596 = x_10305 & x_10306;
assign x_41597 = x_41595 & x_41596;
assign x_41598 = x_41594 & x_41597;
assign x_41599 = x_10307 & x_10308;
assign x_41600 = x_10309 & x_10310;
assign x_41601 = x_41599 & x_41600;
assign x_41602 = x_10311 & x_10312;
assign x_41603 = x_10313 & x_10314;
assign x_41604 = x_41602 & x_41603;
assign x_41605 = x_41601 & x_41604;
assign x_41606 = x_41598 & x_41605;
assign x_41607 = x_10315 & x_10316;
assign x_41608 = x_10317 & x_10318;
assign x_41609 = x_41607 & x_41608;
assign x_41610 = x_10319 & x_10320;
assign x_41611 = x_10321 & x_10322;
assign x_41612 = x_41610 & x_41611;
assign x_41613 = x_41609 & x_41612;
assign x_41614 = x_10323 & x_10324;
assign x_41615 = x_10325 & x_10326;
assign x_41616 = x_41614 & x_41615;
assign x_41617 = x_10327 & x_10328;
assign x_41618 = x_10329 & x_10330;
assign x_41619 = x_41617 & x_41618;
assign x_41620 = x_41616 & x_41619;
assign x_41621 = x_41613 & x_41620;
assign x_41622 = x_41606 & x_41621;
assign x_41623 = x_41592 & x_41622;
assign x_41624 = x_10332 & x_10333;
assign x_41625 = x_10331 & x_41624;
assign x_41626 = x_10334 & x_10335;
assign x_41627 = x_10336 & x_10337;
assign x_41628 = x_41626 & x_41627;
assign x_41629 = x_41625 & x_41628;
assign x_41630 = x_10338 & x_10339;
assign x_41631 = x_10340 & x_10341;
assign x_41632 = x_41630 & x_41631;
assign x_41633 = x_10342 & x_10343;
assign x_41634 = x_10344 & x_10345;
assign x_41635 = x_41633 & x_41634;
assign x_41636 = x_41632 & x_41635;
assign x_41637 = x_41629 & x_41636;
assign x_41638 = x_10347 & x_10348;
assign x_41639 = x_10346 & x_41638;
assign x_41640 = x_10349 & x_10350;
assign x_41641 = x_10351 & x_10352;
assign x_41642 = x_41640 & x_41641;
assign x_41643 = x_41639 & x_41642;
assign x_41644 = x_10353 & x_10354;
assign x_41645 = x_10355 & x_10356;
assign x_41646 = x_41644 & x_41645;
assign x_41647 = x_10357 & x_10358;
assign x_41648 = x_10359 & x_10360;
assign x_41649 = x_41647 & x_41648;
assign x_41650 = x_41646 & x_41649;
assign x_41651 = x_41643 & x_41650;
assign x_41652 = x_41637 & x_41651;
assign x_41653 = x_10362 & x_10363;
assign x_41654 = x_10361 & x_41653;
assign x_41655 = x_10364 & x_10365;
assign x_41656 = x_10366 & x_10367;
assign x_41657 = x_41655 & x_41656;
assign x_41658 = x_41654 & x_41657;
assign x_41659 = x_10368 & x_10369;
assign x_41660 = x_10370 & x_10371;
assign x_41661 = x_41659 & x_41660;
assign x_41662 = x_10372 & x_10373;
assign x_41663 = x_10374 & x_10375;
assign x_41664 = x_41662 & x_41663;
assign x_41665 = x_41661 & x_41664;
assign x_41666 = x_41658 & x_41665;
assign x_41667 = x_10376 & x_10377;
assign x_41668 = x_10378 & x_10379;
assign x_41669 = x_41667 & x_41668;
assign x_41670 = x_10380 & x_10381;
assign x_41671 = x_10382 & x_10383;
assign x_41672 = x_41670 & x_41671;
assign x_41673 = x_41669 & x_41672;
assign x_41674 = x_10384 & x_10385;
assign x_41675 = x_10386 & x_10387;
assign x_41676 = x_41674 & x_41675;
assign x_41677 = x_10388 & x_10389;
assign x_41678 = x_10390 & x_10391;
assign x_41679 = x_41677 & x_41678;
assign x_41680 = x_41676 & x_41679;
assign x_41681 = x_41673 & x_41680;
assign x_41682 = x_41666 & x_41681;
assign x_41683 = x_41652 & x_41682;
assign x_41684 = x_41623 & x_41683;
assign x_41685 = x_10393 & x_10394;
assign x_41686 = x_10392 & x_41685;
assign x_41687 = x_10395 & x_10396;
assign x_41688 = x_10397 & x_10398;
assign x_41689 = x_41687 & x_41688;
assign x_41690 = x_41686 & x_41689;
assign x_41691 = x_10399 & x_10400;
assign x_41692 = x_10401 & x_10402;
assign x_41693 = x_41691 & x_41692;
assign x_41694 = x_10403 & x_10404;
assign x_41695 = x_10405 & x_10406;
assign x_41696 = x_41694 & x_41695;
assign x_41697 = x_41693 & x_41696;
assign x_41698 = x_41690 & x_41697;
assign x_41699 = x_10408 & x_10409;
assign x_41700 = x_10407 & x_41699;
assign x_41701 = x_10410 & x_10411;
assign x_41702 = x_10412 & x_10413;
assign x_41703 = x_41701 & x_41702;
assign x_41704 = x_41700 & x_41703;
assign x_41705 = x_10414 & x_10415;
assign x_41706 = x_10416 & x_10417;
assign x_41707 = x_41705 & x_41706;
assign x_41708 = x_10418 & x_10419;
assign x_41709 = x_10420 & x_10421;
assign x_41710 = x_41708 & x_41709;
assign x_41711 = x_41707 & x_41710;
assign x_41712 = x_41704 & x_41711;
assign x_41713 = x_41698 & x_41712;
assign x_41714 = x_10423 & x_10424;
assign x_41715 = x_10422 & x_41714;
assign x_41716 = x_10425 & x_10426;
assign x_41717 = x_10427 & x_10428;
assign x_41718 = x_41716 & x_41717;
assign x_41719 = x_41715 & x_41718;
assign x_41720 = x_10429 & x_10430;
assign x_41721 = x_10431 & x_10432;
assign x_41722 = x_41720 & x_41721;
assign x_41723 = x_10433 & x_10434;
assign x_41724 = x_10435 & x_10436;
assign x_41725 = x_41723 & x_41724;
assign x_41726 = x_41722 & x_41725;
assign x_41727 = x_41719 & x_41726;
assign x_41728 = x_10437 & x_10438;
assign x_41729 = x_10439 & x_10440;
assign x_41730 = x_41728 & x_41729;
assign x_41731 = x_10441 & x_10442;
assign x_41732 = x_10443 & x_10444;
assign x_41733 = x_41731 & x_41732;
assign x_41734 = x_41730 & x_41733;
assign x_41735 = x_10445 & x_10446;
assign x_41736 = x_10447 & x_10448;
assign x_41737 = x_41735 & x_41736;
assign x_41738 = x_10449 & x_10450;
assign x_41739 = x_10451 & x_10452;
assign x_41740 = x_41738 & x_41739;
assign x_41741 = x_41737 & x_41740;
assign x_41742 = x_41734 & x_41741;
assign x_41743 = x_41727 & x_41742;
assign x_41744 = x_41713 & x_41743;
assign x_41745 = x_10454 & x_10455;
assign x_41746 = x_10453 & x_41745;
assign x_41747 = x_10456 & x_10457;
assign x_41748 = x_10458 & x_10459;
assign x_41749 = x_41747 & x_41748;
assign x_41750 = x_41746 & x_41749;
assign x_41751 = x_10460 & x_10461;
assign x_41752 = x_10462 & x_10463;
assign x_41753 = x_41751 & x_41752;
assign x_41754 = x_10464 & x_10465;
assign x_41755 = x_10466 & x_10467;
assign x_41756 = x_41754 & x_41755;
assign x_41757 = x_41753 & x_41756;
assign x_41758 = x_41750 & x_41757;
assign x_41759 = x_10469 & x_10470;
assign x_41760 = x_10468 & x_41759;
assign x_41761 = x_10471 & x_10472;
assign x_41762 = x_10473 & x_10474;
assign x_41763 = x_41761 & x_41762;
assign x_41764 = x_41760 & x_41763;
assign x_41765 = x_10475 & x_10476;
assign x_41766 = x_10477 & x_10478;
assign x_41767 = x_41765 & x_41766;
assign x_41768 = x_10479 & x_10480;
assign x_41769 = x_10481 & x_10482;
assign x_41770 = x_41768 & x_41769;
assign x_41771 = x_41767 & x_41770;
assign x_41772 = x_41764 & x_41771;
assign x_41773 = x_41758 & x_41772;
assign x_41774 = x_10484 & x_10485;
assign x_41775 = x_10483 & x_41774;
assign x_41776 = x_10486 & x_10487;
assign x_41777 = x_10488 & x_10489;
assign x_41778 = x_41776 & x_41777;
assign x_41779 = x_41775 & x_41778;
assign x_41780 = x_10490 & x_10491;
assign x_41781 = x_10492 & x_10493;
assign x_41782 = x_41780 & x_41781;
assign x_41783 = x_10494 & x_10495;
assign x_41784 = x_10496 & x_10497;
assign x_41785 = x_41783 & x_41784;
assign x_41786 = x_41782 & x_41785;
assign x_41787 = x_41779 & x_41786;
assign x_41788 = x_10498 & x_10499;
assign x_41789 = x_10500 & x_10501;
assign x_41790 = x_41788 & x_41789;
assign x_41791 = x_10502 & x_10503;
assign x_41792 = x_10504 & x_10505;
assign x_41793 = x_41791 & x_41792;
assign x_41794 = x_41790 & x_41793;
assign x_41795 = x_10506 & x_10507;
assign x_41796 = x_10508 & x_10509;
assign x_41797 = x_41795 & x_41796;
assign x_41798 = x_10510 & x_10511;
assign x_41799 = x_10512 & x_10513;
assign x_41800 = x_41798 & x_41799;
assign x_41801 = x_41797 & x_41800;
assign x_41802 = x_41794 & x_41801;
assign x_41803 = x_41787 & x_41802;
assign x_41804 = x_41773 & x_41803;
assign x_41805 = x_41744 & x_41804;
assign x_41806 = x_41684 & x_41805;
assign x_41807 = x_10515 & x_10516;
assign x_41808 = x_10514 & x_41807;
assign x_41809 = x_10517 & x_10518;
assign x_41810 = x_10519 & x_10520;
assign x_41811 = x_41809 & x_41810;
assign x_41812 = x_41808 & x_41811;
assign x_41813 = x_10521 & x_10522;
assign x_41814 = x_10523 & x_10524;
assign x_41815 = x_41813 & x_41814;
assign x_41816 = x_10525 & x_10526;
assign x_41817 = x_10527 & x_10528;
assign x_41818 = x_41816 & x_41817;
assign x_41819 = x_41815 & x_41818;
assign x_41820 = x_41812 & x_41819;
assign x_41821 = x_10530 & x_10531;
assign x_41822 = x_10529 & x_41821;
assign x_41823 = x_10532 & x_10533;
assign x_41824 = x_10534 & x_10535;
assign x_41825 = x_41823 & x_41824;
assign x_41826 = x_41822 & x_41825;
assign x_41827 = x_10536 & x_10537;
assign x_41828 = x_10538 & x_10539;
assign x_41829 = x_41827 & x_41828;
assign x_41830 = x_10540 & x_10541;
assign x_41831 = x_10542 & x_10543;
assign x_41832 = x_41830 & x_41831;
assign x_41833 = x_41829 & x_41832;
assign x_41834 = x_41826 & x_41833;
assign x_41835 = x_41820 & x_41834;
assign x_41836 = x_10545 & x_10546;
assign x_41837 = x_10544 & x_41836;
assign x_41838 = x_10547 & x_10548;
assign x_41839 = x_10549 & x_10550;
assign x_41840 = x_41838 & x_41839;
assign x_41841 = x_41837 & x_41840;
assign x_41842 = x_10551 & x_10552;
assign x_41843 = x_10553 & x_10554;
assign x_41844 = x_41842 & x_41843;
assign x_41845 = x_10555 & x_10556;
assign x_41846 = x_10557 & x_10558;
assign x_41847 = x_41845 & x_41846;
assign x_41848 = x_41844 & x_41847;
assign x_41849 = x_41841 & x_41848;
assign x_41850 = x_10559 & x_10560;
assign x_41851 = x_10561 & x_10562;
assign x_41852 = x_41850 & x_41851;
assign x_41853 = x_10563 & x_10564;
assign x_41854 = x_10565 & x_10566;
assign x_41855 = x_41853 & x_41854;
assign x_41856 = x_41852 & x_41855;
assign x_41857 = x_10567 & x_10568;
assign x_41858 = x_10569 & x_10570;
assign x_41859 = x_41857 & x_41858;
assign x_41860 = x_10571 & x_10572;
assign x_41861 = x_10573 & x_10574;
assign x_41862 = x_41860 & x_41861;
assign x_41863 = x_41859 & x_41862;
assign x_41864 = x_41856 & x_41863;
assign x_41865 = x_41849 & x_41864;
assign x_41866 = x_41835 & x_41865;
assign x_41867 = x_10576 & x_10577;
assign x_41868 = x_10575 & x_41867;
assign x_41869 = x_10578 & x_10579;
assign x_41870 = x_10580 & x_10581;
assign x_41871 = x_41869 & x_41870;
assign x_41872 = x_41868 & x_41871;
assign x_41873 = x_10582 & x_10583;
assign x_41874 = x_10584 & x_10585;
assign x_41875 = x_41873 & x_41874;
assign x_41876 = x_10586 & x_10587;
assign x_41877 = x_10588 & x_10589;
assign x_41878 = x_41876 & x_41877;
assign x_41879 = x_41875 & x_41878;
assign x_41880 = x_41872 & x_41879;
assign x_41881 = x_10591 & x_10592;
assign x_41882 = x_10590 & x_41881;
assign x_41883 = x_10593 & x_10594;
assign x_41884 = x_10595 & x_10596;
assign x_41885 = x_41883 & x_41884;
assign x_41886 = x_41882 & x_41885;
assign x_41887 = x_10597 & x_10598;
assign x_41888 = x_10599 & x_10600;
assign x_41889 = x_41887 & x_41888;
assign x_41890 = x_10601 & x_10602;
assign x_41891 = x_10603 & x_10604;
assign x_41892 = x_41890 & x_41891;
assign x_41893 = x_41889 & x_41892;
assign x_41894 = x_41886 & x_41893;
assign x_41895 = x_41880 & x_41894;
assign x_41896 = x_10606 & x_10607;
assign x_41897 = x_10605 & x_41896;
assign x_41898 = x_10608 & x_10609;
assign x_41899 = x_10610 & x_10611;
assign x_41900 = x_41898 & x_41899;
assign x_41901 = x_41897 & x_41900;
assign x_41902 = x_10612 & x_10613;
assign x_41903 = x_10614 & x_10615;
assign x_41904 = x_41902 & x_41903;
assign x_41905 = x_10616 & x_10617;
assign x_41906 = x_10618 & x_10619;
assign x_41907 = x_41905 & x_41906;
assign x_41908 = x_41904 & x_41907;
assign x_41909 = x_41901 & x_41908;
assign x_41910 = x_10620 & x_10621;
assign x_41911 = x_10622 & x_10623;
assign x_41912 = x_41910 & x_41911;
assign x_41913 = x_10624 & x_10625;
assign x_41914 = x_10626 & x_10627;
assign x_41915 = x_41913 & x_41914;
assign x_41916 = x_41912 & x_41915;
assign x_41917 = x_10628 & x_10629;
assign x_41918 = x_10630 & x_10631;
assign x_41919 = x_41917 & x_41918;
assign x_41920 = x_10632 & x_10633;
assign x_41921 = x_10634 & x_10635;
assign x_41922 = x_41920 & x_41921;
assign x_41923 = x_41919 & x_41922;
assign x_41924 = x_41916 & x_41923;
assign x_41925 = x_41909 & x_41924;
assign x_41926 = x_41895 & x_41925;
assign x_41927 = x_41866 & x_41926;
assign x_41928 = x_10637 & x_10638;
assign x_41929 = x_10636 & x_41928;
assign x_41930 = x_10639 & x_10640;
assign x_41931 = x_10641 & x_10642;
assign x_41932 = x_41930 & x_41931;
assign x_41933 = x_41929 & x_41932;
assign x_41934 = x_10643 & x_10644;
assign x_41935 = x_10645 & x_10646;
assign x_41936 = x_41934 & x_41935;
assign x_41937 = x_10647 & x_10648;
assign x_41938 = x_10649 & x_10650;
assign x_41939 = x_41937 & x_41938;
assign x_41940 = x_41936 & x_41939;
assign x_41941 = x_41933 & x_41940;
assign x_41942 = x_10652 & x_10653;
assign x_41943 = x_10651 & x_41942;
assign x_41944 = x_10654 & x_10655;
assign x_41945 = x_10656 & x_10657;
assign x_41946 = x_41944 & x_41945;
assign x_41947 = x_41943 & x_41946;
assign x_41948 = x_10658 & x_10659;
assign x_41949 = x_10660 & x_10661;
assign x_41950 = x_41948 & x_41949;
assign x_41951 = x_10662 & x_10663;
assign x_41952 = x_10664 & x_10665;
assign x_41953 = x_41951 & x_41952;
assign x_41954 = x_41950 & x_41953;
assign x_41955 = x_41947 & x_41954;
assign x_41956 = x_41941 & x_41955;
assign x_41957 = x_10667 & x_10668;
assign x_41958 = x_10666 & x_41957;
assign x_41959 = x_10669 & x_10670;
assign x_41960 = x_10671 & x_10672;
assign x_41961 = x_41959 & x_41960;
assign x_41962 = x_41958 & x_41961;
assign x_41963 = x_10673 & x_10674;
assign x_41964 = x_10675 & x_10676;
assign x_41965 = x_41963 & x_41964;
assign x_41966 = x_10677 & x_10678;
assign x_41967 = x_10679 & x_10680;
assign x_41968 = x_41966 & x_41967;
assign x_41969 = x_41965 & x_41968;
assign x_41970 = x_41962 & x_41969;
assign x_41971 = x_10681 & x_10682;
assign x_41972 = x_10683 & x_10684;
assign x_41973 = x_41971 & x_41972;
assign x_41974 = x_10685 & x_10686;
assign x_41975 = x_10687 & x_10688;
assign x_41976 = x_41974 & x_41975;
assign x_41977 = x_41973 & x_41976;
assign x_41978 = x_10689 & x_10690;
assign x_41979 = x_10691 & x_10692;
assign x_41980 = x_41978 & x_41979;
assign x_41981 = x_10693 & x_10694;
assign x_41982 = x_10695 & x_10696;
assign x_41983 = x_41981 & x_41982;
assign x_41984 = x_41980 & x_41983;
assign x_41985 = x_41977 & x_41984;
assign x_41986 = x_41970 & x_41985;
assign x_41987 = x_41956 & x_41986;
assign x_41988 = x_10698 & x_10699;
assign x_41989 = x_10697 & x_41988;
assign x_41990 = x_10700 & x_10701;
assign x_41991 = x_10702 & x_10703;
assign x_41992 = x_41990 & x_41991;
assign x_41993 = x_41989 & x_41992;
assign x_41994 = x_10704 & x_10705;
assign x_41995 = x_10706 & x_10707;
assign x_41996 = x_41994 & x_41995;
assign x_41997 = x_10708 & x_10709;
assign x_41998 = x_10710 & x_10711;
assign x_41999 = x_41997 & x_41998;
assign x_42000 = x_41996 & x_41999;
assign x_42001 = x_41993 & x_42000;
assign x_42002 = x_10712 & x_10713;
assign x_42003 = x_10714 & x_10715;
assign x_42004 = x_42002 & x_42003;
assign x_42005 = x_10716 & x_10717;
assign x_42006 = x_10718 & x_10719;
assign x_42007 = x_42005 & x_42006;
assign x_42008 = x_42004 & x_42007;
assign x_42009 = x_10720 & x_10721;
assign x_42010 = x_10722 & x_10723;
assign x_42011 = x_42009 & x_42010;
assign x_42012 = x_10724 & x_10725;
assign x_42013 = x_10726 & x_10727;
assign x_42014 = x_42012 & x_42013;
assign x_42015 = x_42011 & x_42014;
assign x_42016 = x_42008 & x_42015;
assign x_42017 = x_42001 & x_42016;
assign x_42018 = x_10729 & x_10730;
assign x_42019 = x_10728 & x_42018;
assign x_42020 = x_10731 & x_10732;
assign x_42021 = x_10733 & x_10734;
assign x_42022 = x_42020 & x_42021;
assign x_42023 = x_42019 & x_42022;
assign x_42024 = x_10735 & x_10736;
assign x_42025 = x_10737 & x_10738;
assign x_42026 = x_42024 & x_42025;
assign x_42027 = x_10739 & x_10740;
assign x_42028 = x_10741 & x_10742;
assign x_42029 = x_42027 & x_42028;
assign x_42030 = x_42026 & x_42029;
assign x_42031 = x_42023 & x_42030;
assign x_42032 = x_10743 & x_10744;
assign x_42033 = x_10745 & x_10746;
assign x_42034 = x_42032 & x_42033;
assign x_42035 = x_10747 & x_10748;
assign x_42036 = x_10749 & x_10750;
assign x_42037 = x_42035 & x_42036;
assign x_42038 = x_42034 & x_42037;
assign x_42039 = x_10751 & x_10752;
assign x_42040 = x_10753 & x_10754;
assign x_42041 = x_42039 & x_42040;
assign x_42042 = x_10755 & x_10756;
assign x_42043 = x_10757 & x_10758;
assign x_42044 = x_42042 & x_42043;
assign x_42045 = x_42041 & x_42044;
assign x_42046 = x_42038 & x_42045;
assign x_42047 = x_42031 & x_42046;
assign x_42048 = x_42017 & x_42047;
assign x_42049 = x_41987 & x_42048;
assign x_42050 = x_41927 & x_42049;
assign x_42051 = x_41806 & x_42050;
assign x_42052 = x_41563 & x_42051;
assign x_42053 = x_10760 & x_10761;
assign x_42054 = x_10759 & x_42053;
assign x_42055 = x_10762 & x_10763;
assign x_42056 = x_10764 & x_10765;
assign x_42057 = x_42055 & x_42056;
assign x_42058 = x_42054 & x_42057;
assign x_42059 = x_10766 & x_10767;
assign x_42060 = x_10768 & x_10769;
assign x_42061 = x_42059 & x_42060;
assign x_42062 = x_10770 & x_10771;
assign x_42063 = x_10772 & x_10773;
assign x_42064 = x_42062 & x_42063;
assign x_42065 = x_42061 & x_42064;
assign x_42066 = x_42058 & x_42065;
assign x_42067 = x_10775 & x_10776;
assign x_42068 = x_10774 & x_42067;
assign x_42069 = x_10777 & x_10778;
assign x_42070 = x_10779 & x_10780;
assign x_42071 = x_42069 & x_42070;
assign x_42072 = x_42068 & x_42071;
assign x_42073 = x_10781 & x_10782;
assign x_42074 = x_10783 & x_10784;
assign x_42075 = x_42073 & x_42074;
assign x_42076 = x_10785 & x_10786;
assign x_42077 = x_10787 & x_10788;
assign x_42078 = x_42076 & x_42077;
assign x_42079 = x_42075 & x_42078;
assign x_42080 = x_42072 & x_42079;
assign x_42081 = x_42066 & x_42080;
assign x_42082 = x_10790 & x_10791;
assign x_42083 = x_10789 & x_42082;
assign x_42084 = x_10792 & x_10793;
assign x_42085 = x_10794 & x_10795;
assign x_42086 = x_42084 & x_42085;
assign x_42087 = x_42083 & x_42086;
assign x_42088 = x_10796 & x_10797;
assign x_42089 = x_10798 & x_10799;
assign x_42090 = x_42088 & x_42089;
assign x_42091 = x_10800 & x_10801;
assign x_42092 = x_10802 & x_10803;
assign x_42093 = x_42091 & x_42092;
assign x_42094 = x_42090 & x_42093;
assign x_42095 = x_42087 & x_42094;
assign x_42096 = x_10804 & x_10805;
assign x_42097 = x_10806 & x_10807;
assign x_42098 = x_42096 & x_42097;
assign x_42099 = x_10808 & x_10809;
assign x_42100 = x_10810 & x_10811;
assign x_42101 = x_42099 & x_42100;
assign x_42102 = x_42098 & x_42101;
assign x_42103 = x_10812 & x_10813;
assign x_42104 = x_10814 & x_10815;
assign x_42105 = x_42103 & x_42104;
assign x_42106 = x_10816 & x_10817;
assign x_42107 = x_10818 & x_10819;
assign x_42108 = x_42106 & x_42107;
assign x_42109 = x_42105 & x_42108;
assign x_42110 = x_42102 & x_42109;
assign x_42111 = x_42095 & x_42110;
assign x_42112 = x_42081 & x_42111;
assign x_42113 = x_10821 & x_10822;
assign x_42114 = x_10820 & x_42113;
assign x_42115 = x_10823 & x_10824;
assign x_42116 = x_10825 & x_10826;
assign x_42117 = x_42115 & x_42116;
assign x_42118 = x_42114 & x_42117;
assign x_42119 = x_10827 & x_10828;
assign x_42120 = x_10829 & x_10830;
assign x_42121 = x_42119 & x_42120;
assign x_42122 = x_10831 & x_10832;
assign x_42123 = x_10833 & x_10834;
assign x_42124 = x_42122 & x_42123;
assign x_42125 = x_42121 & x_42124;
assign x_42126 = x_42118 & x_42125;
assign x_42127 = x_10836 & x_10837;
assign x_42128 = x_10835 & x_42127;
assign x_42129 = x_10838 & x_10839;
assign x_42130 = x_10840 & x_10841;
assign x_42131 = x_42129 & x_42130;
assign x_42132 = x_42128 & x_42131;
assign x_42133 = x_10842 & x_10843;
assign x_42134 = x_10844 & x_10845;
assign x_42135 = x_42133 & x_42134;
assign x_42136 = x_10846 & x_10847;
assign x_42137 = x_10848 & x_10849;
assign x_42138 = x_42136 & x_42137;
assign x_42139 = x_42135 & x_42138;
assign x_42140 = x_42132 & x_42139;
assign x_42141 = x_42126 & x_42140;
assign x_42142 = x_10851 & x_10852;
assign x_42143 = x_10850 & x_42142;
assign x_42144 = x_10853 & x_10854;
assign x_42145 = x_10855 & x_10856;
assign x_42146 = x_42144 & x_42145;
assign x_42147 = x_42143 & x_42146;
assign x_42148 = x_10857 & x_10858;
assign x_42149 = x_10859 & x_10860;
assign x_42150 = x_42148 & x_42149;
assign x_42151 = x_10861 & x_10862;
assign x_42152 = x_10863 & x_10864;
assign x_42153 = x_42151 & x_42152;
assign x_42154 = x_42150 & x_42153;
assign x_42155 = x_42147 & x_42154;
assign x_42156 = x_10865 & x_10866;
assign x_42157 = x_10867 & x_10868;
assign x_42158 = x_42156 & x_42157;
assign x_42159 = x_10869 & x_10870;
assign x_42160 = x_10871 & x_10872;
assign x_42161 = x_42159 & x_42160;
assign x_42162 = x_42158 & x_42161;
assign x_42163 = x_10873 & x_10874;
assign x_42164 = x_10875 & x_10876;
assign x_42165 = x_42163 & x_42164;
assign x_42166 = x_10877 & x_10878;
assign x_42167 = x_10879 & x_10880;
assign x_42168 = x_42166 & x_42167;
assign x_42169 = x_42165 & x_42168;
assign x_42170 = x_42162 & x_42169;
assign x_42171 = x_42155 & x_42170;
assign x_42172 = x_42141 & x_42171;
assign x_42173 = x_42112 & x_42172;
assign x_42174 = x_10882 & x_10883;
assign x_42175 = x_10881 & x_42174;
assign x_42176 = x_10884 & x_10885;
assign x_42177 = x_10886 & x_10887;
assign x_42178 = x_42176 & x_42177;
assign x_42179 = x_42175 & x_42178;
assign x_42180 = x_10888 & x_10889;
assign x_42181 = x_10890 & x_10891;
assign x_42182 = x_42180 & x_42181;
assign x_42183 = x_10892 & x_10893;
assign x_42184 = x_10894 & x_10895;
assign x_42185 = x_42183 & x_42184;
assign x_42186 = x_42182 & x_42185;
assign x_42187 = x_42179 & x_42186;
assign x_42188 = x_10897 & x_10898;
assign x_42189 = x_10896 & x_42188;
assign x_42190 = x_10899 & x_10900;
assign x_42191 = x_10901 & x_10902;
assign x_42192 = x_42190 & x_42191;
assign x_42193 = x_42189 & x_42192;
assign x_42194 = x_10903 & x_10904;
assign x_42195 = x_10905 & x_10906;
assign x_42196 = x_42194 & x_42195;
assign x_42197 = x_10907 & x_10908;
assign x_42198 = x_10909 & x_10910;
assign x_42199 = x_42197 & x_42198;
assign x_42200 = x_42196 & x_42199;
assign x_42201 = x_42193 & x_42200;
assign x_42202 = x_42187 & x_42201;
assign x_42203 = x_10912 & x_10913;
assign x_42204 = x_10911 & x_42203;
assign x_42205 = x_10914 & x_10915;
assign x_42206 = x_10916 & x_10917;
assign x_42207 = x_42205 & x_42206;
assign x_42208 = x_42204 & x_42207;
assign x_42209 = x_10918 & x_10919;
assign x_42210 = x_10920 & x_10921;
assign x_42211 = x_42209 & x_42210;
assign x_42212 = x_10922 & x_10923;
assign x_42213 = x_10924 & x_10925;
assign x_42214 = x_42212 & x_42213;
assign x_42215 = x_42211 & x_42214;
assign x_42216 = x_42208 & x_42215;
assign x_42217 = x_10926 & x_10927;
assign x_42218 = x_10928 & x_10929;
assign x_42219 = x_42217 & x_42218;
assign x_42220 = x_10930 & x_10931;
assign x_42221 = x_10932 & x_10933;
assign x_42222 = x_42220 & x_42221;
assign x_42223 = x_42219 & x_42222;
assign x_42224 = x_10934 & x_10935;
assign x_42225 = x_10936 & x_10937;
assign x_42226 = x_42224 & x_42225;
assign x_42227 = x_10938 & x_10939;
assign x_42228 = x_10940 & x_10941;
assign x_42229 = x_42227 & x_42228;
assign x_42230 = x_42226 & x_42229;
assign x_42231 = x_42223 & x_42230;
assign x_42232 = x_42216 & x_42231;
assign x_42233 = x_42202 & x_42232;
assign x_42234 = x_10943 & x_10944;
assign x_42235 = x_10942 & x_42234;
assign x_42236 = x_10945 & x_10946;
assign x_42237 = x_10947 & x_10948;
assign x_42238 = x_42236 & x_42237;
assign x_42239 = x_42235 & x_42238;
assign x_42240 = x_10949 & x_10950;
assign x_42241 = x_10951 & x_10952;
assign x_42242 = x_42240 & x_42241;
assign x_42243 = x_10953 & x_10954;
assign x_42244 = x_10955 & x_10956;
assign x_42245 = x_42243 & x_42244;
assign x_42246 = x_42242 & x_42245;
assign x_42247 = x_42239 & x_42246;
assign x_42248 = x_10958 & x_10959;
assign x_42249 = x_10957 & x_42248;
assign x_42250 = x_10960 & x_10961;
assign x_42251 = x_10962 & x_10963;
assign x_42252 = x_42250 & x_42251;
assign x_42253 = x_42249 & x_42252;
assign x_42254 = x_10964 & x_10965;
assign x_42255 = x_10966 & x_10967;
assign x_42256 = x_42254 & x_42255;
assign x_42257 = x_10968 & x_10969;
assign x_42258 = x_10970 & x_10971;
assign x_42259 = x_42257 & x_42258;
assign x_42260 = x_42256 & x_42259;
assign x_42261 = x_42253 & x_42260;
assign x_42262 = x_42247 & x_42261;
assign x_42263 = x_10973 & x_10974;
assign x_42264 = x_10972 & x_42263;
assign x_42265 = x_10975 & x_10976;
assign x_42266 = x_10977 & x_10978;
assign x_42267 = x_42265 & x_42266;
assign x_42268 = x_42264 & x_42267;
assign x_42269 = x_10979 & x_10980;
assign x_42270 = x_10981 & x_10982;
assign x_42271 = x_42269 & x_42270;
assign x_42272 = x_10983 & x_10984;
assign x_42273 = x_10985 & x_10986;
assign x_42274 = x_42272 & x_42273;
assign x_42275 = x_42271 & x_42274;
assign x_42276 = x_42268 & x_42275;
assign x_42277 = x_10987 & x_10988;
assign x_42278 = x_10989 & x_10990;
assign x_42279 = x_42277 & x_42278;
assign x_42280 = x_10991 & x_10992;
assign x_42281 = x_10993 & x_10994;
assign x_42282 = x_42280 & x_42281;
assign x_42283 = x_42279 & x_42282;
assign x_42284 = x_10995 & x_10996;
assign x_42285 = x_10997 & x_10998;
assign x_42286 = x_42284 & x_42285;
assign x_42287 = x_10999 & x_11000;
assign x_42288 = x_11001 & x_11002;
assign x_42289 = x_42287 & x_42288;
assign x_42290 = x_42286 & x_42289;
assign x_42291 = x_42283 & x_42290;
assign x_42292 = x_42276 & x_42291;
assign x_42293 = x_42262 & x_42292;
assign x_42294 = x_42233 & x_42293;
assign x_42295 = x_42173 & x_42294;
assign x_42296 = x_11004 & x_11005;
assign x_42297 = x_11003 & x_42296;
assign x_42298 = x_11006 & x_11007;
assign x_42299 = x_11008 & x_11009;
assign x_42300 = x_42298 & x_42299;
assign x_42301 = x_42297 & x_42300;
assign x_42302 = x_11010 & x_11011;
assign x_42303 = x_11012 & x_11013;
assign x_42304 = x_42302 & x_42303;
assign x_42305 = x_11014 & x_11015;
assign x_42306 = x_11016 & x_11017;
assign x_42307 = x_42305 & x_42306;
assign x_42308 = x_42304 & x_42307;
assign x_42309 = x_42301 & x_42308;
assign x_42310 = x_11019 & x_11020;
assign x_42311 = x_11018 & x_42310;
assign x_42312 = x_11021 & x_11022;
assign x_42313 = x_11023 & x_11024;
assign x_42314 = x_42312 & x_42313;
assign x_42315 = x_42311 & x_42314;
assign x_42316 = x_11025 & x_11026;
assign x_42317 = x_11027 & x_11028;
assign x_42318 = x_42316 & x_42317;
assign x_42319 = x_11029 & x_11030;
assign x_42320 = x_11031 & x_11032;
assign x_42321 = x_42319 & x_42320;
assign x_42322 = x_42318 & x_42321;
assign x_42323 = x_42315 & x_42322;
assign x_42324 = x_42309 & x_42323;
assign x_42325 = x_11034 & x_11035;
assign x_42326 = x_11033 & x_42325;
assign x_42327 = x_11036 & x_11037;
assign x_42328 = x_11038 & x_11039;
assign x_42329 = x_42327 & x_42328;
assign x_42330 = x_42326 & x_42329;
assign x_42331 = x_11040 & x_11041;
assign x_42332 = x_11042 & x_11043;
assign x_42333 = x_42331 & x_42332;
assign x_42334 = x_11044 & x_11045;
assign x_42335 = x_11046 & x_11047;
assign x_42336 = x_42334 & x_42335;
assign x_42337 = x_42333 & x_42336;
assign x_42338 = x_42330 & x_42337;
assign x_42339 = x_11048 & x_11049;
assign x_42340 = x_11050 & x_11051;
assign x_42341 = x_42339 & x_42340;
assign x_42342 = x_11052 & x_11053;
assign x_42343 = x_11054 & x_11055;
assign x_42344 = x_42342 & x_42343;
assign x_42345 = x_42341 & x_42344;
assign x_42346 = x_11056 & x_11057;
assign x_42347 = x_11058 & x_11059;
assign x_42348 = x_42346 & x_42347;
assign x_42349 = x_11060 & x_11061;
assign x_42350 = x_11062 & x_11063;
assign x_42351 = x_42349 & x_42350;
assign x_42352 = x_42348 & x_42351;
assign x_42353 = x_42345 & x_42352;
assign x_42354 = x_42338 & x_42353;
assign x_42355 = x_42324 & x_42354;
assign x_42356 = x_11065 & x_11066;
assign x_42357 = x_11064 & x_42356;
assign x_42358 = x_11067 & x_11068;
assign x_42359 = x_11069 & x_11070;
assign x_42360 = x_42358 & x_42359;
assign x_42361 = x_42357 & x_42360;
assign x_42362 = x_11071 & x_11072;
assign x_42363 = x_11073 & x_11074;
assign x_42364 = x_42362 & x_42363;
assign x_42365 = x_11075 & x_11076;
assign x_42366 = x_11077 & x_11078;
assign x_42367 = x_42365 & x_42366;
assign x_42368 = x_42364 & x_42367;
assign x_42369 = x_42361 & x_42368;
assign x_42370 = x_11080 & x_11081;
assign x_42371 = x_11079 & x_42370;
assign x_42372 = x_11082 & x_11083;
assign x_42373 = x_11084 & x_11085;
assign x_42374 = x_42372 & x_42373;
assign x_42375 = x_42371 & x_42374;
assign x_42376 = x_11086 & x_11087;
assign x_42377 = x_11088 & x_11089;
assign x_42378 = x_42376 & x_42377;
assign x_42379 = x_11090 & x_11091;
assign x_42380 = x_11092 & x_11093;
assign x_42381 = x_42379 & x_42380;
assign x_42382 = x_42378 & x_42381;
assign x_42383 = x_42375 & x_42382;
assign x_42384 = x_42369 & x_42383;
assign x_42385 = x_11095 & x_11096;
assign x_42386 = x_11094 & x_42385;
assign x_42387 = x_11097 & x_11098;
assign x_42388 = x_11099 & x_11100;
assign x_42389 = x_42387 & x_42388;
assign x_42390 = x_42386 & x_42389;
assign x_42391 = x_11101 & x_11102;
assign x_42392 = x_11103 & x_11104;
assign x_42393 = x_42391 & x_42392;
assign x_42394 = x_11105 & x_11106;
assign x_42395 = x_11107 & x_11108;
assign x_42396 = x_42394 & x_42395;
assign x_42397 = x_42393 & x_42396;
assign x_42398 = x_42390 & x_42397;
assign x_42399 = x_11109 & x_11110;
assign x_42400 = x_11111 & x_11112;
assign x_42401 = x_42399 & x_42400;
assign x_42402 = x_11113 & x_11114;
assign x_42403 = x_11115 & x_11116;
assign x_42404 = x_42402 & x_42403;
assign x_42405 = x_42401 & x_42404;
assign x_42406 = x_11117 & x_11118;
assign x_42407 = x_11119 & x_11120;
assign x_42408 = x_42406 & x_42407;
assign x_42409 = x_11121 & x_11122;
assign x_42410 = x_11123 & x_11124;
assign x_42411 = x_42409 & x_42410;
assign x_42412 = x_42408 & x_42411;
assign x_42413 = x_42405 & x_42412;
assign x_42414 = x_42398 & x_42413;
assign x_42415 = x_42384 & x_42414;
assign x_42416 = x_42355 & x_42415;
assign x_42417 = x_11126 & x_11127;
assign x_42418 = x_11125 & x_42417;
assign x_42419 = x_11128 & x_11129;
assign x_42420 = x_11130 & x_11131;
assign x_42421 = x_42419 & x_42420;
assign x_42422 = x_42418 & x_42421;
assign x_42423 = x_11132 & x_11133;
assign x_42424 = x_11134 & x_11135;
assign x_42425 = x_42423 & x_42424;
assign x_42426 = x_11136 & x_11137;
assign x_42427 = x_11138 & x_11139;
assign x_42428 = x_42426 & x_42427;
assign x_42429 = x_42425 & x_42428;
assign x_42430 = x_42422 & x_42429;
assign x_42431 = x_11141 & x_11142;
assign x_42432 = x_11140 & x_42431;
assign x_42433 = x_11143 & x_11144;
assign x_42434 = x_11145 & x_11146;
assign x_42435 = x_42433 & x_42434;
assign x_42436 = x_42432 & x_42435;
assign x_42437 = x_11147 & x_11148;
assign x_42438 = x_11149 & x_11150;
assign x_42439 = x_42437 & x_42438;
assign x_42440 = x_11151 & x_11152;
assign x_42441 = x_11153 & x_11154;
assign x_42442 = x_42440 & x_42441;
assign x_42443 = x_42439 & x_42442;
assign x_42444 = x_42436 & x_42443;
assign x_42445 = x_42430 & x_42444;
assign x_42446 = x_11156 & x_11157;
assign x_42447 = x_11155 & x_42446;
assign x_42448 = x_11158 & x_11159;
assign x_42449 = x_11160 & x_11161;
assign x_42450 = x_42448 & x_42449;
assign x_42451 = x_42447 & x_42450;
assign x_42452 = x_11162 & x_11163;
assign x_42453 = x_11164 & x_11165;
assign x_42454 = x_42452 & x_42453;
assign x_42455 = x_11166 & x_11167;
assign x_42456 = x_11168 & x_11169;
assign x_42457 = x_42455 & x_42456;
assign x_42458 = x_42454 & x_42457;
assign x_42459 = x_42451 & x_42458;
assign x_42460 = x_11170 & x_11171;
assign x_42461 = x_11172 & x_11173;
assign x_42462 = x_42460 & x_42461;
assign x_42463 = x_11174 & x_11175;
assign x_42464 = x_11176 & x_11177;
assign x_42465 = x_42463 & x_42464;
assign x_42466 = x_42462 & x_42465;
assign x_42467 = x_11178 & x_11179;
assign x_42468 = x_11180 & x_11181;
assign x_42469 = x_42467 & x_42468;
assign x_42470 = x_11182 & x_11183;
assign x_42471 = x_11184 & x_11185;
assign x_42472 = x_42470 & x_42471;
assign x_42473 = x_42469 & x_42472;
assign x_42474 = x_42466 & x_42473;
assign x_42475 = x_42459 & x_42474;
assign x_42476 = x_42445 & x_42475;
assign x_42477 = x_11187 & x_11188;
assign x_42478 = x_11186 & x_42477;
assign x_42479 = x_11189 & x_11190;
assign x_42480 = x_11191 & x_11192;
assign x_42481 = x_42479 & x_42480;
assign x_42482 = x_42478 & x_42481;
assign x_42483 = x_11193 & x_11194;
assign x_42484 = x_11195 & x_11196;
assign x_42485 = x_42483 & x_42484;
assign x_42486 = x_11197 & x_11198;
assign x_42487 = x_11199 & x_11200;
assign x_42488 = x_42486 & x_42487;
assign x_42489 = x_42485 & x_42488;
assign x_42490 = x_42482 & x_42489;
assign x_42491 = x_11201 & x_11202;
assign x_42492 = x_11203 & x_11204;
assign x_42493 = x_42491 & x_42492;
assign x_42494 = x_11205 & x_11206;
assign x_42495 = x_11207 & x_11208;
assign x_42496 = x_42494 & x_42495;
assign x_42497 = x_42493 & x_42496;
assign x_42498 = x_11209 & x_11210;
assign x_42499 = x_11211 & x_11212;
assign x_42500 = x_42498 & x_42499;
assign x_42501 = x_11213 & x_11214;
assign x_42502 = x_11215 & x_11216;
assign x_42503 = x_42501 & x_42502;
assign x_42504 = x_42500 & x_42503;
assign x_42505 = x_42497 & x_42504;
assign x_42506 = x_42490 & x_42505;
assign x_42507 = x_11218 & x_11219;
assign x_42508 = x_11217 & x_42507;
assign x_42509 = x_11220 & x_11221;
assign x_42510 = x_11222 & x_11223;
assign x_42511 = x_42509 & x_42510;
assign x_42512 = x_42508 & x_42511;
assign x_42513 = x_11224 & x_11225;
assign x_42514 = x_11226 & x_11227;
assign x_42515 = x_42513 & x_42514;
assign x_42516 = x_11228 & x_11229;
assign x_42517 = x_11230 & x_11231;
assign x_42518 = x_42516 & x_42517;
assign x_42519 = x_42515 & x_42518;
assign x_42520 = x_42512 & x_42519;
assign x_42521 = x_11232 & x_11233;
assign x_42522 = x_11234 & x_11235;
assign x_42523 = x_42521 & x_42522;
assign x_42524 = x_11236 & x_11237;
assign x_42525 = x_11238 & x_11239;
assign x_42526 = x_42524 & x_42525;
assign x_42527 = x_42523 & x_42526;
assign x_42528 = x_11240 & x_11241;
assign x_42529 = x_11242 & x_11243;
assign x_42530 = x_42528 & x_42529;
assign x_42531 = x_11244 & x_11245;
assign x_42532 = x_11246 & x_11247;
assign x_42533 = x_42531 & x_42532;
assign x_42534 = x_42530 & x_42533;
assign x_42535 = x_42527 & x_42534;
assign x_42536 = x_42520 & x_42535;
assign x_42537 = x_42506 & x_42536;
assign x_42538 = x_42476 & x_42537;
assign x_42539 = x_42416 & x_42538;
assign x_42540 = x_42295 & x_42539;
assign x_42541 = x_11249 & x_11250;
assign x_42542 = x_11248 & x_42541;
assign x_42543 = x_11251 & x_11252;
assign x_42544 = x_11253 & x_11254;
assign x_42545 = x_42543 & x_42544;
assign x_42546 = x_42542 & x_42545;
assign x_42547 = x_11255 & x_11256;
assign x_42548 = x_11257 & x_11258;
assign x_42549 = x_42547 & x_42548;
assign x_42550 = x_11259 & x_11260;
assign x_42551 = x_11261 & x_11262;
assign x_42552 = x_42550 & x_42551;
assign x_42553 = x_42549 & x_42552;
assign x_42554 = x_42546 & x_42553;
assign x_42555 = x_11264 & x_11265;
assign x_42556 = x_11263 & x_42555;
assign x_42557 = x_11266 & x_11267;
assign x_42558 = x_11268 & x_11269;
assign x_42559 = x_42557 & x_42558;
assign x_42560 = x_42556 & x_42559;
assign x_42561 = x_11270 & x_11271;
assign x_42562 = x_11272 & x_11273;
assign x_42563 = x_42561 & x_42562;
assign x_42564 = x_11274 & x_11275;
assign x_42565 = x_11276 & x_11277;
assign x_42566 = x_42564 & x_42565;
assign x_42567 = x_42563 & x_42566;
assign x_42568 = x_42560 & x_42567;
assign x_42569 = x_42554 & x_42568;
assign x_42570 = x_11279 & x_11280;
assign x_42571 = x_11278 & x_42570;
assign x_42572 = x_11281 & x_11282;
assign x_42573 = x_11283 & x_11284;
assign x_42574 = x_42572 & x_42573;
assign x_42575 = x_42571 & x_42574;
assign x_42576 = x_11285 & x_11286;
assign x_42577 = x_11287 & x_11288;
assign x_42578 = x_42576 & x_42577;
assign x_42579 = x_11289 & x_11290;
assign x_42580 = x_11291 & x_11292;
assign x_42581 = x_42579 & x_42580;
assign x_42582 = x_42578 & x_42581;
assign x_42583 = x_42575 & x_42582;
assign x_42584 = x_11293 & x_11294;
assign x_42585 = x_11295 & x_11296;
assign x_42586 = x_42584 & x_42585;
assign x_42587 = x_11297 & x_11298;
assign x_42588 = x_11299 & x_11300;
assign x_42589 = x_42587 & x_42588;
assign x_42590 = x_42586 & x_42589;
assign x_42591 = x_11301 & x_11302;
assign x_42592 = x_11303 & x_11304;
assign x_42593 = x_42591 & x_42592;
assign x_42594 = x_11305 & x_11306;
assign x_42595 = x_11307 & x_11308;
assign x_42596 = x_42594 & x_42595;
assign x_42597 = x_42593 & x_42596;
assign x_42598 = x_42590 & x_42597;
assign x_42599 = x_42583 & x_42598;
assign x_42600 = x_42569 & x_42599;
assign x_42601 = x_11310 & x_11311;
assign x_42602 = x_11309 & x_42601;
assign x_42603 = x_11312 & x_11313;
assign x_42604 = x_11314 & x_11315;
assign x_42605 = x_42603 & x_42604;
assign x_42606 = x_42602 & x_42605;
assign x_42607 = x_11316 & x_11317;
assign x_42608 = x_11318 & x_11319;
assign x_42609 = x_42607 & x_42608;
assign x_42610 = x_11320 & x_11321;
assign x_42611 = x_11322 & x_11323;
assign x_42612 = x_42610 & x_42611;
assign x_42613 = x_42609 & x_42612;
assign x_42614 = x_42606 & x_42613;
assign x_42615 = x_11325 & x_11326;
assign x_42616 = x_11324 & x_42615;
assign x_42617 = x_11327 & x_11328;
assign x_42618 = x_11329 & x_11330;
assign x_42619 = x_42617 & x_42618;
assign x_42620 = x_42616 & x_42619;
assign x_42621 = x_11331 & x_11332;
assign x_42622 = x_11333 & x_11334;
assign x_42623 = x_42621 & x_42622;
assign x_42624 = x_11335 & x_11336;
assign x_42625 = x_11337 & x_11338;
assign x_42626 = x_42624 & x_42625;
assign x_42627 = x_42623 & x_42626;
assign x_42628 = x_42620 & x_42627;
assign x_42629 = x_42614 & x_42628;
assign x_42630 = x_11340 & x_11341;
assign x_42631 = x_11339 & x_42630;
assign x_42632 = x_11342 & x_11343;
assign x_42633 = x_11344 & x_11345;
assign x_42634 = x_42632 & x_42633;
assign x_42635 = x_42631 & x_42634;
assign x_42636 = x_11346 & x_11347;
assign x_42637 = x_11348 & x_11349;
assign x_42638 = x_42636 & x_42637;
assign x_42639 = x_11350 & x_11351;
assign x_42640 = x_11352 & x_11353;
assign x_42641 = x_42639 & x_42640;
assign x_42642 = x_42638 & x_42641;
assign x_42643 = x_42635 & x_42642;
assign x_42644 = x_11354 & x_11355;
assign x_42645 = x_11356 & x_11357;
assign x_42646 = x_42644 & x_42645;
assign x_42647 = x_11358 & x_11359;
assign x_42648 = x_11360 & x_11361;
assign x_42649 = x_42647 & x_42648;
assign x_42650 = x_42646 & x_42649;
assign x_42651 = x_11362 & x_11363;
assign x_42652 = x_11364 & x_11365;
assign x_42653 = x_42651 & x_42652;
assign x_42654 = x_11366 & x_11367;
assign x_42655 = x_11368 & x_11369;
assign x_42656 = x_42654 & x_42655;
assign x_42657 = x_42653 & x_42656;
assign x_42658 = x_42650 & x_42657;
assign x_42659 = x_42643 & x_42658;
assign x_42660 = x_42629 & x_42659;
assign x_42661 = x_42600 & x_42660;
assign x_42662 = x_11371 & x_11372;
assign x_42663 = x_11370 & x_42662;
assign x_42664 = x_11373 & x_11374;
assign x_42665 = x_11375 & x_11376;
assign x_42666 = x_42664 & x_42665;
assign x_42667 = x_42663 & x_42666;
assign x_42668 = x_11377 & x_11378;
assign x_42669 = x_11379 & x_11380;
assign x_42670 = x_42668 & x_42669;
assign x_42671 = x_11381 & x_11382;
assign x_42672 = x_11383 & x_11384;
assign x_42673 = x_42671 & x_42672;
assign x_42674 = x_42670 & x_42673;
assign x_42675 = x_42667 & x_42674;
assign x_42676 = x_11386 & x_11387;
assign x_42677 = x_11385 & x_42676;
assign x_42678 = x_11388 & x_11389;
assign x_42679 = x_11390 & x_11391;
assign x_42680 = x_42678 & x_42679;
assign x_42681 = x_42677 & x_42680;
assign x_42682 = x_11392 & x_11393;
assign x_42683 = x_11394 & x_11395;
assign x_42684 = x_42682 & x_42683;
assign x_42685 = x_11396 & x_11397;
assign x_42686 = x_11398 & x_11399;
assign x_42687 = x_42685 & x_42686;
assign x_42688 = x_42684 & x_42687;
assign x_42689 = x_42681 & x_42688;
assign x_42690 = x_42675 & x_42689;
assign x_42691 = x_11401 & x_11402;
assign x_42692 = x_11400 & x_42691;
assign x_42693 = x_11403 & x_11404;
assign x_42694 = x_11405 & x_11406;
assign x_42695 = x_42693 & x_42694;
assign x_42696 = x_42692 & x_42695;
assign x_42697 = x_11407 & x_11408;
assign x_42698 = x_11409 & x_11410;
assign x_42699 = x_42697 & x_42698;
assign x_42700 = x_11411 & x_11412;
assign x_42701 = x_11413 & x_11414;
assign x_42702 = x_42700 & x_42701;
assign x_42703 = x_42699 & x_42702;
assign x_42704 = x_42696 & x_42703;
assign x_42705 = x_11415 & x_11416;
assign x_42706 = x_11417 & x_11418;
assign x_42707 = x_42705 & x_42706;
assign x_42708 = x_11419 & x_11420;
assign x_42709 = x_11421 & x_11422;
assign x_42710 = x_42708 & x_42709;
assign x_42711 = x_42707 & x_42710;
assign x_42712 = x_11423 & x_11424;
assign x_42713 = x_11425 & x_11426;
assign x_42714 = x_42712 & x_42713;
assign x_42715 = x_11427 & x_11428;
assign x_42716 = x_11429 & x_11430;
assign x_42717 = x_42715 & x_42716;
assign x_42718 = x_42714 & x_42717;
assign x_42719 = x_42711 & x_42718;
assign x_42720 = x_42704 & x_42719;
assign x_42721 = x_42690 & x_42720;
assign x_42722 = x_11432 & x_11433;
assign x_42723 = x_11431 & x_42722;
assign x_42724 = x_11434 & x_11435;
assign x_42725 = x_11436 & x_11437;
assign x_42726 = x_42724 & x_42725;
assign x_42727 = x_42723 & x_42726;
assign x_42728 = x_11438 & x_11439;
assign x_42729 = x_11440 & x_11441;
assign x_42730 = x_42728 & x_42729;
assign x_42731 = x_11442 & x_11443;
assign x_42732 = x_11444 & x_11445;
assign x_42733 = x_42731 & x_42732;
assign x_42734 = x_42730 & x_42733;
assign x_42735 = x_42727 & x_42734;
assign x_42736 = x_11447 & x_11448;
assign x_42737 = x_11446 & x_42736;
assign x_42738 = x_11449 & x_11450;
assign x_42739 = x_11451 & x_11452;
assign x_42740 = x_42738 & x_42739;
assign x_42741 = x_42737 & x_42740;
assign x_42742 = x_11453 & x_11454;
assign x_42743 = x_11455 & x_11456;
assign x_42744 = x_42742 & x_42743;
assign x_42745 = x_11457 & x_11458;
assign x_42746 = x_11459 & x_11460;
assign x_42747 = x_42745 & x_42746;
assign x_42748 = x_42744 & x_42747;
assign x_42749 = x_42741 & x_42748;
assign x_42750 = x_42735 & x_42749;
assign x_42751 = x_11462 & x_11463;
assign x_42752 = x_11461 & x_42751;
assign x_42753 = x_11464 & x_11465;
assign x_42754 = x_11466 & x_11467;
assign x_42755 = x_42753 & x_42754;
assign x_42756 = x_42752 & x_42755;
assign x_42757 = x_11468 & x_11469;
assign x_42758 = x_11470 & x_11471;
assign x_42759 = x_42757 & x_42758;
assign x_42760 = x_11472 & x_11473;
assign x_42761 = x_11474 & x_11475;
assign x_42762 = x_42760 & x_42761;
assign x_42763 = x_42759 & x_42762;
assign x_42764 = x_42756 & x_42763;
assign x_42765 = x_11476 & x_11477;
assign x_42766 = x_11478 & x_11479;
assign x_42767 = x_42765 & x_42766;
assign x_42768 = x_11480 & x_11481;
assign x_42769 = x_11482 & x_11483;
assign x_42770 = x_42768 & x_42769;
assign x_42771 = x_42767 & x_42770;
assign x_42772 = x_11484 & x_11485;
assign x_42773 = x_11486 & x_11487;
assign x_42774 = x_42772 & x_42773;
assign x_42775 = x_11488 & x_11489;
assign x_42776 = x_11490 & x_11491;
assign x_42777 = x_42775 & x_42776;
assign x_42778 = x_42774 & x_42777;
assign x_42779 = x_42771 & x_42778;
assign x_42780 = x_42764 & x_42779;
assign x_42781 = x_42750 & x_42780;
assign x_42782 = x_42721 & x_42781;
assign x_42783 = x_42661 & x_42782;
assign x_42784 = x_11493 & x_11494;
assign x_42785 = x_11492 & x_42784;
assign x_42786 = x_11495 & x_11496;
assign x_42787 = x_11497 & x_11498;
assign x_42788 = x_42786 & x_42787;
assign x_42789 = x_42785 & x_42788;
assign x_42790 = x_11499 & x_11500;
assign x_42791 = x_11501 & x_11502;
assign x_42792 = x_42790 & x_42791;
assign x_42793 = x_11503 & x_11504;
assign x_42794 = x_11505 & x_11506;
assign x_42795 = x_42793 & x_42794;
assign x_42796 = x_42792 & x_42795;
assign x_42797 = x_42789 & x_42796;
assign x_42798 = x_11508 & x_11509;
assign x_42799 = x_11507 & x_42798;
assign x_42800 = x_11510 & x_11511;
assign x_42801 = x_11512 & x_11513;
assign x_42802 = x_42800 & x_42801;
assign x_42803 = x_42799 & x_42802;
assign x_42804 = x_11514 & x_11515;
assign x_42805 = x_11516 & x_11517;
assign x_42806 = x_42804 & x_42805;
assign x_42807 = x_11518 & x_11519;
assign x_42808 = x_11520 & x_11521;
assign x_42809 = x_42807 & x_42808;
assign x_42810 = x_42806 & x_42809;
assign x_42811 = x_42803 & x_42810;
assign x_42812 = x_42797 & x_42811;
assign x_42813 = x_11523 & x_11524;
assign x_42814 = x_11522 & x_42813;
assign x_42815 = x_11525 & x_11526;
assign x_42816 = x_11527 & x_11528;
assign x_42817 = x_42815 & x_42816;
assign x_42818 = x_42814 & x_42817;
assign x_42819 = x_11529 & x_11530;
assign x_42820 = x_11531 & x_11532;
assign x_42821 = x_42819 & x_42820;
assign x_42822 = x_11533 & x_11534;
assign x_42823 = x_11535 & x_11536;
assign x_42824 = x_42822 & x_42823;
assign x_42825 = x_42821 & x_42824;
assign x_42826 = x_42818 & x_42825;
assign x_42827 = x_11537 & x_11538;
assign x_42828 = x_11539 & x_11540;
assign x_42829 = x_42827 & x_42828;
assign x_42830 = x_11541 & x_11542;
assign x_42831 = x_11543 & x_11544;
assign x_42832 = x_42830 & x_42831;
assign x_42833 = x_42829 & x_42832;
assign x_42834 = x_11545 & x_11546;
assign x_42835 = x_11547 & x_11548;
assign x_42836 = x_42834 & x_42835;
assign x_42837 = x_11549 & x_11550;
assign x_42838 = x_11551 & x_11552;
assign x_42839 = x_42837 & x_42838;
assign x_42840 = x_42836 & x_42839;
assign x_42841 = x_42833 & x_42840;
assign x_42842 = x_42826 & x_42841;
assign x_42843 = x_42812 & x_42842;
assign x_42844 = x_11554 & x_11555;
assign x_42845 = x_11553 & x_42844;
assign x_42846 = x_11556 & x_11557;
assign x_42847 = x_11558 & x_11559;
assign x_42848 = x_42846 & x_42847;
assign x_42849 = x_42845 & x_42848;
assign x_42850 = x_11560 & x_11561;
assign x_42851 = x_11562 & x_11563;
assign x_42852 = x_42850 & x_42851;
assign x_42853 = x_11564 & x_11565;
assign x_42854 = x_11566 & x_11567;
assign x_42855 = x_42853 & x_42854;
assign x_42856 = x_42852 & x_42855;
assign x_42857 = x_42849 & x_42856;
assign x_42858 = x_11569 & x_11570;
assign x_42859 = x_11568 & x_42858;
assign x_42860 = x_11571 & x_11572;
assign x_42861 = x_11573 & x_11574;
assign x_42862 = x_42860 & x_42861;
assign x_42863 = x_42859 & x_42862;
assign x_42864 = x_11575 & x_11576;
assign x_42865 = x_11577 & x_11578;
assign x_42866 = x_42864 & x_42865;
assign x_42867 = x_11579 & x_11580;
assign x_42868 = x_11581 & x_11582;
assign x_42869 = x_42867 & x_42868;
assign x_42870 = x_42866 & x_42869;
assign x_42871 = x_42863 & x_42870;
assign x_42872 = x_42857 & x_42871;
assign x_42873 = x_11584 & x_11585;
assign x_42874 = x_11583 & x_42873;
assign x_42875 = x_11586 & x_11587;
assign x_42876 = x_11588 & x_11589;
assign x_42877 = x_42875 & x_42876;
assign x_42878 = x_42874 & x_42877;
assign x_42879 = x_11590 & x_11591;
assign x_42880 = x_11592 & x_11593;
assign x_42881 = x_42879 & x_42880;
assign x_42882 = x_11594 & x_11595;
assign x_42883 = x_11596 & x_11597;
assign x_42884 = x_42882 & x_42883;
assign x_42885 = x_42881 & x_42884;
assign x_42886 = x_42878 & x_42885;
assign x_42887 = x_11598 & x_11599;
assign x_42888 = x_11600 & x_11601;
assign x_42889 = x_42887 & x_42888;
assign x_42890 = x_11602 & x_11603;
assign x_42891 = x_11604 & x_11605;
assign x_42892 = x_42890 & x_42891;
assign x_42893 = x_42889 & x_42892;
assign x_42894 = x_11606 & x_11607;
assign x_42895 = x_11608 & x_11609;
assign x_42896 = x_42894 & x_42895;
assign x_42897 = x_11610 & x_11611;
assign x_42898 = x_11612 & x_11613;
assign x_42899 = x_42897 & x_42898;
assign x_42900 = x_42896 & x_42899;
assign x_42901 = x_42893 & x_42900;
assign x_42902 = x_42886 & x_42901;
assign x_42903 = x_42872 & x_42902;
assign x_42904 = x_42843 & x_42903;
assign x_42905 = x_11615 & x_11616;
assign x_42906 = x_11614 & x_42905;
assign x_42907 = x_11617 & x_11618;
assign x_42908 = x_11619 & x_11620;
assign x_42909 = x_42907 & x_42908;
assign x_42910 = x_42906 & x_42909;
assign x_42911 = x_11621 & x_11622;
assign x_42912 = x_11623 & x_11624;
assign x_42913 = x_42911 & x_42912;
assign x_42914 = x_11625 & x_11626;
assign x_42915 = x_11627 & x_11628;
assign x_42916 = x_42914 & x_42915;
assign x_42917 = x_42913 & x_42916;
assign x_42918 = x_42910 & x_42917;
assign x_42919 = x_11630 & x_11631;
assign x_42920 = x_11629 & x_42919;
assign x_42921 = x_11632 & x_11633;
assign x_42922 = x_11634 & x_11635;
assign x_42923 = x_42921 & x_42922;
assign x_42924 = x_42920 & x_42923;
assign x_42925 = x_11636 & x_11637;
assign x_42926 = x_11638 & x_11639;
assign x_42927 = x_42925 & x_42926;
assign x_42928 = x_11640 & x_11641;
assign x_42929 = x_11642 & x_11643;
assign x_42930 = x_42928 & x_42929;
assign x_42931 = x_42927 & x_42930;
assign x_42932 = x_42924 & x_42931;
assign x_42933 = x_42918 & x_42932;
assign x_42934 = x_11645 & x_11646;
assign x_42935 = x_11644 & x_42934;
assign x_42936 = x_11647 & x_11648;
assign x_42937 = x_11649 & x_11650;
assign x_42938 = x_42936 & x_42937;
assign x_42939 = x_42935 & x_42938;
assign x_42940 = x_11651 & x_11652;
assign x_42941 = x_11653 & x_11654;
assign x_42942 = x_42940 & x_42941;
assign x_42943 = x_11655 & x_11656;
assign x_42944 = x_11657 & x_11658;
assign x_42945 = x_42943 & x_42944;
assign x_42946 = x_42942 & x_42945;
assign x_42947 = x_42939 & x_42946;
assign x_42948 = x_11659 & x_11660;
assign x_42949 = x_11661 & x_11662;
assign x_42950 = x_42948 & x_42949;
assign x_42951 = x_11663 & x_11664;
assign x_42952 = x_11665 & x_11666;
assign x_42953 = x_42951 & x_42952;
assign x_42954 = x_42950 & x_42953;
assign x_42955 = x_11667 & x_11668;
assign x_42956 = x_11669 & x_11670;
assign x_42957 = x_42955 & x_42956;
assign x_42958 = x_11671 & x_11672;
assign x_42959 = x_11673 & x_11674;
assign x_42960 = x_42958 & x_42959;
assign x_42961 = x_42957 & x_42960;
assign x_42962 = x_42954 & x_42961;
assign x_42963 = x_42947 & x_42962;
assign x_42964 = x_42933 & x_42963;
assign x_42965 = x_11676 & x_11677;
assign x_42966 = x_11675 & x_42965;
assign x_42967 = x_11678 & x_11679;
assign x_42968 = x_11680 & x_11681;
assign x_42969 = x_42967 & x_42968;
assign x_42970 = x_42966 & x_42969;
assign x_42971 = x_11682 & x_11683;
assign x_42972 = x_11684 & x_11685;
assign x_42973 = x_42971 & x_42972;
assign x_42974 = x_11686 & x_11687;
assign x_42975 = x_11688 & x_11689;
assign x_42976 = x_42974 & x_42975;
assign x_42977 = x_42973 & x_42976;
assign x_42978 = x_42970 & x_42977;
assign x_42979 = x_11690 & x_11691;
assign x_42980 = x_11692 & x_11693;
assign x_42981 = x_42979 & x_42980;
assign x_42982 = x_11694 & x_11695;
assign x_42983 = x_11696 & x_11697;
assign x_42984 = x_42982 & x_42983;
assign x_42985 = x_42981 & x_42984;
assign x_42986 = x_11698 & x_11699;
assign x_42987 = x_11700 & x_11701;
assign x_42988 = x_42986 & x_42987;
assign x_42989 = x_11702 & x_11703;
assign x_42990 = x_11704 & x_11705;
assign x_42991 = x_42989 & x_42990;
assign x_42992 = x_42988 & x_42991;
assign x_42993 = x_42985 & x_42992;
assign x_42994 = x_42978 & x_42993;
assign x_42995 = x_11707 & x_11708;
assign x_42996 = x_11706 & x_42995;
assign x_42997 = x_11709 & x_11710;
assign x_42998 = x_11711 & x_11712;
assign x_42999 = x_42997 & x_42998;
assign x_43000 = x_42996 & x_42999;
assign x_43001 = x_11713 & x_11714;
assign x_43002 = x_11715 & x_11716;
assign x_43003 = x_43001 & x_43002;
assign x_43004 = x_11717 & x_11718;
assign x_43005 = x_11719 & x_11720;
assign x_43006 = x_43004 & x_43005;
assign x_43007 = x_43003 & x_43006;
assign x_43008 = x_43000 & x_43007;
assign x_43009 = x_11721 & x_11722;
assign x_43010 = x_11723 & x_11724;
assign x_43011 = x_43009 & x_43010;
assign x_43012 = x_11725 & x_11726;
assign x_43013 = x_11727 & x_11728;
assign x_43014 = x_43012 & x_43013;
assign x_43015 = x_43011 & x_43014;
assign x_43016 = x_11729 & x_11730;
assign x_43017 = x_11731 & x_11732;
assign x_43018 = x_43016 & x_43017;
assign x_43019 = x_11733 & x_11734;
assign x_43020 = x_11735 & x_11736;
assign x_43021 = x_43019 & x_43020;
assign x_43022 = x_43018 & x_43021;
assign x_43023 = x_43015 & x_43022;
assign x_43024 = x_43008 & x_43023;
assign x_43025 = x_42994 & x_43024;
assign x_43026 = x_42964 & x_43025;
assign x_43027 = x_42904 & x_43026;
assign x_43028 = x_42783 & x_43027;
assign x_43029 = x_42540 & x_43028;
assign x_43030 = x_42052 & x_43029;
assign x_43031 = x_41075 & x_43030;
assign x_43032 = x_11738 & x_11739;
assign x_43033 = x_11737 & x_43032;
assign x_43034 = x_11740 & x_11741;
assign x_43035 = x_11742 & x_11743;
assign x_43036 = x_43034 & x_43035;
assign x_43037 = x_43033 & x_43036;
assign x_43038 = x_11744 & x_11745;
assign x_43039 = x_11746 & x_11747;
assign x_43040 = x_43038 & x_43039;
assign x_43041 = x_11748 & x_11749;
assign x_43042 = x_11750 & x_11751;
assign x_43043 = x_43041 & x_43042;
assign x_43044 = x_43040 & x_43043;
assign x_43045 = x_43037 & x_43044;
assign x_43046 = x_11753 & x_11754;
assign x_43047 = x_11752 & x_43046;
assign x_43048 = x_11755 & x_11756;
assign x_43049 = x_11757 & x_11758;
assign x_43050 = x_43048 & x_43049;
assign x_43051 = x_43047 & x_43050;
assign x_43052 = x_11759 & x_11760;
assign x_43053 = x_11761 & x_11762;
assign x_43054 = x_43052 & x_43053;
assign x_43055 = x_11763 & x_11764;
assign x_43056 = x_11765 & x_11766;
assign x_43057 = x_43055 & x_43056;
assign x_43058 = x_43054 & x_43057;
assign x_43059 = x_43051 & x_43058;
assign x_43060 = x_43045 & x_43059;
assign x_43061 = x_11768 & x_11769;
assign x_43062 = x_11767 & x_43061;
assign x_43063 = x_11770 & x_11771;
assign x_43064 = x_11772 & x_11773;
assign x_43065 = x_43063 & x_43064;
assign x_43066 = x_43062 & x_43065;
assign x_43067 = x_11774 & x_11775;
assign x_43068 = x_11776 & x_11777;
assign x_43069 = x_43067 & x_43068;
assign x_43070 = x_11778 & x_11779;
assign x_43071 = x_11780 & x_11781;
assign x_43072 = x_43070 & x_43071;
assign x_43073 = x_43069 & x_43072;
assign x_43074 = x_43066 & x_43073;
assign x_43075 = x_11782 & x_11783;
assign x_43076 = x_11784 & x_11785;
assign x_43077 = x_43075 & x_43076;
assign x_43078 = x_11786 & x_11787;
assign x_43079 = x_11788 & x_11789;
assign x_43080 = x_43078 & x_43079;
assign x_43081 = x_43077 & x_43080;
assign x_43082 = x_11790 & x_11791;
assign x_43083 = x_11792 & x_11793;
assign x_43084 = x_43082 & x_43083;
assign x_43085 = x_11794 & x_11795;
assign x_43086 = x_11796 & x_11797;
assign x_43087 = x_43085 & x_43086;
assign x_43088 = x_43084 & x_43087;
assign x_43089 = x_43081 & x_43088;
assign x_43090 = x_43074 & x_43089;
assign x_43091 = x_43060 & x_43090;
assign x_43092 = x_11799 & x_11800;
assign x_43093 = x_11798 & x_43092;
assign x_43094 = x_11801 & x_11802;
assign x_43095 = x_11803 & x_11804;
assign x_43096 = x_43094 & x_43095;
assign x_43097 = x_43093 & x_43096;
assign x_43098 = x_11805 & x_11806;
assign x_43099 = x_11807 & x_11808;
assign x_43100 = x_43098 & x_43099;
assign x_43101 = x_11809 & x_11810;
assign x_43102 = x_11811 & x_11812;
assign x_43103 = x_43101 & x_43102;
assign x_43104 = x_43100 & x_43103;
assign x_43105 = x_43097 & x_43104;
assign x_43106 = x_11814 & x_11815;
assign x_43107 = x_11813 & x_43106;
assign x_43108 = x_11816 & x_11817;
assign x_43109 = x_11818 & x_11819;
assign x_43110 = x_43108 & x_43109;
assign x_43111 = x_43107 & x_43110;
assign x_43112 = x_11820 & x_11821;
assign x_43113 = x_11822 & x_11823;
assign x_43114 = x_43112 & x_43113;
assign x_43115 = x_11824 & x_11825;
assign x_43116 = x_11826 & x_11827;
assign x_43117 = x_43115 & x_43116;
assign x_43118 = x_43114 & x_43117;
assign x_43119 = x_43111 & x_43118;
assign x_43120 = x_43105 & x_43119;
assign x_43121 = x_11829 & x_11830;
assign x_43122 = x_11828 & x_43121;
assign x_43123 = x_11831 & x_11832;
assign x_43124 = x_11833 & x_11834;
assign x_43125 = x_43123 & x_43124;
assign x_43126 = x_43122 & x_43125;
assign x_43127 = x_11835 & x_11836;
assign x_43128 = x_11837 & x_11838;
assign x_43129 = x_43127 & x_43128;
assign x_43130 = x_11839 & x_11840;
assign x_43131 = x_11841 & x_11842;
assign x_43132 = x_43130 & x_43131;
assign x_43133 = x_43129 & x_43132;
assign x_43134 = x_43126 & x_43133;
assign x_43135 = x_11843 & x_11844;
assign x_43136 = x_11845 & x_11846;
assign x_43137 = x_43135 & x_43136;
assign x_43138 = x_11847 & x_11848;
assign x_43139 = x_11849 & x_11850;
assign x_43140 = x_43138 & x_43139;
assign x_43141 = x_43137 & x_43140;
assign x_43142 = x_11851 & x_11852;
assign x_43143 = x_11853 & x_11854;
assign x_43144 = x_43142 & x_43143;
assign x_43145 = x_11855 & x_11856;
assign x_43146 = x_11857 & x_11858;
assign x_43147 = x_43145 & x_43146;
assign x_43148 = x_43144 & x_43147;
assign x_43149 = x_43141 & x_43148;
assign x_43150 = x_43134 & x_43149;
assign x_43151 = x_43120 & x_43150;
assign x_43152 = x_43091 & x_43151;
assign x_43153 = x_11860 & x_11861;
assign x_43154 = x_11859 & x_43153;
assign x_43155 = x_11862 & x_11863;
assign x_43156 = x_11864 & x_11865;
assign x_43157 = x_43155 & x_43156;
assign x_43158 = x_43154 & x_43157;
assign x_43159 = x_11866 & x_11867;
assign x_43160 = x_11868 & x_11869;
assign x_43161 = x_43159 & x_43160;
assign x_43162 = x_11870 & x_11871;
assign x_43163 = x_11872 & x_11873;
assign x_43164 = x_43162 & x_43163;
assign x_43165 = x_43161 & x_43164;
assign x_43166 = x_43158 & x_43165;
assign x_43167 = x_11875 & x_11876;
assign x_43168 = x_11874 & x_43167;
assign x_43169 = x_11877 & x_11878;
assign x_43170 = x_11879 & x_11880;
assign x_43171 = x_43169 & x_43170;
assign x_43172 = x_43168 & x_43171;
assign x_43173 = x_11881 & x_11882;
assign x_43174 = x_11883 & x_11884;
assign x_43175 = x_43173 & x_43174;
assign x_43176 = x_11885 & x_11886;
assign x_43177 = x_11887 & x_11888;
assign x_43178 = x_43176 & x_43177;
assign x_43179 = x_43175 & x_43178;
assign x_43180 = x_43172 & x_43179;
assign x_43181 = x_43166 & x_43180;
assign x_43182 = x_11890 & x_11891;
assign x_43183 = x_11889 & x_43182;
assign x_43184 = x_11892 & x_11893;
assign x_43185 = x_11894 & x_11895;
assign x_43186 = x_43184 & x_43185;
assign x_43187 = x_43183 & x_43186;
assign x_43188 = x_11896 & x_11897;
assign x_43189 = x_11898 & x_11899;
assign x_43190 = x_43188 & x_43189;
assign x_43191 = x_11900 & x_11901;
assign x_43192 = x_11902 & x_11903;
assign x_43193 = x_43191 & x_43192;
assign x_43194 = x_43190 & x_43193;
assign x_43195 = x_43187 & x_43194;
assign x_43196 = x_11904 & x_11905;
assign x_43197 = x_11906 & x_11907;
assign x_43198 = x_43196 & x_43197;
assign x_43199 = x_11908 & x_11909;
assign x_43200 = x_11910 & x_11911;
assign x_43201 = x_43199 & x_43200;
assign x_43202 = x_43198 & x_43201;
assign x_43203 = x_11912 & x_11913;
assign x_43204 = x_11914 & x_11915;
assign x_43205 = x_43203 & x_43204;
assign x_43206 = x_11916 & x_11917;
assign x_43207 = x_11918 & x_11919;
assign x_43208 = x_43206 & x_43207;
assign x_43209 = x_43205 & x_43208;
assign x_43210 = x_43202 & x_43209;
assign x_43211 = x_43195 & x_43210;
assign x_43212 = x_43181 & x_43211;
assign x_43213 = x_11921 & x_11922;
assign x_43214 = x_11920 & x_43213;
assign x_43215 = x_11923 & x_11924;
assign x_43216 = x_11925 & x_11926;
assign x_43217 = x_43215 & x_43216;
assign x_43218 = x_43214 & x_43217;
assign x_43219 = x_11927 & x_11928;
assign x_43220 = x_11929 & x_11930;
assign x_43221 = x_43219 & x_43220;
assign x_43222 = x_11931 & x_11932;
assign x_43223 = x_11933 & x_11934;
assign x_43224 = x_43222 & x_43223;
assign x_43225 = x_43221 & x_43224;
assign x_43226 = x_43218 & x_43225;
assign x_43227 = x_11936 & x_11937;
assign x_43228 = x_11935 & x_43227;
assign x_43229 = x_11938 & x_11939;
assign x_43230 = x_11940 & x_11941;
assign x_43231 = x_43229 & x_43230;
assign x_43232 = x_43228 & x_43231;
assign x_43233 = x_11942 & x_11943;
assign x_43234 = x_11944 & x_11945;
assign x_43235 = x_43233 & x_43234;
assign x_43236 = x_11946 & x_11947;
assign x_43237 = x_11948 & x_11949;
assign x_43238 = x_43236 & x_43237;
assign x_43239 = x_43235 & x_43238;
assign x_43240 = x_43232 & x_43239;
assign x_43241 = x_43226 & x_43240;
assign x_43242 = x_11951 & x_11952;
assign x_43243 = x_11950 & x_43242;
assign x_43244 = x_11953 & x_11954;
assign x_43245 = x_11955 & x_11956;
assign x_43246 = x_43244 & x_43245;
assign x_43247 = x_43243 & x_43246;
assign x_43248 = x_11957 & x_11958;
assign x_43249 = x_11959 & x_11960;
assign x_43250 = x_43248 & x_43249;
assign x_43251 = x_11961 & x_11962;
assign x_43252 = x_11963 & x_11964;
assign x_43253 = x_43251 & x_43252;
assign x_43254 = x_43250 & x_43253;
assign x_43255 = x_43247 & x_43254;
assign x_43256 = x_11965 & x_11966;
assign x_43257 = x_11967 & x_11968;
assign x_43258 = x_43256 & x_43257;
assign x_43259 = x_11969 & x_11970;
assign x_43260 = x_11971 & x_11972;
assign x_43261 = x_43259 & x_43260;
assign x_43262 = x_43258 & x_43261;
assign x_43263 = x_11973 & x_11974;
assign x_43264 = x_11975 & x_11976;
assign x_43265 = x_43263 & x_43264;
assign x_43266 = x_11977 & x_11978;
assign x_43267 = x_11979 & x_11980;
assign x_43268 = x_43266 & x_43267;
assign x_43269 = x_43265 & x_43268;
assign x_43270 = x_43262 & x_43269;
assign x_43271 = x_43255 & x_43270;
assign x_43272 = x_43241 & x_43271;
assign x_43273 = x_43212 & x_43272;
assign x_43274 = x_43152 & x_43273;
assign x_43275 = x_11982 & x_11983;
assign x_43276 = x_11981 & x_43275;
assign x_43277 = x_11984 & x_11985;
assign x_43278 = x_11986 & x_11987;
assign x_43279 = x_43277 & x_43278;
assign x_43280 = x_43276 & x_43279;
assign x_43281 = x_11988 & x_11989;
assign x_43282 = x_11990 & x_11991;
assign x_43283 = x_43281 & x_43282;
assign x_43284 = x_11992 & x_11993;
assign x_43285 = x_11994 & x_11995;
assign x_43286 = x_43284 & x_43285;
assign x_43287 = x_43283 & x_43286;
assign x_43288 = x_43280 & x_43287;
assign x_43289 = x_11997 & x_11998;
assign x_43290 = x_11996 & x_43289;
assign x_43291 = x_11999 & x_12000;
assign x_43292 = x_12001 & x_12002;
assign x_43293 = x_43291 & x_43292;
assign x_43294 = x_43290 & x_43293;
assign x_43295 = x_12003 & x_12004;
assign x_43296 = x_12005 & x_12006;
assign x_43297 = x_43295 & x_43296;
assign x_43298 = x_12007 & x_12008;
assign x_43299 = x_12009 & x_12010;
assign x_43300 = x_43298 & x_43299;
assign x_43301 = x_43297 & x_43300;
assign x_43302 = x_43294 & x_43301;
assign x_43303 = x_43288 & x_43302;
assign x_43304 = x_12012 & x_12013;
assign x_43305 = x_12011 & x_43304;
assign x_43306 = x_12014 & x_12015;
assign x_43307 = x_12016 & x_12017;
assign x_43308 = x_43306 & x_43307;
assign x_43309 = x_43305 & x_43308;
assign x_43310 = x_12018 & x_12019;
assign x_43311 = x_12020 & x_12021;
assign x_43312 = x_43310 & x_43311;
assign x_43313 = x_12022 & x_12023;
assign x_43314 = x_12024 & x_12025;
assign x_43315 = x_43313 & x_43314;
assign x_43316 = x_43312 & x_43315;
assign x_43317 = x_43309 & x_43316;
assign x_43318 = x_12026 & x_12027;
assign x_43319 = x_12028 & x_12029;
assign x_43320 = x_43318 & x_43319;
assign x_43321 = x_12030 & x_12031;
assign x_43322 = x_12032 & x_12033;
assign x_43323 = x_43321 & x_43322;
assign x_43324 = x_43320 & x_43323;
assign x_43325 = x_12034 & x_12035;
assign x_43326 = x_12036 & x_12037;
assign x_43327 = x_43325 & x_43326;
assign x_43328 = x_12038 & x_12039;
assign x_43329 = x_12040 & x_12041;
assign x_43330 = x_43328 & x_43329;
assign x_43331 = x_43327 & x_43330;
assign x_43332 = x_43324 & x_43331;
assign x_43333 = x_43317 & x_43332;
assign x_43334 = x_43303 & x_43333;
assign x_43335 = x_12043 & x_12044;
assign x_43336 = x_12042 & x_43335;
assign x_43337 = x_12045 & x_12046;
assign x_43338 = x_12047 & x_12048;
assign x_43339 = x_43337 & x_43338;
assign x_43340 = x_43336 & x_43339;
assign x_43341 = x_12049 & x_12050;
assign x_43342 = x_12051 & x_12052;
assign x_43343 = x_43341 & x_43342;
assign x_43344 = x_12053 & x_12054;
assign x_43345 = x_12055 & x_12056;
assign x_43346 = x_43344 & x_43345;
assign x_43347 = x_43343 & x_43346;
assign x_43348 = x_43340 & x_43347;
assign x_43349 = x_12058 & x_12059;
assign x_43350 = x_12057 & x_43349;
assign x_43351 = x_12060 & x_12061;
assign x_43352 = x_12062 & x_12063;
assign x_43353 = x_43351 & x_43352;
assign x_43354 = x_43350 & x_43353;
assign x_43355 = x_12064 & x_12065;
assign x_43356 = x_12066 & x_12067;
assign x_43357 = x_43355 & x_43356;
assign x_43358 = x_12068 & x_12069;
assign x_43359 = x_12070 & x_12071;
assign x_43360 = x_43358 & x_43359;
assign x_43361 = x_43357 & x_43360;
assign x_43362 = x_43354 & x_43361;
assign x_43363 = x_43348 & x_43362;
assign x_43364 = x_12073 & x_12074;
assign x_43365 = x_12072 & x_43364;
assign x_43366 = x_12075 & x_12076;
assign x_43367 = x_12077 & x_12078;
assign x_43368 = x_43366 & x_43367;
assign x_43369 = x_43365 & x_43368;
assign x_43370 = x_12079 & x_12080;
assign x_43371 = x_12081 & x_12082;
assign x_43372 = x_43370 & x_43371;
assign x_43373 = x_12083 & x_12084;
assign x_43374 = x_12085 & x_12086;
assign x_43375 = x_43373 & x_43374;
assign x_43376 = x_43372 & x_43375;
assign x_43377 = x_43369 & x_43376;
assign x_43378 = x_12087 & x_12088;
assign x_43379 = x_12089 & x_12090;
assign x_43380 = x_43378 & x_43379;
assign x_43381 = x_12091 & x_12092;
assign x_43382 = x_12093 & x_12094;
assign x_43383 = x_43381 & x_43382;
assign x_43384 = x_43380 & x_43383;
assign x_43385 = x_12095 & x_12096;
assign x_43386 = x_12097 & x_12098;
assign x_43387 = x_43385 & x_43386;
assign x_43388 = x_12099 & x_12100;
assign x_43389 = x_12101 & x_12102;
assign x_43390 = x_43388 & x_43389;
assign x_43391 = x_43387 & x_43390;
assign x_43392 = x_43384 & x_43391;
assign x_43393 = x_43377 & x_43392;
assign x_43394 = x_43363 & x_43393;
assign x_43395 = x_43334 & x_43394;
assign x_43396 = x_12104 & x_12105;
assign x_43397 = x_12103 & x_43396;
assign x_43398 = x_12106 & x_12107;
assign x_43399 = x_12108 & x_12109;
assign x_43400 = x_43398 & x_43399;
assign x_43401 = x_43397 & x_43400;
assign x_43402 = x_12110 & x_12111;
assign x_43403 = x_12112 & x_12113;
assign x_43404 = x_43402 & x_43403;
assign x_43405 = x_12114 & x_12115;
assign x_43406 = x_12116 & x_12117;
assign x_43407 = x_43405 & x_43406;
assign x_43408 = x_43404 & x_43407;
assign x_43409 = x_43401 & x_43408;
assign x_43410 = x_12119 & x_12120;
assign x_43411 = x_12118 & x_43410;
assign x_43412 = x_12121 & x_12122;
assign x_43413 = x_12123 & x_12124;
assign x_43414 = x_43412 & x_43413;
assign x_43415 = x_43411 & x_43414;
assign x_43416 = x_12125 & x_12126;
assign x_43417 = x_12127 & x_12128;
assign x_43418 = x_43416 & x_43417;
assign x_43419 = x_12129 & x_12130;
assign x_43420 = x_12131 & x_12132;
assign x_43421 = x_43419 & x_43420;
assign x_43422 = x_43418 & x_43421;
assign x_43423 = x_43415 & x_43422;
assign x_43424 = x_43409 & x_43423;
assign x_43425 = x_12134 & x_12135;
assign x_43426 = x_12133 & x_43425;
assign x_43427 = x_12136 & x_12137;
assign x_43428 = x_12138 & x_12139;
assign x_43429 = x_43427 & x_43428;
assign x_43430 = x_43426 & x_43429;
assign x_43431 = x_12140 & x_12141;
assign x_43432 = x_12142 & x_12143;
assign x_43433 = x_43431 & x_43432;
assign x_43434 = x_12144 & x_12145;
assign x_43435 = x_12146 & x_12147;
assign x_43436 = x_43434 & x_43435;
assign x_43437 = x_43433 & x_43436;
assign x_43438 = x_43430 & x_43437;
assign x_43439 = x_12148 & x_12149;
assign x_43440 = x_12150 & x_12151;
assign x_43441 = x_43439 & x_43440;
assign x_43442 = x_12152 & x_12153;
assign x_43443 = x_12154 & x_12155;
assign x_43444 = x_43442 & x_43443;
assign x_43445 = x_43441 & x_43444;
assign x_43446 = x_12156 & x_12157;
assign x_43447 = x_12158 & x_12159;
assign x_43448 = x_43446 & x_43447;
assign x_43449 = x_12160 & x_12161;
assign x_43450 = x_12162 & x_12163;
assign x_43451 = x_43449 & x_43450;
assign x_43452 = x_43448 & x_43451;
assign x_43453 = x_43445 & x_43452;
assign x_43454 = x_43438 & x_43453;
assign x_43455 = x_43424 & x_43454;
assign x_43456 = x_12165 & x_12166;
assign x_43457 = x_12164 & x_43456;
assign x_43458 = x_12167 & x_12168;
assign x_43459 = x_12169 & x_12170;
assign x_43460 = x_43458 & x_43459;
assign x_43461 = x_43457 & x_43460;
assign x_43462 = x_12171 & x_12172;
assign x_43463 = x_12173 & x_12174;
assign x_43464 = x_43462 & x_43463;
assign x_43465 = x_12175 & x_12176;
assign x_43466 = x_12177 & x_12178;
assign x_43467 = x_43465 & x_43466;
assign x_43468 = x_43464 & x_43467;
assign x_43469 = x_43461 & x_43468;
assign x_43470 = x_12179 & x_12180;
assign x_43471 = x_12181 & x_12182;
assign x_43472 = x_43470 & x_43471;
assign x_43473 = x_12183 & x_12184;
assign x_43474 = x_12185 & x_12186;
assign x_43475 = x_43473 & x_43474;
assign x_43476 = x_43472 & x_43475;
assign x_43477 = x_12187 & x_12188;
assign x_43478 = x_12189 & x_12190;
assign x_43479 = x_43477 & x_43478;
assign x_43480 = x_12191 & x_12192;
assign x_43481 = x_12193 & x_12194;
assign x_43482 = x_43480 & x_43481;
assign x_43483 = x_43479 & x_43482;
assign x_43484 = x_43476 & x_43483;
assign x_43485 = x_43469 & x_43484;
assign x_43486 = x_12196 & x_12197;
assign x_43487 = x_12195 & x_43486;
assign x_43488 = x_12198 & x_12199;
assign x_43489 = x_12200 & x_12201;
assign x_43490 = x_43488 & x_43489;
assign x_43491 = x_43487 & x_43490;
assign x_43492 = x_12202 & x_12203;
assign x_43493 = x_12204 & x_12205;
assign x_43494 = x_43492 & x_43493;
assign x_43495 = x_12206 & x_12207;
assign x_43496 = x_12208 & x_12209;
assign x_43497 = x_43495 & x_43496;
assign x_43498 = x_43494 & x_43497;
assign x_43499 = x_43491 & x_43498;
assign x_43500 = x_12210 & x_12211;
assign x_43501 = x_12212 & x_12213;
assign x_43502 = x_43500 & x_43501;
assign x_43503 = x_12214 & x_12215;
assign x_43504 = x_12216 & x_12217;
assign x_43505 = x_43503 & x_43504;
assign x_43506 = x_43502 & x_43505;
assign x_43507 = x_12218 & x_12219;
assign x_43508 = x_12220 & x_12221;
assign x_43509 = x_43507 & x_43508;
assign x_43510 = x_12222 & x_12223;
assign x_43511 = x_12224 & x_12225;
assign x_43512 = x_43510 & x_43511;
assign x_43513 = x_43509 & x_43512;
assign x_43514 = x_43506 & x_43513;
assign x_43515 = x_43499 & x_43514;
assign x_43516 = x_43485 & x_43515;
assign x_43517 = x_43455 & x_43516;
assign x_43518 = x_43395 & x_43517;
assign x_43519 = x_43274 & x_43518;
assign x_43520 = x_12227 & x_12228;
assign x_43521 = x_12226 & x_43520;
assign x_43522 = x_12229 & x_12230;
assign x_43523 = x_12231 & x_12232;
assign x_43524 = x_43522 & x_43523;
assign x_43525 = x_43521 & x_43524;
assign x_43526 = x_12233 & x_12234;
assign x_43527 = x_12235 & x_12236;
assign x_43528 = x_43526 & x_43527;
assign x_43529 = x_12237 & x_12238;
assign x_43530 = x_12239 & x_12240;
assign x_43531 = x_43529 & x_43530;
assign x_43532 = x_43528 & x_43531;
assign x_43533 = x_43525 & x_43532;
assign x_43534 = x_12242 & x_12243;
assign x_43535 = x_12241 & x_43534;
assign x_43536 = x_12244 & x_12245;
assign x_43537 = x_12246 & x_12247;
assign x_43538 = x_43536 & x_43537;
assign x_43539 = x_43535 & x_43538;
assign x_43540 = x_12248 & x_12249;
assign x_43541 = x_12250 & x_12251;
assign x_43542 = x_43540 & x_43541;
assign x_43543 = x_12252 & x_12253;
assign x_43544 = x_12254 & x_12255;
assign x_43545 = x_43543 & x_43544;
assign x_43546 = x_43542 & x_43545;
assign x_43547 = x_43539 & x_43546;
assign x_43548 = x_43533 & x_43547;
assign x_43549 = x_12257 & x_12258;
assign x_43550 = x_12256 & x_43549;
assign x_43551 = x_12259 & x_12260;
assign x_43552 = x_12261 & x_12262;
assign x_43553 = x_43551 & x_43552;
assign x_43554 = x_43550 & x_43553;
assign x_43555 = x_12263 & x_12264;
assign x_43556 = x_12265 & x_12266;
assign x_43557 = x_43555 & x_43556;
assign x_43558 = x_12267 & x_12268;
assign x_43559 = x_12269 & x_12270;
assign x_43560 = x_43558 & x_43559;
assign x_43561 = x_43557 & x_43560;
assign x_43562 = x_43554 & x_43561;
assign x_43563 = x_12271 & x_12272;
assign x_43564 = x_12273 & x_12274;
assign x_43565 = x_43563 & x_43564;
assign x_43566 = x_12275 & x_12276;
assign x_43567 = x_12277 & x_12278;
assign x_43568 = x_43566 & x_43567;
assign x_43569 = x_43565 & x_43568;
assign x_43570 = x_12279 & x_12280;
assign x_43571 = x_12281 & x_12282;
assign x_43572 = x_43570 & x_43571;
assign x_43573 = x_12283 & x_12284;
assign x_43574 = x_12285 & x_12286;
assign x_43575 = x_43573 & x_43574;
assign x_43576 = x_43572 & x_43575;
assign x_43577 = x_43569 & x_43576;
assign x_43578 = x_43562 & x_43577;
assign x_43579 = x_43548 & x_43578;
assign x_43580 = x_12288 & x_12289;
assign x_43581 = x_12287 & x_43580;
assign x_43582 = x_12290 & x_12291;
assign x_43583 = x_12292 & x_12293;
assign x_43584 = x_43582 & x_43583;
assign x_43585 = x_43581 & x_43584;
assign x_43586 = x_12294 & x_12295;
assign x_43587 = x_12296 & x_12297;
assign x_43588 = x_43586 & x_43587;
assign x_43589 = x_12298 & x_12299;
assign x_43590 = x_12300 & x_12301;
assign x_43591 = x_43589 & x_43590;
assign x_43592 = x_43588 & x_43591;
assign x_43593 = x_43585 & x_43592;
assign x_43594 = x_12303 & x_12304;
assign x_43595 = x_12302 & x_43594;
assign x_43596 = x_12305 & x_12306;
assign x_43597 = x_12307 & x_12308;
assign x_43598 = x_43596 & x_43597;
assign x_43599 = x_43595 & x_43598;
assign x_43600 = x_12309 & x_12310;
assign x_43601 = x_12311 & x_12312;
assign x_43602 = x_43600 & x_43601;
assign x_43603 = x_12313 & x_12314;
assign x_43604 = x_12315 & x_12316;
assign x_43605 = x_43603 & x_43604;
assign x_43606 = x_43602 & x_43605;
assign x_43607 = x_43599 & x_43606;
assign x_43608 = x_43593 & x_43607;
assign x_43609 = x_12318 & x_12319;
assign x_43610 = x_12317 & x_43609;
assign x_43611 = x_12320 & x_12321;
assign x_43612 = x_12322 & x_12323;
assign x_43613 = x_43611 & x_43612;
assign x_43614 = x_43610 & x_43613;
assign x_43615 = x_12324 & x_12325;
assign x_43616 = x_12326 & x_12327;
assign x_43617 = x_43615 & x_43616;
assign x_43618 = x_12328 & x_12329;
assign x_43619 = x_12330 & x_12331;
assign x_43620 = x_43618 & x_43619;
assign x_43621 = x_43617 & x_43620;
assign x_43622 = x_43614 & x_43621;
assign x_43623 = x_12332 & x_12333;
assign x_43624 = x_12334 & x_12335;
assign x_43625 = x_43623 & x_43624;
assign x_43626 = x_12336 & x_12337;
assign x_43627 = x_12338 & x_12339;
assign x_43628 = x_43626 & x_43627;
assign x_43629 = x_43625 & x_43628;
assign x_43630 = x_12340 & x_12341;
assign x_43631 = x_12342 & x_12343;
assign x_43632 = x_43630 & x_43631;
assign x_43633 = x_12344 & x_12345;
assign x_43634 = x_12346 & x_12347;
assign x_43635 = x_43633 & x_43634;
assign x_43636 = x_43632 & x_43635;
assign x_43637 = x_43629 & x_43636;
assign x_43638 = x_43622 & x_43637;
assign x_43639 = x_43608 & x_43638;
assign x_43640 = x_43579 & x_43639;
assign x_43641 = x_12349 & x_12350;
assign x_43642 = x_12348 & x_43641;
assign x_43643 = x_12351 & x_12352;
assign x_43644 = x_12353 & x_12354;
assign x_43645 = x_43643 & x_43644;
assign x_43646 = x_43642 & x_43645;
assign x_43647 = x_12355 & x_12356;
assign x_43648 = x_12357 & x_12358;
assign x_43649 = x_43647 & x_43648;
assign x_43650 = x_12359 & x_12360;
assign x_43651 = x_12361 & x_12362;
assign x_43652 = x_43650 & x_43651;
assign x_43653 = x_43649 & x_43652;
assign x_43654 = x_43646 & x_43653;
assign x_43655 = x_12364 & x_12365;
assign x_43656 = x_12363 & x_43655;
assign x_43657 = x_12366 & x_12367;
assign x_43658 = x_12368 & x_12369;
assign x_43659 = x_43657 & x_43658;
assign x_43660 = x_43656 & x_43659;
assign x_43661 = x_12370 & x_12371;
assign x_43662 = x_12372 & x_12373;
assign x_43663 = x_43661 & x_43662;
assign x_43664 = x_12374 & x_12375;
assign x_43665 = x_12376 & x_12377;
assign x_43666 = x_43664 & x_43665;
assign x_43667 = x_43663 & x_43666;
assign x_43668 = x_43660 & x_43667;
assign x_43669 = x_43654 & x_43668;
assign x_43670 = x_12379 & x_12380;
assign x_43671 = x_12378 & x_43670;
assign x_43672 = x_12381 & x_12382;
assign x_43673 = x_12383 & x_12384;
assign x_43674 = x_43672 & x_43673;
assign x_43675 = x_43671 & x_43674;
assign x_43676 = x_12385 & x_12386;
assign x_43677 = x_12387 & x_12388;
assign x_43678 = x_43676 & x_43677;
assign x_43679 = x_12389 & x_12390;
assign x_43680 = x_12391 & x_12392;
assign x_43681 = x_43679 & x_43680;
assign x_43682 = x_43678 & x_43681;
assign x_43683 = x_43675 & x_43682;
assign x_43684 = x_12393 & x_12394;
assign x_43685 = x_12395 & x_12396;
assign x_43686 = x_43684 & x_43685;
assign x_43687 = x_12397 & x_12398;
assign x_43688 = x_12399 & x_12400;
assign x_43689 = x_43687 & x_43688;
assign x_43690 = x_43686 & x_43689;
assign x_43691 = x_12401 & x_12402;
assign x_43692 = x_12403 & x_12404;
assign x_43693 = x_43691 & x_43692;
assign x_43694 = x_12405 & x_12406;
assign x_43695 = x_12407 & x_12408;
assign x_43696 = x_43694 & x_43695;
assign x_43697 = x_43693 & x_43696;
assign x_43698 = x_43690 & x_43697;
assign x_43699 = x_43683 & x_43698;
assign x_43700 = x_43669 & x_43699;
assign x_43701 = x_12410 & x_12411;
assign x_43702 = x_12409 & x_43701;
assign x_43703 = x_12412 & x_12413;
assign x_43704 = x_12414 & x_12415;
assign x_43705 = x_43703 & x_43704;
assign x_43706 = x_43702 & x_43705;
assign x_43707 = x_12416 & x_12417;
assign x_43708 = x_12418 & x_12419;
assign x_43709 = x_43707 & x_43708;
assign x_43710 = x_12420 & x_12421;
assign x_43711 = x_12422 & x_12423;
assign x_43712 = x_43710 & x_43711;
assign x_43713 = x_43709 & x_43712;
assign x_43714 = x_43706 & x_43713;
assign x_43715 = x_12425 & x_12426;
assign x_43716 = x_12424 & x_43715;
assign x_43717 = x_12427 & x_12428;
assign x_43718 = x_12429 & x_12430;
assign x_43719 = x_43717 & x_43718;
assign x_43720 = x_43716 & x_43719;
assign x_43721 = x_12431 & x_12432;
assign x_43722 = x_12433 & x_12434;
assign x_43723 = x_43721 & x_43722;
assign x_43724 = x_12435 & x_12436;
assign x_43725 = x_12437 & x_12438;
assign x_43726 = x_43724 & x_43725;
assign x_43727 = x_43723 & x_43726;
assign x_43728 = x_43720 & x_43727;
assign x_43729 = x_43714 & x_43728;
assign x_43730 = x_12440 & x_12441;
assign x_43731 = x_12439 & x_43730;
assign x_43732 = x_12442 & x_12443;
assign x_43733 = x_12444 & x_12445;
assign x_43734 = x_43732 & x_43733;
assign x_43735 = x_43731 & x_43734;
assign x_43736 = x_12446 & x_12447;
assign x_43737 = x_12448 & x_12449;
assign x_43738 = x_43736 & x_43737;
assign x_43739 = x_12450 & x_12451;
assign x_43740 = x_12452 & x_12453;
assign x_43741 = x_43739 & x_43740;
assign x_43742 = x_43738 & x_43741;
assign x_43743 = x_43735 & x_43742;
assign x_43744 = x_12454 & x_12455;
assign x_43745 = x_12456 & x_12457;
assign x_43746 = x_43744 & x_43745;
assign x_43747 = x_12458 & x_12459;
assign x_43748 = x_12460 & x_12461;
assign x_43749 = x_43747 & x_43748;
assign x_43750 = x_43746 & x_43749;
assign x_43751 = x_12462 & x_12463;
assign x_43752 = x_12464 & x_12465;
assign x_43753 = x_43751 & x_43752;
assign x_43754 = x_12466 & x_12467;
assign x_43755 = x_12468 & x_12469;
assign x_43756 = x_43754 & x_43755;
assign x_43757 = x_43753 & x_43756;
assign x_43758 = x_43750 & x_43757;
assign x_43759 = x_43743 & x_43758;
assign x_43760 = x_43729 & x_43759;
assign x_43761 = x_43700 & x_43760;
assign x_43762 = x_43640 & x_43761;
assign x_43763 = x_12471 & x_12472;
assign x_43764 = x_12470 & x_43763;
assign x_43765 = x_12473 & x_12474;
assign x_43766 = x_12475 & x_12476;
assign x_43767 = x_43765 & x_43766;
assign x_43768 = x_43764 & x_43767;
assign x_43769 = x_12477 & x_12478;
assign x_43770 = x_12479 & x_12480;
assign x_43771 = x_43769 & x_43770;
assign x_43772 = x_12481 & x_12482;
assign x_43773 = x_12483 & x_12484;
assign x_43774 = x_43772 & x_43773;
assign x_43775 = x_43771 & x_43774;
assign x_43776 = x_43768 & x_43775;
assign x_43777 = x_12486 & x_12487;
assign x_43778 = x_12485 & x_43777;
assign x_43779 = x_12488 & x_12489;
assign x_43780 = x_12490 & x_12491;
assign x_43781 = x_43779 & x_43780;
assign x_43782 = x_43778 & x_43781;
assign x_43783 = x_12492 & x_12493;
assign x_43784 = x_12494 & x_12495;
assign x_43785 = x_43783 & x_43784;
assign x_43786 = x_12496 & x_12497;
assign x_43787 = x_12498 & x_12499;
assign x_43788 = x_43786 & x_43787;
assign x_43789 = x_43785 & x_43788;
assign x_43790 = x_43782 & x_43789;
assign x_43791 = x_43776 & x_43790;
assign x_43792 = x_12501 & x_12502;
assign x_43793 = x_12500 & x_43792;
assign x_43794 = x_12503 & x_12504;
assign x_43795 = x_12505 & x_12506;
assign x_43796 = x_43794 & x_43795;
assign x_43797 = x_43793 & x_43796;
assign x_43798 = x_12507 & x_12508;
assign x_43799 = x_12509 & x_12510;
assign x_43800 = x_43798 & x_43799;
assign x_43801 = x_12511 & x_12512;
assign x_43802 = x_12513 & x_12514;
assign x_43803 = x_43801 & x_43802;
assign x_43804 = x_43800 & x_43803;
assign x_43805 = x_43797 & x_43804;
assign x_43806 = x_12515 & x_12516;
assign x_43807 = x_12517 & x_12518;
assign x_43808 = x_43806 & x_43807;
assign x_43809 = x_12519 & x_12520;
assign x_43810 = x_12521 & x_12522;
assign x_43811 = x_43809 & x_43810;
assign x_43812 = x_43808 & x_43811;
assign x_43813 = x_12523 & x_12524;
assign x_43814 = x_12525 & x_12526;
assign x_43815 = x_43813 & x_43814;
assign x_43816 = x_12527 & x_12528;
assign x_43817 = x_12529 & x_12530;
assign x_43818 = x_43816 & x_43817;
assign x_43819 = x_43815 & x_43818;
assign x_43820 = x_43812 & x_43819;
assign x_43821 = x_43805 & x_43820;
assign x_43822 = x_43791 & x_43821;
assign x_43823 = x_12532 & x_12533;
assign x_43824 = x_12531 & x_43823;
assign x_43825 = x_12534 & x_12535;
assign x_43826 = x_12536 & x_12537;
assign x_43827 = x_43825 & x_43826;
assign x_43828 = x_43824 & x_43827;
assign x_43829 = x_12538 & x_12539;
assign x_43830 = x_12540 & x_12541;
assign x_43831 = x_43829 & x_43830;
assign x_43832 = x_12542 & x_12543;
assign x_43833 = x_12544 & x_12545;
assign x_43834 = x_43832 & x_43833;
assign x_43835 = x_43831 & x_43834;
assign x_43836 = x_43828 & x_43835;
assign x_43837 = x_12547 & x_12548;
assign x_43838 = x_12546 & x_43837;
assign x_43839 = x_12549 & x_12550;
assign x_43840 = x_12551 & x_12552;
assign x_43841 = x_43839 & x_43840;
assign x_43842 = x_43838 & x_43841;
assign x_43843 = x_12553 & x_12554;
assign x_43844 = x_12555 & x_12556;
assign x_43845 = x_43843 & x_43844;
assign x_43846 = x_12557 & x_12558;
assign x_43847 = x_12559 & x_12560;
assign x_43848 = x_43846 & x_43847;
assign x_43849 = x_43845 & x_43848;
assign x_43850 = x_43842 & x_43849;
assign x_43851 = x_43836 & x_43850;
assign x_43852 = x_12562 & x_12563;
assign x_43853 = x_12561 & x_43852;
assign x_43854 = x_12564 & x_12565;
assign x_43855 = x_12566 & x_12567;
assign x_43856 = x_43854 & x_43855;
assign x_43857 = x_43853 & x_43856;
assign x_43858 = x_12568 & x_12569;
assign x_43859 = x_12570 & x_12571;
assign x_43860 = x_43858 & x_43859;
assign x_43861 = x_12572 & x_12573;
assign x_43862 = x_12574 & x_12575;
assign x_43863 = x_43861 & x_43862;
assign x_43864 = x_43860 & x_43863;
assign x_43865 = x_43857 & x_43864;
assign x_43866 = x_12576 & x_12577;
assign x_43867 = x_12578 & x_12579;
assign x_43868 = x_43866 & x_43867;
assign x_43869 = x_12580 & x_12581;
assign x_43870 = x_12582 & x_12583;
assign x_43871 = x_43869 & x_43870;
assign x_43872 = x_43868 & x_43871;
assign x_43873 = x_12584 & x_12585;
assign x_43874 = x_12586 & x_12587;
assign x_43875 = x_43873 & x_43874;
assign x_43876 = x_12588 & x_12589;
assign x_43877 = x_12590 & x_12591;
assign x_43878 = x_43876 & x_43877;
assign x_43879 = x_43875 & x_43878;
assign x_43880 = x_43872 & x_43879;
assign x_43881 = x_43865 & x_43880;
assign x_43882 = x_43851 & x_43881;
assign x_43883 = x_43822 & x_43882;
assign x_43884 = x_12593 & x_12594;
assign x_43885 = x_12592 & x_43884;
assign x_43886 = x_12595 & x_12596;
assign x_43887 = x_12597 & x_12598;
assign x_43888 = x_43886 & x_43887;
assign x_43889 = x_43885 & x_43888;
assign x_43890 = x_12599 & x_12600;
assign x_43891 = x_12601 & x_12602;
assign x_43892 = x_43890 & x_43891;
assign x_43893 = x_12603 & x_12604;
assign x_43894 = x_12605 & x_12606;
assign x_43895 = x_43893 & x_43894;
assign x_43896 = x_43892 & x_43895;
assign x_43897 = x_43889 & x_43896;
assign x_43898 = x_12608 & x_12609;
assign x_43899 = x_12607 & x_43898;
assign x_43900 = x_12610 & x_12611;
assign x_43901 = x_12612 & x_12613;
assign x_43902 = x_43900 & x_43901;
assign x_43903 = x_43899 & x_43902;
assign x_43904 = x_12614 & x_12615;
assign x_43905 = x_12616 & x_12617;
assign x_43906 = x_43904 & x_43905;
assign x_43907 = x_12618 & x_12619;
assign x_43908 = x_12620 & x_12621;
assign x_43909 = x_43907 & x_43908;
assign x_43910 = x_43906 & x_43909;
assign x_43911 = x_43903 & x_43910;
assign x_43912 = x_43897 & x_43911;
assign x_43913 = x_12623 & x_12624;
assign x_43914 = x_12622 & x_43913;
assign x_43915 = x_12625 & x_12626;
assign x_43916 = x_12627 & x_12628;
assign x_43917 = x_43915 & x_43916;
assign x_43918 = x_43914 & x_43917;
assign x_43919 = x_12629 & x_12630;
assign x_43920 = x_12631 & x_12632;
assign x_43921 = x_43919 & x_43920;
assign x_43922 = x_12633 & x_12634;
assign x_43923 = x_12635 & x_12636;
assign x_43924 = x_43922 & x_43923;
assign x_43925 = x_43921 & x_43924;
assign x_43926 = x_43918 & x_43925;
assign x_43927 = x_12637 & x_12638;
assign x_43928 = x_12639 & x_12640;
assign x_43929 = x_43927 & x_43928;
assign x_43930 = x_12641 & x_12642;
assign x_43931 = x_12643 & x_12644;
assign x_43932 = x_43930 & x_43931;
assign x_43933 = x_43929 & x_43932;
assign x_43934 = x_12645 & x_12646;
assign x_43935 = x_12647 & x_12648;
assign x_43936 = x_43934 & x_43935;
assign x_43937 = x_12649 & x_12650;
assign x_43938 = x_12651 & x_12652;
assign x_43939 = x_43937 & x_43938;
assign x_43940 = x_43936 & x_43939;
assign x_43941 = x_43933 & x_43940;
assign x_43942 = x_43926 & x_43941;
assign x_43943 = x_43912 & x_43942;
assign x_43944 = x_12654 & x_12655;
assign x_43945 = x_12653 & x_43944;
assign x_43946 = x_12656 & x_12657;
assign x_43947 = x_12658 & x_12659;
assign x_43948 = x_43946 & x_43947;
assign x_43949 = x_43945 & x_43948;
assign x_43950 = x_12660 & x_12661;
assign x_43951 = x_12662 & x_12663;
assign x_43952 = x_43950 & x_43951;
assign x_43953 = x_12664 & x_12665;
assign x_43954 = x_12666 & x_12667;
assign x_43955 = x_43953 & x_43954;
assign x_43956 = x_43952 & x_43955;
assign x_43957 = x_43949 & x_43956;
assign x_43958 = x_12668 & x_12669;
assign x_43959 = x_12670 & x_12671;
assign x_43960 = x_43958 & x_43959;
assign x_43961 = x_12672 & x_12673;
assign x_43962 = x_12674 & x_12675;
assign x_43963 = x_43961 & x_43962;
assign x_43964 = x_43960 & x_43963;
assign x_43965 = x_12676 & x_12677;
assign x_43966 = x_12678 & x_12679;
assign x_43967 = x_43965 & x_43966;
assign x_43968 = x_12680 & x_12681;
assign x_43969 = x_12682 & x_12683;
assign x_43970 = x_43968 & x_43969;
assign x_43971 = x_43967 & x_43970;
assign x_43972 = x_43964 & x_43971;
assign x_43973 = x_43957 & x_43972;
assign x_43974 = x_12685 & x_12686;
assign x_43975 = x_12684 & x_43974;
assign x_43976 = x_12687 & x_12688;
assign x_43977 = x_12689 & x_12690;
assign x_43978 = x_43976 & x_43977;
assign x_43979 = x_43975 & x_43978;
assign x_43980 = x_12691 & x_12692;
assign x_43981 = x_12693 & x_12694;
assign x_43982 = x_43980 & x_43981;
assign x_43983 = x_12695 & x_12696;
assign x_43984 = x_12697 & x_12698;
assign x_43985 = x_43983 & x_43984;
assign x_43986 = x_43982 & x_43985;
assign x_43987 = x_43979 & x_43986;
assign x_43988 = x_12699 & x_12700;
assign x_43989 = x_12701 & x_12702;
assign x_43990 = x_43988 & x_43989;
assign x_43991 = x_12703 & x_12704;
assign x_43992 = x_12705 & x_12706;
assign x_43993 = x_43991 & x_43992;
assign x_43994 = x_43990 & x_43993;
assign x_43995 = x_12707 & x_12708;
assign x_43996 = x_12709 & x_12710;
assign x_43997 = x_43995 & x_43996;
assign x_43998 = x_12711 & x_12712;
assign x_43999 = x_12713 & x_12714;
assign x_44000 = x_43998 & x_43999;
assign x_44001 = x_43997 & x_44000;
assign x_44002 = x_43994 & x_44001;
assign x_44003 = x_43987 & x_44002;
assign x_44004 = x_43973 & x_44003;
assign x_44005 = x_43943 & x_44004;
assign x_44006 = x_43883 & x_44005;
assign x_44007 = x_43762 & x_44006;
assign x_44008 = x_43519 & x_44007;
assign x_44009 = x_12716 & x_12717;
assign x_44010 = x_12715 & x_44009;
assign x_44011 = x_12718 & x_12719;
assign x_44012 = x_12720 & x_12721;
assign x_44013 = x_44011 & x_44012;
assign x_44014 = x_44010 & x_44013;
assign x_44015 = x_12722 & x_12723;
assign x_44016 = x_12724 & x_12725;
assign x_44017 = x_44015 & x_44016;
assign x_44018 = x_12726 & x_12727;
assign x_44019 = x_12728 & x_12729;
assign x_44020 = x_44018 & x_44019;
assign x_44021 = x_44017 & x_44020;
assign x_44022 = x_44014 & x_44021;
assign x_44023 = x_12731 & x_12732;
assign x_44024 = x_12730 & x_44023;
assign x_44025 = x_12733 & x_12734;
assign x_44026 = x_12735 & x_12736;
assign x_44027 = x_44025 & x_44026;
assign x_44028 = x_44024 & x_44027;
assign x_44029 = x_12737 & x_12738;
assign x_44030 = x_12739 & x_12740;
assign x_44031 = x_44029 & x_44030;
assign x_44032 = x_12741 & x_12742;
assign x_44033 = x_12743 & x_12744;
assign x_44034 = x_44032 & x_44033;
assign x_44035 = x_44031 & x_44034;
assign x_44036 = x_44028 & x_44035;
assign x_44037 = x_44022 & x_44036;
assign x_44038 = x_12746 & x_12747;
assign x_44039 = x_12745 & x_44038;
assign x_44040 = x_12748 & x_12749;
assign x_44041 = x_12750 & x_12751;
assign x_44042 = x_44040 & x_44041;
assign x_44043 = x_44039 & x_44042;
assign x_44044 = x_12752 & x_12753;
assign x_44045 = x_12754 & x_12755;
assign x_44046 = x_44044 & x_44045;
assign x_44047 = x_12756 & x_12757;
assign x_44048 = x_12758 & x_12759;
assign x_44049 = x_44047 & x_44048;
assign x_44050 = x_44046 & x_44049;
assign x_44051 = x_44043 & x_44050;
assign x_44052 = x_12760 & x_12761;
assign x_44053 = x_12762 & x_12763;
assign x_44054 = x_44052 & x_44053;
assign x_44055 = x_12764 & x_12765;
assign x_44056 = x_12766 & x_12767;
assign x_44057 = x_44055 & x_44056;
assign x_44058 = x_44054 & x_44057;
assign x_44059 = x_12768 & x_12769;
assign x_44060 = x_12770 & x_12771;
assign x_44061 = x_44059 & x_44060;
assign x_44062 = x_12772 & x_12773;
assign x_44063 = x_12774 & x_12775;
assign x_44064 = x_44062 & x_44063;
assign x_44065 = x_44061 & x_44064;
assign x_44066 = x_44058 & x_44065;
assign x_44067 = x_44051 & x_44066;
assign x_44068 = x_44037 & x_44067;
assign x_44069 = x_12777 & x_12778;
assign x_44070 = x_12776 & x_44069;
assign x_44071 = x_12779 & x_12780;
assign x_44072 = x_12781 & x_12782;
assign x_44073 = x_44071 & x_44072;
assign x_44074 = x_44070 & x_44073;
assign x_44075 = x_12783 & x_12784;
assign x_44076 = x_12785 & x_12786;
assign x_44077 = x_44075 & x_44076;
assign x_44078 = x_12787 & x_12788;
assign x_44079 = x_12789 & x_12790;
assign x_44080 = x_44078 & x_44079;
assign x_44081 = x_44077 & x_44080;
assign x_44082 = x_44074 & x_44081;
assign x_44083 = x_12792 & x_12793;
assign x_44084 = x_12791 & x_44083;
assign x_44085 = x_12794 & x_12795;
assign x_44086 = x_12796 & x_12797;
assign x_44087 = x_44085 & x_44086;
assign x_44088 = x_44084 & x_44087;
assign x_44089 = x_12798 & x_12799;
assign x_44090 = x_12800 & x_12801;
assign x_44091 = x_44089 & x_44090;
assign x_44092 = x_12802 & x_12803;
assign x_44093 = x_12804 & x_12805;
assign x_44094 = x_44092 & x_44093;
assign x_44095 = x_44091 & x_44094;
assign x_44096 = x_44088 & x_44095;
assign x_44097 = x_44082 & x_44096;
assign x_44098 = x_12807 & x_12808;
assign x_44099 = x_12806 & x_44098;
assign x_44100 = x_12809 & x_12810;
assign x_44101 = x_12811 & x_12812;
assign x_44102 = x_44100 & x_44101;
assign x_44103 = x_44099 & x_44102;
assign x_44104 = x_12813 & x_12814;
assign x_44105 = x_12815 & x_12816;
assign x_44106 = x_44104 & x_44105;
assign x_44107 = x_12817 & x_12818;
assign x_44108 = x_12819 & x_12820;
assign x_44109 = x_44107 & x_44108;
assign x_44110 = x_44106 & x_44109;
assign x_44111 = x_44103 & x_44110;
assign x_44112 = x_12821 & x_12822;
assign x_44113 = x_12823 & x_12824;
assign x_44114 = x_44112 & x_44113;
assign x_44115 = x_12825 & x_12826;
assign x_44116 = x_12827 & x_12828;
assign x_44117 = x_44115 & x_44116;
assign x_44118 = x_44114 & x_44117;
assign x_44119 = x_12829 & x_12830;
assign x_44120 = x_12831 & x_12832;
assign x_44121 = x_44119 & x_44120;
assign x_44122 = x_12833 & x_12834;
assign x_44123 = x_12835 & x_12836;
assign x_44124 = x_44122 & x_44123;
assign x_44125 = x_44121 & x_44124;
assign x_44126 = x_44118 & x_44125;
assign x_44127 = x_44111 & x_44126;
assign x_44128 = x_44097 & x_44127;
assign x_44129 = x_44068 & x_44128;
assign x_44130 = x_12838 & x_12839;
assign x_44131 = x_12837 & x_44130;
assign x_44132 = x_12840 & x_12841;
assign x_44133 = x_12842 & x_12843;
assign x_44134 = x_44132 & x_44133;
assign x_44135 = x_44131 & x_44134;
assign x_44136 = x_12844 & x_12845;
assign x_44137 = x_12846 & x_12847;
assign x_44138 = x_44136 & x_44137;
assign x_44139 = x_12848 & x_12849;
assign x_44140 = x_12850 & x_12851;
assign x_44141 = x_44139 & x_44140;
assign x_44142 = x_44138 & x_44141;
assign x_44143 = x_44135 & x_44142;
assign x_44144 = x_12853 & x_12854;
assign x_44145 = x_12852 & x_44144;
assign x_44146 = x_12855 & x_12856;
assign x_44147 = x_12857 & x_12858;
assign x_44148 = x_44146 & x_44147;
assign x_44149 = x_44145 & x_44148;
assign x_44150 = x_12859 & x_12860;
assign x_44151 = x_12861 & x_12862;
assign x_44152 = x_44150 & x_44151;
assign x_44153 = x_12863 & x_12864;
assign x_44154 = x_12865 & x_12866;
assign x_44155 = x_44153 & x_44154;
assign x_44156 = x_44152 & x_44155;
assign x_44157 = x_44149 & x_44156;
assign x_44158 = x_44143 & x_44157;
assign x_44159 = x_12868 & x_12869;
assign x_44160 = x_12867 & x_44159;
assign x_44161 = x_12870 & x_12871;
assign x_44162 = x_12872 & x_12873;
assign x_44163 = x_44161 & x_44162;
assign x_44164 = x_44160 & x_44163;
assign x_44165 = x_12874 & x_12875;
assign x_44166 = x_12876 & x_12877;
assign x_44167 = x_44165 & x_44166;
assign x_44168 = x_12878 & x_12879;
assign x_44169 = x_12880 & x_12881;
assign x_44170 = x_44168 & x_44169;
assign x_44171 = x_44167 & x_44170;
assign x_44172 = x_44164 & x_44171;
assign x_44173 = x_12882 & x_12883;
assign x_44174 = x_12884 & x_12885;
assign x_44175 = x_44173 & x_44174;
assign x_44176 = x_12886 & x_12887;
assign x_44177 = x_12888 & x_12889;
assign x_44178 = x_44176 & x_44177;
assign x_44179 = x_44175 & x_44178;
assign x_44180 = x_12890 & x_12891;
assign x_44181 = x_12892 & x_12893;
assign x_44182 = x_44180 & x_44181;
assign x_44183 = x_12894 & x_12895;
assign x_44184 = x_12896 & x_12897;
assign x_44185 = x_44183 & x_44184;
assign x_44186 = x_44182 & x_44185;
assign x_44187 = x_44179 & x_44186;
assign x_44188 = x_44172 & x_44187;
assign x_44189 = x_44158 & x_44188;
assign x_44190 = x_12899 & x_12900;
assign x_44191 = x_12898 & x_44190;
assign x_44192 = x_12901 & x_12902;
assign x_44193 = x_12903 & x_12904;
assign x_44194 = x_44192 & x_44193;
assign x_44195 = x_44191 & x_44194;
assign x_44196 = x_12905 & x_12906;
assign x_44197 = x_12907 & x_12908;
assign x_44198 = x_44196 & x_44197;
assign x_44199 = x_12909 & x_12910;
assign x_44200 = x_12911 & x_12912;
assign x_44201 = x_44199 & x_44200;
assign x_44202 = x_44198 & x_44201;
assign x_44203 = x_44195 & x_44202;
assign x_44204 = x_12914 & x_12915;
assign x_44205 = x_12913 & x_44204;
assign x_44206 = x_12916 & x_12917;
assign x_44207 = x_12918 & x_12919;
assign x_44208 = x_44206 & x_44207;
assign x_44209 = x_44205 & x_44208;
assign x_44210 = x_12920 & x_12921;
assign x_44211 = x_12922 & x_12923;
assign x_44212 = x_44210 & x_44211;
assign x_44213 = x_12924 & x_12925;
assign x_44214 = x_12926 & x_12927;
assign x_44215 = x_44213 & x_44214;
assign x_44216 = x_44212 & x_44215;
assign x_44217 = x_44209 & x_44216;
assign x_44218 = x_44203 & x_44217;
assign x_44219 = x_12929 & x_12930;
assign x_44220 = x_12928 & x_44219;
assign x_44221 = x_12931 & x_12932;
assign x_44222 = x_12933 & x_12934;
assign x_44223 = x_44221 & x_44222;
assign x_44224 = x_44220 & x_44223;
assign x_44225 = x_12935 & x_12936;
assign x_44226 = x_12937 & x_12938;
assign x_44227 = x_44225 & x_44226;
assign x_44228 = x_12939 & x_12940;
assign x_44229 = x_12941 & x_12942;
assign x_44230 = x_44228 & x_44229;
assign x_44231 = x_44227 & x_44230;
assign x_44232 = x_44224 & x_44231;
assign x_44233 = x_12943 & x_12944;
assign x_44234 = x_12945 & x_12946;
assign x_44235 = x_44233 & x_44234;
assign x_44236 = x_12947 & x_12948;
assign x_44237 = x_12949 & x_12950;
assign x_44238 = x_44236 & x_44237;
assign x_44239 = x_44235 & x_44238;
assign x_44240 = x_12951 & x_12952;
assign x_44241 = x_12953 & x_12954;
assign x_44242 = x_44240 & x_44241;
assign x_44243 = x_12955 & x_12956;
assign x_44244 = x_12957 & x_12958;
assign x_44245 = x_44243 & x_44244;
assign x_44246 = x_44242 & x_44245;
assign x_44247 = x_44239 & x_44246;
assign x_44248 = x_44232 & x_44247;
assign x_44249 = x_44218 & x_44248;
assign x_44250 = x_44189 & x_44249;
assign x_44251 = x_44129 & x_44250;
assign x_44252 = x_12960 & x_12961;
assign x_44253 = x_12959 & x_44252;
assign x_44254 = x_12962 & x_12963;
assign x_44255 = x_12964 & x_12965;
assign x_44256 = x_44254 & x_44255;
assign x_44257 = x_44253 & x_44256;
assign x_44258 = x_12966 & x_12967;
assign x_44259 = x_12968 & x_12969;
assign x_44260 = x_44258 & x_44259;
assign x_44261 = x_12970 & x_12971;
assign x_44262 = x_12972 & x_12973;
assign x_44263 = x_44261 & x_44262;
assign x_44264 = x_44260 & x_44263;
assign x_44265 = x_44257 & x_44264;
assign x_44266 = x_12975 & x_12976;
assign x_44267 = x_12974 & x_44266;
assign x_44268 = x_12977 & x_12978;
assign x_44269 = x_12979 & x_12980;
assign x_44270 = x_44268 & x_44269;
assign x_44271 = x_44267 & x_44270;
assign x_44272 = x_12981 & x_12982;
assign x_44273 = x_12983 & x_12984;
assign x_44274 = x_44272 & x_44273;
assign x_44275 = x_12985 & x_12986;
assign x_44276 = x_12987 & x_12988;
assign x_44277 = x_44275 & x_44276;
assign x_44278 = x_44274 & x_44277;
assign x_44279 = x_44271 & x_44278;
assign x_44280 = x_44265 & x_44279;
assign x_44281 = x_12990 & x_12991;
assign x_44282 = x_12989 & x_44281;
assign x_44283 = x_12992 & x_12993;
assign x_44284 = x_12994 & x_12995;
assign x_44285 = x_44283 & x_44284;
assign x_44286 = x_44282 & x_44285;
assign x_44287 = x_12996 & x_12997;
assign x_44288 = x_12998 & x_12999;
assign x_44289 = x_44287 & x_44288;
assign x_44290 = x_13000 & x_13001;
assign x_44291 = x_13002 & x_13003;
assign x_44292 = x_44290 & x_44291;
assign x_44293 = x_44289 & x_44292;
assign x_44294 = x_44286 & x_44293;
assign x_44295 = x_13004 & x_13005;
assign x_44296 = x_13006 & x_13007;
assign x_44297 = x_44295 & x_44296;
assign x_44298 = x_13008 & x_13009;
assign x_44299 = x_13010 & x_13011;
assign x_44300 = x_44298 & x_44299;
assign x_44301 = x_44297 & x_44300;
assign x_44302 = x_13012 & x_13013;
assign x_44303 = x_13014 & x_13015;
assign x_44304 = x_44302 & x_44303;
assign x_44305 = x_13016 & x_13017;
assign x_44306 = x_13018 & x_13019;
assign x_44307 = x_44305 & x_44306;
assign x_44308 = x_44304 & x_44307;
assign x_44309 = x_44301 & x_44308;
assign x_44310 = x_44294 & x_44309;
assign x_44311 = x_44280 & x_44310;
assign x_44312 = x_13021 & x_13022;
assign x_44313 = x_13020 & x_44312;
assign x_44314 = x_13023 & x_13024;
assign x_44315 = x_13025 & x_13026;
assign x_44316 = x_44314 & x_44315;
assign x_44317 = x_44313 & x_44316;
assign x_44318 = x_13027 & x_13028;
assign x_44319 = x_13029 & x_13030;
assign x_44320 = x_44318 & x_44319;
assign x_44321 = x_13031 & x_13032;
assign x_44322 = x_13033 & x_13034;
assign x_44323 = x_44321 & x_44322;
assign x_44324 = x_44320 & x_44323;
assign x_44325 = x_44317 & x_44324;
assign x_44326 = x_13036 & x_13037;
assign x_44327 = x_13035 & x_44326;
assign x_44328 = x_13038 & x_13039;
assign x_44329 = x_13040 & x_13041;
assign x_44330 = x_44328 & x_44329;
assign x_44331 = x_44327 & x_44330;
assign x_44332 = x_13042 & x_13043;
assign x_44333 = x_13044 & x_13045;
assign x_44334 = x_44332 & x_44333;
assign x_44335 = x_13046 & x_13047;
assign x_44336 = x_13048 & x_13049;
assign x_44337 = x_44335 & x_44336;
assign x_44338 = x_44334 & x_44337;
assign x_44339 = x_44331 & x_44338;
assign x_44340 = x_44325 & x_44339;
assign x_44341 = x_13051 & x_13052;
assign x_44342 = x_13050 & x_44341;
assign x_44343 = x_13053 & x_13054;
assign x_44344 = x_13055 & x_13056;
assign x_44345 = x_44343 & x_44344;
assign x_44346 = x_44342 & x_44345;
assign x_44347 = x_13057 & x_13058;
assign x_44348 = x_13059 & x_13060;
assign x_44349 = x_44347 & x_44348;
assign x_44350 = x_13061 & x_13062;
assign x_44351 = x_13063 & x_13064;
assign x_44352 = x_44350 & x_44351;
assign x_44353 = x_44349 & x_44352;
assign x_44354 = x_44346 & x_44353;
assign x_44355 = x_13065 & x_13066;
assign x_44356 = x_13067 & x_13068;
assign x_44357 = x_44355 & x_44356;
assign x_44358 = x_13069 & x_13070;
assign x_44359 = x_13071 & x_13072;
assign x_44360 = x_44358 & x_44359;
assign x_44361 = x_44357 & x_44360;
assign x_44362 = x_13073 & x_13074;
assign x_44363 = x_13075 & x_13076;
assign x_44364 = x_44362 & x_44363;
assign x_44365 = x_13077 & x_13078;
assign x_44366 = x_13079 & x_13080;
assign x_44367 = x_44365 & x_44366;
assign x_44368 = x_44364 & x_44367;
assign x_44369 = x_44361 & x_44368;
assign x_44370 = x_44354 & x_44369;
assign x_44371 = x_44340 & x_44370;
assign x_44372 = x_44311 & x_44371;
assign x_44373 = x_13082 & x_13083;
assign x_44374 = x_13081 & x_44373;
assign x_44375 = x_13084 & x_13085;
assign x_44376 = x_13086 & x_13087;
assign x_44377 = x_44375 & x_44376;
assign x_44378 = x_44374 & x_44377;
assign x_44379 = x_13088 & x_13089;
assign x_44380 = x_13090 & x_13091;
assign x_44381 = x_44379 & x_44380;
assign x_44382 = x_13092 & x_13093;
assign x_44383 = x_13094 & x_13095;
assign x_44384 = x_44382 & x_44383;
assign x_44385 = x_44381 & x_44384;
assign x_44386 = x_44378 & x_44385;
assign x_44387 = x_13097 & x_13098;
assign x_44388 = x_13096 & x_44387;
assign x_44389 = x_13099 & x_13100;
assign x_44390 = x_13101 & x_13102;
assign x_44391 = x_44389 & x_44390;
assign x_44392 = x_44388 & x_44391;
assign x_44393 = x_13103 & x_13104;
assign x_44394 = x_13105 & x_13106;
assign x_44395 = x_44393 & x_44394;
assign x_44396 = x_13107 & x_13108;
assign x_44397 = x_13109 & x_13110;
assign x_44398 = x_44396 & x_44397;
assign x_44399 = x_44395 & x_44398;
assign x_44400 = x_44392 & x_44399;
assign x_44401 = x_44386 & x_44400;
assign x_44402 = x_13112 & x_13113;
assign x_44403 = x_13111 & x_44402;
assign x_44404 = x_13114 & x_13115;
assign x_44405 = x_13116 & x_13117;
assign x_44406 = x_44404 & x_44405;
assign x_44407 = x_44403 & x_44406;
assign x_44408 = x_13118 & x_13119;
assign x_44409 = x_13120 & x_13121;
assign x_44410 = x_44408 & x_44409;
assign x_44411 = x_13122 & x_13123;
assign x_44412 = x_13124 & x_13125;
assign x_44413 = x_44411 & x_44412;
assign x_44414 = x_44410 & x_44413;
assign x_44415 = x_44407 & x_44414;
assign x_44416 = x_13126 & x_13127;
assign x_44417 = x_13128 & x_13129;
assign x_44418 = x_44416 & x_44417;
assign x_44419 = x_13130 & x_13131;
assign x_44420 = x_13132 & x_13133;
assign x_44421 = x_44419 & x_44420;
assign x_44422 = x_44418 & x_44421;
assign x_44423 = x_13134 & x_13135;
assign x_44424 = x_13136 & x_13137;
assign x_44425 = x_44423 & x_44424;
assign x_44426 = x_13138 & x_13139;
assign x_44427 = x_13140 & x_13141;
assign x_44428 = x_44426 & x_44427;
assign x_44429 = x_44425 & x_44428;
assign x_44430 = x_44422 & x_44429;
assign x_44431 = x_44415 & x_44430;
assign x_44432 = x_44401 & x_44431;
assign x_44433 = x_13143 & x_13144;
assign x_44434 = x_13142 & x_44433;
assign x_44435 = x_13145 & x_13146;
assign x_44436 = x_13147 & x_13148;
assign x_44437 = x_44435 & x_44436;
assign x_44438 = x_44434 & x_44437;
assign x_44439 = x_13149 & x_13150;
assign x_44440 = x_13151 & x_13152;
assign x_44441 = x_44439 & x_44440;
assign x_44442 = x_13153 & x_13154;
assign x_44443 = x_13155 & x_13156;
assign x_44444 = x_44442 & x_44443;
assign x_44445 = x_44441 & x_44444;
assign x_44446 = x_44438 & x_44445;
assign x_44447 = x_13157 & x_13158;
assign x_44448 = x_13159 & x_13160;
assign x_44449 = x_44447 & x_44448;
assign x_44450 = x_13161 & x_13162;
assign x_44451 = x_13163 & x_13164;
assign x_44452 = x_44450 & x_44451;
assign x_44453 = x_44449 & x_44452;
assign x_44454 = x_13165 & x_13166;
assign x_44455 = x_13167 & x_13168;
assign x_44456 = x_44454 & x_44455;
assign x_44457 = x_13169 & x_13170;
assign x_44458 = x_13171 & x_13172;
assign x_44459 = x_44457 & x_44458;
assign x_44460 = x_44456 & x_44459;
assign x_44461 = x_44453 & x_44460;
assign x_44462 = x_44446 & x_44461;
assign x_44463 = x_13174 & x_13175;
assign x_44464 = x_13173 & x_44463;
assign x_44465 = x_13176 & x_13177;
assign x_44466 = x_13178 & x_13179;
assign x_44467 = x_44465 & x_44466;
assign x_44468 = x_44464 & x_44467;
assign x_44469 = x_13180 & x_13181;
assign x_44470 = x_13182 & x_13183;
assign x_44471 = x_44469 & x_44470;
assign x_44472 = x_13184 & x_13185;
assign x_44473 = x_13186 & x_13187;
assign x_44474 = x_44472 & x_44473;
assign x_44475 = x_44471 & x_44474;
assign x_44476 = x_44468 & x_44475;
assign x_44477 = x_13188 & x_13189;
assign x_44478 = x_13190 & x_13191;
assign x_44479 = x_44477 & x_44478;
assign x_44480 = x_13192 & x_13193;
assign x_44481 = x_13194 & x_13195;
assign x_44482 = x_44480 & x_44481;
assign x_44483 = x_44479 & x_44482;
assign x_44484 = x_13196 & x_13197;
assign x_44485 = x_13198 & x_13199;
assign x_44486 = x_44484 & x_44485;
assign x_44487 = x_13200 & x_13201;
assign x_44488 = x_13202 & x_13203;
assign x_44489 = x_44487 & x_44488;
assign x_44490 = x_44486 & x_44489;
assign x_44491 = x_44483 & x_44490;
assign x_44492 = x_44476 & x_44491;
assign x_44493 = x_44462 & x_44492;
assign x_44494 = x_44432 & x_44493;
assign x_44495 = x_44372 & x_44494;
assign x_44496 = x_44251 & x_44495;
assign x_44497 = x_13205 & x_13206;
assign x_44498 = x_13204 & x_44497;
assign x_44499 = x_13207 & x_13208;
assign x_44500 = x_13209 & x_13210;
assign x_44501 = x_44499 & x_44500;
assign x_44502 = x_44498 & x_44501;
assign x_44503 = x_13211 & x_13212;
assign x_44504 = x_13213 & x_13214;
assign x_44505 = x_44503 & x_44504;
assign x_44506 = x_13215 & x_13216;
assign x_44507 = x_13217 & x_13218;
assign x_44508 = x_44506 & x_44507;
assign x_44509 = x_44505 & x_44508;
assign x_44510 = x_44502 & x_44509;
assign x_44511 = x_13220 & x_13221;
assign x_44512 = x_13219 & x_44511;
assign x_44513 = x_13222 & x_13223;
assign x_44514 = x_13224 & x_13225;
assign x_44515 = x_44513 & x_44514;
assign x_44516 = x_44512 & x_44515;
assign x_44517 = x_13226 & x_13227;
assign x_44518 = x_13228 & x_13229;
assign x_44519 = x_44517 & x_44518;
assign x_44520 = x_13230 & x_13231;
assign x_44521 = x_13232 & x_13233;
assign x_44522 = x_44520 & x_44521;
assign x_44523 = x_44519 & x_44522;
assign x_44524 = x_44516 & x_44523;
assign x_44525 = x_44510 & x_44524;
assign x_44526 = x_13235 & x_13236;
assign x_44527 = x_13234 & x_44526;
assign x_44528 = x_13237 & x_13238;
assign x_44529 = x_13239 & x_13240;
assign x_44530 = x_44528 & x_44529;
assign x_44531 = x_44527 & x_44530;
assign x_44532 = x_13241 & x_13242;
assign x_44533 = x_13243 & x_13244;
assign x_44534 = x_44532 & x_44533;
assign x_44535 = x_13245 & x_13246;
assign x_44536 = x_13247 & x_13248;
assign x_44537 = x_44535 & x_44536;
assign x_44538 = x_44534 & x_44537;
assign x_44539 = x_44531 & x_44538;
assign x_44540 = x_13249 & x_13250;
assign x_44541 = x_13251 & x_13252;
assign x_44542 = x_44540 & x_44541;
assign x_44543 = x_13253 & x_13254;
assign x_44544 = x_13255 & x_13256;
assign x_44545 = x_44543 & x_44544;
assign x_44546 = x_44542 & x_44545;
assign x_44547 = x_13257 & x_13258;
assign x_44548 = x_13259 & x_13260;
assign x_44549 = x_44547 & x_44548;
assign x_44550 = x_13261 & x_13262;
assign x_44551 = x_13263 & x_13264;
assign x_44552 = x_44550 & x_44551;
assign x_44553 = x_44549 & x_44552;
assign x_44554 = x_44546 & x_44553;
assign x_44555 = x_44539 & x_44554;
assign x_44556 = x_44525 & x_44555;
assign x_44557 = x_13266 & x_13267;
assign x_44558 = x_13265 & x_44557;
assign x_44559 = x_13268 & x_13269;
assign x_44560 = x_13270 & x_13271;
assign x_44561 = x_44559 & x_44560;
assign x_44562 = x_44558 & x_44561;
assign x_44563 = x_13272 & x_13273;
assign x_44564 = x_13274 & x_13275;
assign x_44565 = x_44563 & x_44564;
assign x_44566 = x_13276 & x_13277;
assign x_44567 = x_13278 & x_13279;
assign x_44568 = x_44566 & x_44567;
assign x_44569 = x_44565 & x_44568;
assign x_44570 = x_44562 & x_44569;
assign x_44571 = x_13281 & x_13282;
assign x_44572 = x_13280 & x_44571;
assign x_44573 = x_13283 & x_13284;
assign x_44574 = x_13285 & x_13286;
assign x_44575 = x_44573 & x_44574;
assign x_44576 = x_44572 & x_44575;
assign x_44577 = x_13287 & x_13288;
assign x_44578 = x_13289 & x_13290;
assign x_44579 = x_44577 & x_44578;
assign x_44580 = x_13291 & x_13292;
assign x_44581 = x_13293 & x_13294;
assign x_44582 = x_44580 & x_44581;
assign x_44583 = x_44579 & x_44582;
assign x_44584 = x_44576 & x_44583;
assign x_44585 = x_44570 & x_44584;
assign x_44586 = x_13296 & x_13297;
assign x_44587 = x_13295 & x_44586;
assign x_44588 = x_13298 & x_13299;
assign x_44589 = x_13300 & x_13301;
assign x_44590 = x_44588 & x_44589;
assign x_44591 = x_44587 & x_44590;
assign x_44592 = x_13302 & x_13303;
assign x_44593 = x_13304 & x_13305;
assign x_44594 = x_44592 & x_44593;
assign x_44595 = x_13306 & x_13307;
assign x_44596 = x_13308 & x_13309;
assign x_44597 = x_44595 & x_44596;
assign x_44598 = x_44594 & x_44597;
assign x_44599 = x_44591 & x_44598;
assign x_44600 = x_13310 & x_13311;
assign x_44601 = x_13312 & x_13313;
assign x_44602 = x_44600 & x_44601;
assign x_44603 = x_13314 & x_13315;
assign x_44604 = x_13316 & x_13317;
assign x_44605 = x_44603 & x_44604;
assign x_44606 = x_44602 & x_44605;
assign x_44607 = x_13318 & x_13319;
assign x_44608 = x_13320 & x_13321;
assign x_44609 = x_44607 & x_44608;
assign x_44610 = x_13322 & x_13323;
assign x_44611 = x_13324 & x_13325;
assign x_44612 = x_44610 & x_44611;
assign x_44613 = x_44609 & x_44612;
assign x_44614 = x_44606 & x_44613;
assign x_44615 = x_44599 & x_44614;
assign x_44616 = x_44585 & x_44615;
assign x_44617 = x_44556 & x_44616;
assign x_44618 = x_13327 & x_13328;
assign x_44619 = x_13326 & x_44618;
assign x_44620 = x_13329 & x_13330;
assign x_44621 = x_13331 & x_13332;
assign x_44622 = x_44620 & x_44621;
assign x_44623 = x_44619 & x_44622;
assign x_44624 = x_13333 & x_13334;
assign x_44625 = x_13335 & x_13336;
assign x_44626 = x_44624 & x_44625;
assign x_44627 = x_13337 & x_13338;
assign x_44628 = x_13339 & x_13340;
assign x_44629 = x_44627 & x_44628;
assign x_44630 = x_44626 & x_44629;
assign x_44631 = x_44623 & x_44630;
assign x_44632 = x_13342 & x_13343;
assign x_44633 = x_13341 & x_44632;
assign x_44634 = x_13344 & x_13345;
assign x_44635 = x_13346 & x_13347;
assign x_44636 = x_44634 & x_44635;
assign x_44637 = x_44633 & x_44636;
assign x_44638 = x_13348 & x_13349;
assign x_44639 = x_13350 & x_13351;
assign x_44640 = x_44638 & x_44639;
assign x_44641 = x_13352 & x_13353;
assign x_44642 = x_13354 & x_13355;
assign x_44643 = x_44641 & x_44642;
assign x_44644 = x_44640 & x_44643;
assign x_44645 = x_44637 & x_44644;
assign x_44646 = x_44631 & x_44645;
assign x_44647 = x_13357 & x_13358;
assign x_44648 = x_13356 & x_44647;
assign x_44649 = x_13359 & x_13360;
assign x_44650 = x_13361 & x_13362;
assign x_44651 = x_44649 & x_44650;
assign x_44652 = x_44648 & x_44651;
assign x_44653 = x_13363 & x_13364;
assign x_44654 = x_13365 & x_13366;
assign x_44655 = x_44653 & x_44654;
assign x_44656 = x_13367 & x_13368;
assign x_44657 = x_13369 & x_13370;
assign x_44658 = x_44656 & x_44657;
assign x_44659 = x_44655 & x_44658;
assign x_44660 = x_44652 & x_44659;
assign x_44661 = x_13371 & x_13372;
assign x_44662 = x_13373 & x_13374;
assign x_44663 = x_44661 & x_44662;
assign x_44664 = x_13375 & x_13376;
assign x_44665 = x_13377 & x_13378;
assign x_44666 = x_44664 & x_44665;
assign x_44667 = x_44663 & x_44666;
assign x_44668 = x_13379 & x_13380;
assign x_44669 = x_13381 & x_13382;
assign x_44670 = x_44668 & x_44669;
assign x_44671 = x_13383 & x_13384;
assign x_44672 = x_13385 & x_13386;
assign x_44673 = x_44671 & x_44672;
assign x_44674 = x_44670 & x_44673;
assign x_44675 = x_44667 & x_44674;
assign x_44676 = x_44660 & x_44675;
assign x_44677 = x_44646 & x_44676;
assign x_44678 = x_13388 & x_13389;
assign x_44679 = x_13387 & x_44678;
assign x_44680 = x_13390 & x_13391;
assign x_44681 = x_13392 & x_13393;
assign x_44682 = x_44680 & x_44681;
assign x_44683 = x_44679 & x_44682;
assign x_44684 = x_13394 & x_13395;
assign x_44685 = x_13396 & x_13397;
assign x_44686 = x_44684 & x_44685;
assign x_44687 = x_13398 & x_13399;
assign x_44688 = x_13400 & x_13401;
assign x_44689 = x_44687 & x_44688;
assign x_44690 = x_44686 & x_44689;
assign x_44691 = x_44683 & x_44690;
assign x_44692 = x_13403 & x_13404;
assign x_44693 = x_13402 & x_44692;
assign x_44694 = x_13405 & x_13406;
assign x_44695 = x_13407 & x_13408;
assign x_44696 = x_44694 & x_44695;
assign x_44697 = x_44693 & x_44696;
assign x_44698 = x_13409 & x_13410;
assign x_44699 = x_13411 & x_13412;
assign x_44700 = x_44698 & x_44699;
assign x_44701 = x_13413 & x_13414;
assign x_44702 = x_13415 & x_13416;
assign x_44703 = x_44701 & x_44702;
assign x_44704 = x_44700 & x_44703;
assign x_44705 = x_44697 & x_44704;
assign x_44706 = x_44691 & x_44705;
assign x_44707 = x_13418 & x_13419;
assign x_44708 = x_13417 & x_44707;
assign x_44709 = x_13420 & x_13421;
assign x_44710 = x_13422 & x_13423;
assign x_44711 = x_44709 & x_44710;
assign x_44712 = x_44708 & x_44711;
assign x_44713 = x_13424 & x_13425;
assign x_44714 = x_13426 & x_13427;
assign x_44715 = x_44713 & x_44714;
assign x_44716 = x_13428 & x_13429;
assign x_44717 = x_13430 & x_13431;
assign x_44718 = x_44716 & x_44717;
assign x_44719 = x_44715 & x_44718;
assign x_44720 = x_44712 & x_44719;
assign x_44721 = x_13432 & x_13433;
assign x_44722 = x_13434 & x_13435;
assign x_44723 = x_44721 & x_44722;
assign x_44724 = x_13436 & x_13437;
assign x_44725 = x_13438 & x_13439;
assign x_44726 = x_44724 & x_44725;
assign x_44727 = x_44723 & x_44726;
assign x_44728 = x_13440 & x_13441;
assign x_44729 = x_13442 & x_13443;
assign x_44730 = x_44728 & x_44729;
assign x_44731 = x_13444 & x_13445;
assign x_44732 = x_13446 & x_13447;
assign x_44733 = x_44731 & x_44732;
assign x_44734 = x_44730 & x_44733;
assign x_44735 = x_44727 & x_44734;
assign x_44736 = x_44720 & x_44735;
assign x_44737 = x_44706 & x_44736;
assign x_44738 = x_44677 & x_44737;
assign x_44739 = x_44617 & x_44738;
assign x_44740 = x_13449 & x_13450;
assign x_44741 = x_13448 & x_44740;
assign x_44742 = x_13451 & x_13452;
assign x_44743 = x_13453 & x_13454;
assign x_44744 = x_44742 & x_44743;
assign x_44745 = x_44741 & x_44744;
assign x_44746 = x_13455 & x_13456;
assign x_44747 = x_13457 & x_13458;
assign x_44748 = x_44746 & x_44747;
assign x_44749 = x_13459 & x_13460;
assign x_44750 = x_13461 & x_13462;
assign x_44751 = x_44749 & x_44750;
assign x_44752 = x_44748 & x_44751;
assign x_44753 = x_44745 & x_44752;
assign x_44754 = x_13464 & x_13465;
assign x_44755 = x_13463 & x_44754;
assign x_44756 = x_13466 & x_13467;
assign x_44757 = x_13468 & x_13469;
assign x_44758 = x_44756 & x_44757;
assign x_44759 = x_44755 & x_44758;
assign x_44760 = x_13470 & x_13471;
assign x_44761 = x_13472 & x_13473;
assign x_44762 = x_44760 & x_44761;
assign x_44763 = x_13474 & x_13475;
assign x_44764 = x_13476 & x_13477;
assign x_44765 = x_44763 & x_44764;
assign x_44766 = x_44762 & x_44765;
assign x_44767 = x_44759 & x_44766;
assign x_44768 = x_44753 & x_44767;
assign x_44769 = x_13479 & x_13480;
assign x_44770 = x_13478 & x_44769;
assign x_44771 = x_13481 & x_13482;
assign x_44772 = x_13483 & x_13484;
assign x_44773 = x_44771 & x_44772;
assign x_44774 = x_44770 & x_44773;
assign x_44775 = x_13485 & x_13486;
assign x_44776 = x_13487 & x_13488;
assign x_44777 = x_44775 & x_44776;
assign x_44778 = x_13489 & x_13490;
assign x_44779 = x_13491 & x_13492;
assign x_44780 = x_44778 & x_44779;
assign x_44781 = x_44777 & x_44780;
assign x_44782 = x_44774 & x_44781;
assign x_44783 = x_13493 & x_13494;
assign x_44784 = x_13495 & x_13496;
assign x_44785 = x_44783 & x_44784;
assign x_44786 = x_13497 & x_13498;
assign x_44787 = x_13499 & x_13500;
assign x_44788 = x_44786 & x_44787;
assign x_44789 = x_44785 & x_44788;
assign x_44790 = x_13501 & x_13502;
assign x_44791 = x_13503 & x_13504;
assign x_44792 = x_44790 & x_44791;
assign x_44793 = x_13505 & x_13506;
assign x_44794 = x_13507 & x_13508;
assign x_44795 = x_44793 & x_44794;
assign x_44796 = x_44792 & x_44795;
assign x_44797 = x_44789 & x_44796;
assign x_44798 = x_44782 & x_44797;
assign x_44799 = x_44768 & x_44798;
assign x_44800 = x_13510 & x_13511;
assign x_44801 = x_13509 & x_44800;
assign x_44802 = x_13512 & x_13513;
assign x_44803 = x_13514 & x_13515;
assign x_44804 = x_44802 & x_44803;
assign x_44805 = x_44801 & x_44804;
assign x_44806 = x_13516 & x_13517;
assign x_44807 = x_13518 & x_13519;
assign x_44808 = x_44806 & x_44807;
assign x_44809 = x_13520 & x_13521;
assign x_44810 = x_13522 & x_13523;
assign x_44811 = x_44809 & x_44810;
assign x_44812 = x_44808 & x_44811;
assign x_44813 = x_44805 & x_44812;
assign x_44814 = x_13525 & x_13526;
assign x_44815 = x_13524 & x_44814;
assign x_44816 = x_13527 & x_13528;
assign x_44817 = x_13529 & x_13530;
assign x_44818 = x_44816 & x_44817;
assign x_44819 = x_44815 & x_44818;
assign x_44820 = x_13531 & x_13532;
assign x_44821 = x_13533 & x_13534;
assign x_44822 = x_44820 & x_44821;
assign x_44823 = x_13535 & x_13536;
assign x_44824 = x_13537 & x_13538;
assign x_44825 = x_44823 & x_44824;
assign x_44826 = x_44822 & x_44825;
assign x_44827 = x_44819 & x_44826;
assign x_44828 = x_44813 & x_44827;
assign x_44829 = x_13540 & x_13541;
assign x_44830 = x_13539 & x_44829;
assign x_44831 = x_13542 & x_13543;
assign x_44832 = x_13544 & x_13545;
assign x_44833 = x_44831 & x_44832;
assign x_44834 = x_44830 & x_44833;
assign x_44835 = x_13546 & x_13547;
assign x_44836 = x_13548 & x_13549;
assign x_44837 = x_44835 & x_44836;
assign x_44838 = x_13550 & x_13551;
assign x_44839 = x_13552 & x_13553;
assign x_44840 = x_44838 & x_44839;
assign x_44841 = x_44837 & x_44840;
assign x_44842 = x_44834 & x_44841;
assign x_44843 = x_13554 & x_13555;
assign x_44844 = x_13556 & x_13557;
assign x_44845 = x_44843 & x_44844;
assign x_44846 = x_13558 & x_13559;
assign x_44847 = x_13560 & x_13561;
assign x_44848 = x_44846 & x_44847;
assign x_44849 = x_44845 & x_44848;
assign x_44850 = x_13562 & x_13563;
assign x_44851 = x_13564 & x_13565;
assign x_44852 = x_44850 & x_44851;
assign x_44853 = x_13566 & x_13567;
assign x_44854 = x_13568 & x_13569;
assign x_44855 = x_44853 & x_44854;
assign x_44856 = x_44852 & x_44855;
assign x_44857 = x_44849 & x_44856;
assign x_44858 = x_44842 & x_44857;
assign x_44859 = x_44828 & x_44858;
assign x_44860 = x_44799 & x_44859;
assign x_44861 = x_13571 & x_13572;
assign x_44862 = x_13570 & x_44861;
assign x_44863 = x_13573 & x_13574;
assign x_44864 = x_13575 & x_13576;
assign x_44865 = x_44863 & x_44864;
assign x_44866 = x_44862 & x_44865;
assign x_44867 = x_13577 & x_13578;
assign x_44868 = x_13579 & x_13580;
assign x_44869 = x_44867 & x_44868;
assign x_44870 = x_13581 & x_13582;
assign x_44871 = x_13583 & x_13584;
assign x_44872 = x_44870 & x_44871;
assign x_44873 = x_44869 & x_44872;
assign x_44874 = x_44866 & x_44873;
assign x_44875 = x_13586 & x_13587;
assign x_44876 = x_13585 & x_44875;
assign x_44877 = x_13588 & x_13589;
assign x_44878 = x_13590 & x_13591;
assign x_44879 = x_44877 & x_44878;
assign x_44880 = x_44876 & x_44879;
assign x_44881 = x_13592 & x_13593;
assign x_44882 = x_13594 & x_13595;
assign x_44883 = x_44881 & x_44882;
assign x_44884 = x_13596 & x_13597;
assign x_44885 = x_13598 & x_13599;
assign x_44886 = x_44884 & x_44885;
assign x_44887 = x_44883 & x_44886;
assign x_44888 = x_44880 & x_44887;
assign x_44889 = x_44874 & x_44888;
assign x_44890 = x_13601 & x_13602;
assign x_44891 = x_13600 & x_44890;
assign x_44892 = x_13603 & x_13604;
assign x_44893 = x_13605 & x_13606;
assign x_44894 = x_44892 & x_44893;
assign x_44895 = x_44891 & x_44894;
assign x_44896 = x_13607 & x_13608;
assign x_44897 = x_13609 & x_13610;
assign x_44898 = x_44896 & x_44897;
assign x_44899 = x_13611 & x_13612;
assign x_44900 = x_13613 & x_13614;
assign x_44901 = x_44899 & x_44900;
assign x_44902 = x_44898 & x_44901;
assign x_44903 = x_44895 & x_44902;
assign x_44904 = x_13615 & x_13616;
assign x_44905 = x_13617 & x_13618;
assign x_44906 = x_44904 & x_44905;
assign x_44907 = x_13619 & x_13620;
assign x_44908 = x_13621 & x_13622;
assign x_44909 = x_44907 & x_44908;
assign x_44910 = x_44906 & x_44909;
assign x_44911 = x_13623 & x_13624;
assign x_44912 = x_13625 & x_13626;
assign x_44913 = x_44911 & x_44912;
assign x_44914 = x_13627 & x_13628;
assign x_44915 = x_13629 & x_13630;
assign x_44916 = x_44914 & x_44915;
assign x_44917 = x_44913 & x_44916;
assign x_44918 = x_44910 & x_44917;
assign x_44919 = x_44903 & x_44918;
assign x_44920 = x_44889 & x_44919;
assign x_44921 = x_13632 & x_13633;
assign x_44922 = x_13631 & x_44921;
assign x_44923 = x_13634 & x_13635;
assign x_44924 = x_13636 & x_13637;
assign x_44925 = x_44923 & x_44924;
assign x_44926 = x_44922 & x_44925;
assign x_44927 = x_13638 & x_13639;
assign x_44928 = x_13640 & x_13641;
assign x_44929 = x_44927 & x_44928;
assign x_44930 = x_13642 & x_13643;
assign x_44931 = x_13644 & x_13645;
assign x_44932 = x_44930 & x_44931;
assign x_44933 = x_44929 & x_44932;
assign x_44934 = x_44926 & x_44933;
assign x_44935 = x_13646 & x_13647;
assign x_44936 = x_13648 & x_13649;
assign x_44937 = x_44935 & x_44936;
assign x_44938 = x_13650 & x_13651;
assign x_44939 = x_13652 & x_13653;
assign x_44940 = x_44938 & x_44939;
assign x_44941 = x_44937 & x_44940;
assign x_44942 = x_13654 & x_13655;
assign x_44943 = x_13656 & x_13657;
assign x_44944 = x_44942 & x_44943;
assign x_44945 = x_13658 & x_13659;
assign x_44946 = x_13660 & x_13661;
assign x_44947 = x_44945 & x_44946;
assign x_44948 = x_44944 & x_44947;
assign x_44949 = x_44941 & x_44948;
assign x_44950 = x_44934 & x_44949;
assign x_44951 = x_13663 & x_13664;
assign x_44952 = x_13662 & x_44951;
assign x_44953 = x_13665 & x_13666;
assign x_44954 = x_13667 & x_13668;
assign x_44955 = x_44953 & x_44954;
assign x_44956 = x_44952 & x_44955;
assign x_44957 = x_13669 & x_13670;
assign x_44958 = x_13671 & x_13672;
assign x_44959 = x_44957 & x_44958;
assign x_44960 = x_13673 & x_13674;
assign x_44961 = x_13675 & x_13676;
assign x_44962 = x_44960 & x_44961;
assign x_44963 = x_44959 & x_44962;
assign x_44964 = x_44956 & x_44963;
assign x_44965 = x_13677 & x_13678;
assign x_44966 = x_13679 & x_13680;
assign x_44967 = x_44965 & x_44966;
assign x_44968 = x_13681 & x_13682;
assign x_44969 = x_13683 & x_13684;
assign x_44970 = x_44968 & x_44969;
assign x_44971 = x_44967 & x_44970;
assign x_44972 = x_13685 & x_13686;
assign x_44973 = x_13687 & x_13688;
assign x_44974 = x_44972 & x_44973;
assign x_44975 = x_13689 & x_13690;
assign x_44976 = x_13691 & x_13692;
assign x_44977 = x_44975 & x_44976;
assign x_44978 = x_44974 & x_44977;
assign x_44979 = x_44971 & x_44978;
assign x_44980 = x_44964 & x_44979;
assign x_44981 = x_44950 & x_44980;
assign x_44982 = x_44920 & x_44981;
assign x_44983 = x_44860 & x_44982;
assign x_44984 = x_44739 & x_44983;
assign x_44985 = x_44496 & x_44984;
assign x_44986 = x_44008 & x_44985;
assign x_44987 = x_13694 & x_13695;
assign x_44988 = x_13693 & x_44987;
assign x_44989 = x_13696 & x_13697;
assign x_44990 = x_13698 & x_13699;
assign x_44991 = x_44989 & x_44990;
assign x_44992 = x_44988 & x_44991;
assign x_44993 = x_13700 & x_13701;
assign x_44994 = x_13702 & x_13703;
assign x_44995 = x_44993 & x_44994;
assign x_44996 = x_13704 & x_13705;
assign x_44997 = x_13706 & x_13707;
assign x_44998 = x_44996 & x_44997;
assign x_44999 = x_44995 & x_44998;
assign x_45000 = x_44992 & x_44999;
assign x_45001 = x_13709 & x_13710;
assign x_45002 = x_13708 & x_45001;
assign x_45003 = x_13711 & x_13712;
assign x_45004 = x_13713 & x_13714;
assign x_45005 = x_45003 & x_45004;
assign x_45006 = x_45002 & x_45005;
assign x_45007 = x_13715 & x_13716;
assign x_45008 = x_13717 & x_13718;
assign x_45009 = x_45007 & x_45008;
assign x_45010 = x_13719 & x_13720;
assign x_45011 = x_13721 & x_13722;
assign x_45012 = x_45010 & x_45011;
assign x_45013 = x_45009 & x_45012;
assign x_45014 = x_45006 & x_45013;
assign x_45015 = x_45000 & x_45014;
assign x_45016 = x_13724 & x_13725;
assign x_45017 = x_13723 & x_45016;
assign x_45018 = x_13726 & x_13727;
assign x_45019 = x_13728 & x_13729;
assign x_45020 = x_45018 & x_45019;
assign x_45021 = x_45017 & x_45020;
assign x_45022 = x_13730 & x_13731;
assign x_45023 = x_13732 & x_13733;
assign x_45024 = x_45022 & x_45023;
assign x_45025 = x_13734 & x_13735;
assign x_45026 = x_13736 & x_13737;
assign x_45027 = x_45025 & x_45026;
assign x_45028 = x_45024 & x_45027;
assign x_45029 = x_45021 & x_45028;
assign x_45030 = x_13738 & x_13739;
assign x_45031 = x_13740 & x_13741;
assign x_45032 = x_45030 & x_45031;
assign x_45033 = x_13742 & x_13743;
assign x_45034 = x_13744 & x_13745;
assign x_45035 = x_45033 & x_45034;
assign x_45036 = x_45032 & x_45035;
assign x_45037 = x_13746 & x_13747;
assign x_45038 = x_13748 & x_13749;
assign x_45039 = x_45037 & x_45038;
assign x_45040 = x_13750 & x_13751;
assign x_45041 = x_13752 & x_13753;
assign x_45042 = x_45040 & x_45041;
assign x_45043 = x_45039 & x_45042;
assign x_45044 = x_45036 & x_45043;
assign x_45045 = x_45029 & x_45044;
assign x_45046 = x_45015 & x_45045;
assign x_45047 = x_13755 & x_13756;
assign x_45048 = x_13754 & x_45047;
assign x_45049 = x_13757 & x_13758;
assign x_45050 = x_13759 & x_13760;
assign x_45051 = x_45049 & x_45050;
assign x_45052 = x_45048 & x_45051;
assign x_45053 = x_13761 & x_13762;
assign x_45054 = x_13763 & x_13764;
assign x_45055 = x_45053 & x_45054;
assign x_45056 = x_13765 & x_13766;
assign x_45057 = x_13767 & x_13768;
assign x_45058 = x_45056 & x_45057;
assign x_45059 = x_45055 & x_45058;
assign x_45060 = x_45052 & x_45059;
assign x_45061 = x_13770 & x_13771;
assign x_45062 = x_13769 & x_45061;
assign x_45063 = x_13772 & x_13773;
assign x_45064 = x_13774 & x_13775;
assign x_45065 = x_45063 & x_45064;
assign x_45066 = x_45062 & x_45065;
assign x_45067 = x_13776 & x_13777;
assign x_45068 = x_13778 & x_13779;
assign x_45069 = x_45067 & x_45068;
assign x_45070 = x_13780 & x_13781;
assign x_45071 = x_13782 & x_13783;
assign x_45072 = x_45070 & x_45071;
assign x_45073 = x_45069 & x_45072;
assign x_45074 = x_45066 & x_45073;
assign x_45075 = x_45060 & x_45074;
assign x_45076 = x_13785 & x_13786;
assign x_45077 = x_13784 & x_45076;
assign x_45078 = x_13787 & x_13788;
assign x_45079 = x_13789 & x_13790;
assign x_45080 = x_45078 & x_45079;
assign x_45081 = x_45077 & x_45080;
assign x_45082 = x_13791 & x_13792;
assign x_45083 = x_13793 & x_13794;
assign x_45084 = x_45082 & x_45083;
assign x_45085 = x_13795 & x_13796;
assign x_45086 = x_13797 & x_13798;
assign x_45087 = x_45085 & x_45086;
assign x_45088 = x_45084 & x_45087;
assign x_45089 = x_45081 & x_45088;
assign x_45090 = x_13799 & x_13800;
assign x_45091 = x_13801 & x_13802;
assign x_45092 = x_45090 & x_45091;
assign x_45093 = x_13803 & x_13804;
assign x_45094 = x_13805 & x_13806;
assign x_45095 = x_45093 & x_45094;
assign x_45096 = x_45092 & x_45095;
assign x_45097 = x_13807 & x_13808;
assign x_45098 = x_13809 & x_13810;
assign x_45099 = x_45097 & x_45098;
assign x_45100 = x_13811 & x_13812;
assign x_45101 = x_13813 & x_13814;
assign x_45102 = x_45100 & x_45101;
assign x_45103 = x_45099 & x_45102;
assign x_45104 = x_45096 & x_45103;
assign x_45105 = x_45089 & x_45104;
assign x_45106 = x_45075 & x_45105;
assign x_45107 = x_45046 & x_45106;
assign x_45108 = x_13816 & x_13817;
assign x_45109 = x_13815 & x_45108;
assign x_45110 = x_13818 & x_13819;
assign x_45111 = x_13820 & x_13821;
assign x_45112 = x_45110 & x_45111;
assign x_45113 = x_45109 & x_45112;
assign x_45114 = x_13822 & x_13823;
assign x_45115 = x_13824 & x_13825;
assign x_45116 = x_45114 & x_45115;
assign x_45117 = x_13826 & x_13827;
assign x_45118 = x_13828 & x_13829;
assign x_45119 = x_45117 & x_45118;
assign x_45120 = x_45116 & x_45119;
assign x_45121 = x_45113 & x_45120;
assign x_45122 = x_13831 & x_13832;
assign x_45123 = x_13830 & x_45122;
assign x_45124 = x_13833 & x_13834;
assign x_45125 = x_13835 & x_13836;
assign x_45126 = x_45124 & x_45125;
assign x_45127 = x_45123 & x_45126;
assign x_45128 = x_13837 & x_13838;
assign x_45129 = x_13839 & x_13840;
assign x_45130 = x_45128 & x_45129;
assign x_45131 = x_13841 & x_13842;
assign x_45132 = x_13843 & x_13844;
assign x_45133 = x_45131 & x_45132;
assign x_45134 = x_45130 & x_45133;
assign x_45135 = x_45127 & x_45134;
assign x_45136 = x_45121 & x_45135;
assign x_45137 = x_13846 & x_13847;
assign x_45138 = x_13845 & x_45137;
assign x_45139 = x_13848 & x_13849;
assign x_45140 = x_13850 & x_13851;
assign x_45141 = x_45139 & x_45140;
assign x_45142 = x_45138 & x_45141;
assign x_45143 = x_13852 & x_13853;
assign x_45144 = x_13854 & x_13855;
assign x_45145 = x_45143 & x_45144;
assign x_45146 = x_13856 & x_13857;
assign x_45147 = x_13858 & x_13859;
assign x_45148 = x_45146 & x_45147;
assign x_45149 = x_45145 & x_45148;
assign x_45150 = x_45142 & x_45149;
assign x_45151 = x_13860 & x_13861;
assign x_45152 = x_13862 & x_13863;
assign x_45153 = x_45151 & x_45152;
assign x_45154 = x_13864 & x_13865;
assign x_45155 = x_13866 & x_13867;
assign x_45156 = x_45154 & x_45155;
assign x_45157 = x_45153 & x_45156;
assign x_45158 = x_13868 & x_13869;
assign x_45159 = x_13870 & x_13871;
assign x_45160 = x_45158 & x_45159;
assign x_45161 = x_13872 & x_13873;
assign x_45162 = x_13874 & x_13875;
assign x_45163 = x_45161 & x_45162;
assign x_45164 = x_45160 & x_45163;
assign x_45165 = x_45157 & x_45164;
assign x_45166 = x_45150 & x_45165;
assign x_45167 = x_45136 & x_45166;
assign x_45168 = x_13877 & x_13878;
assign x_45169 = x_13876 & x_45168;
assign x_45170 = x_13879 & x_13880;
assign x_45171 = x_13881 & x_13882;
assign x_45172 = x_45170 & x_45171;
assign x_45173 = x_45169 & x_45172;
assign x_45174 = x_13883 & x_13884;
assign x_45175 = x_13885 & x_13886;
assign x_45176 = x_45174 & x_45175;
assign x_45177 = x_13887 & x_13888;
assign x_45178 = x_13889 & x_13890;
assign x_45179 = x_45177 & x_45178;
assign x_45180 = x_45176 & x_45179;
assign x_45181 = x_45173 & x_45180;
assign x_45182 = x_13892 & x_13893;
assign x_45183 = x_13891 & x_45182;
assign x_45184 = x_13894 & x_13895;
assign x_45185 = x_13896 & x_13897;
assign x_45186 = x_45184 & x_45185;
assign x_45187 = x_45183 & x_45186;
assign x_45188 = x_13898 & x_13899;
assign x_45189 = x_13900 & x_13901;
assign x_45190 = x_45188 & x_45189;
assign x_45191 = x_13902 & x_13903;
assign x_45192 = x_13904 & x_13905;
assign x_45193 = x_45191 & x_45192;
assign x_45194 = x_45190 & x_45193;
assign x_45195 = x_45187 & x_45194;
assign x_45196 = x_45181 & x_45195;
assign x_45197 = x_13907 & x_13908;
assign x_45198 = x_13906 & x_45197;
assign x_45199 = x_13909 & x_13910;
assign x_45200 = x_13911 & x_13912;
assign x_45201 = x_45199 & x_45200;
assign x_45202 = x_45198 & x_45201;
assign x_45203 = x_13913 & x_13914;
assign x_45204 = x_13915 & x_13916;
assign x_45205 = x_45203 & x_45204;
assign x_45206 = x_13917 & x_13918;
assign x_45207 = x_13919 & x_13920;
assign x_45208 = x_45206 & x_45207;
assign x_45209 = x_45205 & x_45208;
assign x_45210 = x_45202 & x_45209;
assign x_45211 = x_13921 & x_13922;
assign x_45212 = x_13923 & x_13924;
assign x_45213 = x_45211 & x_45212;
assign x_45214 = x_13925 & x_13926;
assign x_45215 = x_13927 & x_13928;
assign x_45216 = x_45214 & x_45215;
assign x_45217 = x_45213 & x_45216;
assign x_45218 = x_13929 & x_13930;
assign x_45219 = x_13931 & x_13932;
assign x_45220 = x_45218 & x_45219;
assign x_45221 = x_13933 & x_13934;
assign x_45222 = x_13935 & x_13936;
assign x_45223 = x_45221 & x_45222;
assign x_45224 = x_45220 & x_45223;
assign x_45225 = x_45217 & x_45224;
assign x_45226 = x_45210 & x_45225;
assign x_45227 = x_45196 & x_45226;
assign x_45228 = x_45167 & x_45227;
assign x_45229 = x_45107 & x_45228;
assign x_45230 = x_13938 & x_13939;
assign x_45231 = x_13937 & x_45230;
assign x_45232 = x_13940 & x_13941;
assign x_45233 = x_13942 & x_13943;
assign x_45234 = x_45232 & x_45233;
assign x_45235 = x_45231 & x_45234;
assign x_45236 = x_13944 & x_13945;
assign x_45237 = x_13946 & x_13947;
assign x_45238 = x_45236 & x_45237;
assign x_45239 = x_13948 & x_13949;
assign x_45240 = x_13950 & x_13951;
assign x_45241 = x_45239 & x_45240;
assign x_45242 = x_45238 & x_45241;
assign x_45243 = x_45235 & x_45242;
assign x_45244 = x_13953 & x_13954;
assign x_45245 = x_13952 & x_45244;
assign x_45246 = x_13955 & x_13956;
assign x_45247 = x_13957 & x_13958;
assign x_45248 = x_45246 & x_45247;
assign x_45249 = x_45245 & x_45248;
assign x_45250 = x_13959 & x_13960;
assign x_45251 = x_13961 & x_13962;
assign x_45252 = x_45250 & x_45251;
assign x_45253 = x_13963 & x_13964;
assign x_45254 = x_13965 & x_13966;
assign x_45255 = x_45253 & x_45254;
assign x_45256 = x_45252 & x_45255;
assign x_45257 = x_45249 & x_45256;
assign x_45258 = x_45243 & x_45257;
assign x_45259 = x_13968 & x_13969;
assign x_45260 = x_13967 & x_45259;
assign x_45261 = x_13970 & x_13971;
assign x_45262 = x_13972 & x_13973;
assign x_45263 = x_45261 & x_45262;
assign x_45264 = x_45260 & x_45263;
assign x_45265 = x_13974 & x_13975;
assign x_45266 = x_13976 & x_13977;
assign x_45267 = x_45265 & x_45266;
assign x_45268 = x_13978 & x_13979;
assign x_45269 = x_13980 & x_13981;
assign x_45270 = x_45268 & x_45269;
assign x_45271 = x_45267 & x_45270;
assign x_45272 = x_45264 & x_45271;
assign x_45273 = x_13982 & x_13983;
assign x_45274 = x_13984 & x_13985;
assign x_45275 = x_45273 & x_45274;
assign x_45276 = x_13986 & x_13987;
assign x_45277 = x_13988 & x_13989;
assign x_45278 = x_45276 & x_45277;
assign x_45279 = x_45275 & x_45278;
assign x_45280 = x_13990 & x_13991;
assign x_45281 = x_13992 & x_13993;
assign x_45282 = x_45280 & x_45281;
assign x_45283 = x_13994 & x_13995;
assign x_45284 = x_13996 & x_13997;
assign x_45285 = x_45283 & x_45284;
assign x_45286 = x_45282 & x_45285;
assign x_45287 = x_45279 & x_45286;
assign x_45288 = x_45272 & x_45287;
assign x_45289 = x_45258 & x_45288;
assign x_45290 = x_13999 & x_14000;
assign x_45291 = x_13998 & x_45290;
assign x_45292 = x_14001 & x_14002;
assign x_45293 = x_14003 & x_14004;
assign x_45294 = x_45292 & x_45293;
assign x_45295 = x_45291 & x_45294;
assign x_45296 = x_14005 & x_14006;
assign x_45297 = x_14007 & x_14008;
assign x_45298 = x_45296 & x_45297;
assign x_45299 = x_14009 & x_14010;
assign x_45300 = x_14011 & x_14012;
assign x_45301 = x_45299 & x_45300;
assign x_45302 = x_45298 & x_45301;
assign x_45303 = x_45295 & x_45302;
assign x_45304 = x_14014 & x_14015;
assign x_45305 = x_14013 & x_45304;
assign x_45306 = x_14016 & x_14017;
assign x_45307 = x_14018 & x_14019;
assign x_45308 = x_45306 & x_45307;
assign x_45309 = x_45305 & x_45308;
assign x_45310 = x_14020 & x_14021;
assign x_45311 = x_14022 & x_14023;
assign x_45312 = x_45310 & x_45311;
assign x_45313 = x_14024 & x_14025;
assign x_45314 = x_14026 & x_14027;
assign x_45315 = x_45313 & x_45314;
assign x_45316 = x_45312 & x_45315;
assign x_45317 = x_45309 & x_45316;
assign x_45318 = x_45303 & x_45317;
assign x_45319 = x_14029 & x_14030;
assign x_45320 = x_14028 & x_45319;
assign x_45321 = x_14031 & x_14032;
assign x_45322 = x_14033 & x_14034;
assign x_45323 = x_45321 & x_45322;
assign x_45324 = x_45320 & x_45323;
assign x_45325 = x_14035 & x_14036;
assign x_45326 = x_14037 & x_14038;
assign x_45327 = x_45325 & x_45326;
assign x_45328 = x_14039 & x_14040;
assign x_45329 = x_14041 & x_14042;
assign x_45330 = x_45328 & x_45329;
assign x_45331 = x_45327 & x_45330;
assign x_45332 = x_45324 & x_45331;
assign x_45333 = x_14043 & x_14044;
assign x_45334 = x_14045 & x_14046;
assign x_45335 = x_45333 & x_45334;
assign x_45336 = x_14047 & x_14048;
assign x_45337 = x_14049 & x_14050;
assign x_45338 = x_45336 & x_45337;
assign x_45339 = x_45335 & x_45338;
assign x_45340 = x_14051 & x_14052;
assign x_45341 = x_14053 & x_14054;
assign x_45342 = x_45340 & x_45341;
assign x_45343 = x_14055 & x_14056;
assign x_45344 = x_14057 & x_14058;
assign x_45345 = x_45343 & x_45344;
assign x_45346 = x_45342 & x_45345;
assign x_45347 = x_45339 & x_45346;
assign x_45348 = x_45332 & x_45347;
assign x_45349 = x_45318 & x_45348;
assign x_45350 = x_45289 & x_45349;
assign x_45351 = x_14060 & x_14061;
assign x_45352 = x_14059 & x_45351;
assign x_45353 = x_14062 & x_14063;
assign x_45354 = x_14064 & x_14065;
assign x_45355 = x_45353 & x_45354;
assign x_45356 = x_45352 & x_45355;
assign x_45357 = x_14066 & x_14067;
assign x_45358 = x_14068 & x_14069;
assign x_45359 = x_45357 & x_45358;
assign x_45360 = x_14070 & x_14071;
assign x_45361 = x_14072 & x_14073;
assign x_45362 = x_45360 & x_45361;
assign x_45363 = x_45359 & x_45362;
assign x_45364 = x_45356 & x_45363;
assign x_45365 = x_14075 & x_14076;
assign x_45366 = x_14074 & x_45365;
assign x_45367 = x_14077 & x_14078;
assign x_45368 = x_14079 & x_14080;
assign x_45369 = x_45367 & x_45368;
assign x_45370 = x_45366 & x_45369;
assign x_45371 = x_14081 & x_14082;
assign x_45372 = x_14083 & x_14084;
assign x_45373 = x_45371 & x_45372;
assign x_45374 = x_14085 & x_14086;
assign x_45375 = x_14087 & x_14088;
assign x_45376 = x_45374 & x_45375;
assign x_45377 = x_45373 & x_45376;
assign x_45378 = x_45370 & x_45377;
assign x_45379 = x_45364 & x_45378;
assign x_45380 = x_14090 & x_14091;
assign x_45381 = x_14089 & x_45380;
assign x_45382 = x_14092 & x_14093;
assign x_45383 = x_14094 & x_14095;
assign x_45384 = x_45382 & x_45383;
assign x_45385 = x_45381 & x_45384;
assign x_45386 = x_14096 & x_14097;
assign x_45387 = x_14098 & x_14099;
assign x_45388 = x_45386 & x_45387;
assign x_45389 = x_14100 & x_14101;
assign x_45390 = x_14102 & x_14103;
assign x_45391 = x_45389 & x_45390;
assign x_45392 = x_45388 & x_45391;
assign x_45393 = x_45385 & x_45392;
assign x_45394 = x_14104 & x_14105;
assign x_45395 = x_14106 & x_14107;
assign x_45396 = x_45394 & x_45395;
assign x_45397 = x_14108 & x_14109;
assign x_45398 = x_14110 & x_14111;
assign x_45399 = x_45397 & x_45398;
assign x_45400 = x_45396 & x_45399;
assign x_45401 = x_14112 & x_14113;
assign x_45402 = x_14114 & x_14115;
assign x_45403 = x_45401 & x_45402;
assign x_45404 = x_14116 & x_14117;
assign x_45405 = x_14118 & x_14119;
assign x_45406 = x_45404 & x_45405;
assign x_45407 = x_45403 & x_45406;
assign x_45408 = x_45400 & x_45407;
assign x_45409 = x_45393 & x_45408;
assign x_45410 = x_45379 & x_45409;
assign x_45411 = x_14121 & x_14122;
assign x_45412 = x_14120 & x_45411;
assign x_45413 = x_14123 & x_14124;
assign x_45414 = x_14125 & x_14126;
assign x_45415 = x_45413 & x_45414;
assign x_45416 = x_45412 & x_45415;
assign x_45417 = x_14127 & x_14128;
assign x_45418 = x_14129 & x_14130;
assign x_45419 = x_45417 & x_45418;
assign x_45420 = x_14131 & x_14132;
assign x_45421 = x_14133 & x_14134;
assign x_45422 = x_45420 & x_45421;
assign x_45423 = x_45419 & x_45422;
assign x_45424 = x_45416 & x_45423;
assign x_45425 = x_14135 & x_14136;
assign x_45426 = x_14137 & x_14138;
assign x_45427 = x_45425 & x_45426;
assign x_45428 = x_14139 & x_14140;
assign x_45429 = x_14141 & x_14142;
assign x_45430 = x_45428 & x_45429;
assign x_45431 = x_45427 & x_45430;
assign x_45432 = x_14143 & x_14144;
assign x_45433 = x_14145 & x_14146;
assign x_45434 = x_45432 & x_45433;
assign x_45435 = x_14147 & x_14148;
assign x_45436 = x_14149 & x_14150;
assign x_45437 = x_45435 & x_45436;
assign x_45438 = x_45434 & x_45437;
assign x_45439 = x_45431 & x_45438;
assign x_45440 = x_45424 & x_45439;
assign x_45441 = x_14152 & x_14153;
assign x_45442 = x_14151 & x_45441;
assign x_45443 = x_14154 & x_14155;
assign x_45444 = x_14156 & x_14157;
assign x_45445 = x_45443 & x_45444;
assign x_45446 = x_45442 & x_45445;
assign x_45447 = x_14158 & x_14159;
assign x_45448 = x_14160 & x_14161;
assign x_45449 = x_45447 & x_45448;
assign x_45450 = x_14162 & x_14163;
assign x_45451 = x_14164 & x_14165;
assign x_45452 = x_45450 & x_45451;
assign x_45453 = x_45449 & x_45452;
assign x_45454 = x_45446 & x_45453;
assign x_45455 = x_14166 & x_14167;
assign x_45456 = x_14168 & x_14169;
assign x_45457 = x_45455 & x_45456;
assign x_45458 = x_14170 & x_14171;
assign x_45459 = x_14172 & x_14173;
assign x_45460 = x_45458 & x_45459;
assign x_45461 = x_45457 & x_45460;
assign x_45462 = x_14174 & x_14175;
assign x_45463 = x_14176 & x_14177;
assign x_45464 = x_45462 & x_45463;
assign x_45465 = x_14178 & x_14179;
assign x_45466 = x_14180 & x_14181;
assign x_45467 = x_45465 & x_45466;
assign x_45468 = x_45464 & x_45467;
assign x_45469 = x_45461 & x_45468;
assign x_45470 = x_45454 & x_45469;
assign x_45471 = x_45440 & x_45470;
assign x_45472 = x_45410 & x_45471;
assign x_45473 = x_45350 & x_45472;
assign x_45474 = x_45229 & x_45473;
assign x_45475 = x_14183 & x_14184;
assign x_45476 = x_14182 & x_45475;
assign x_45477 = x_14185 & x_14186;
assign x_45478 = x_14187 & x_14188;
assign x_45479 = x_45477 & x_45478;
assign x_45480 = x_45476 & x_45479;
assign x_45481 = x_14189 & x_14190;
assign x_45482 = x_14191 & x_14192;
assign x_45483 = x_45481 & x_45482;
assign x_45484 = x_14193 & x_14194;
assign x_45485 = x_14195 & x_14196;
assign x_45486 = x_45484 & x_45485;
assign x_45487 = x_45483 & x_45486;
assign x_45488 = x_45480 & x_45487;
assign x_45489 = x_14198 & x_14199;
assign x_45490 = x_14197 & x_45489;
assign x_45491 = x_14200 & x_14201;
assign x_45492 = x_14202 & x_14203;
assign x_45493 = x_45491 & x_45492;
assign x_45494 = x_45490 & x_45493;
assign x_45495 = x_14204 & x_14205;
assign x_45496 = x_14206 & x_14207;
assign x_45497 = x_45495 & x_45496;
assign x_45498 = x_14208 & x_14209;
assign x_45499 = x_14210 & x_14211;
assign x_45500 = x_45498 & x_45499;
assign x_45501 = x_45497 & x_45500;
assign x_45502 = x_45494 & x_45501;
assign x_45503 = x_45488 & x_45502;
assign x_45504 = x_14213 & x_14214;
assign x_45505 = x_14212 & x_45504;
assign x_45506 = x_14215 & x_14216;
assign x_45507 = x_14217 & x_14218;
assign x_45508 = x_45506 & x_45507;
assign x_45509 = x_45505 & x_45508;
assign x_45510 = x_14219 & x_14220;
assign x_45511 = x_14221 & x_14222;
assign x_45512 = x_45510 & x_45511;
assign x_45513 = x_14223 & x_14224;
assign x_45514 = x_14225 & x_14226;
assign x_45515 = x_45513 & x_45514;
assign x_45516 = x_45512 & x_45515;
assign x_45517 = x_45509 & x_45516;
assign x_45518 = x_14227 & x_14228;
assign x_45519 = x_14229 & x_14230;
assign x_45520 = x_45518 & x_45519;
assign x_45521 = x_14231 & x_14232;
assign x_45522 = x_14233 & x_14234;
assign x_45523 = x_45521 & x_45522;
assign x_45524 = x_45520 & x_45523;
assign x_45525 = x_14235 & x_14236;
assign x_45526 = x_14237 & x_14238;
assign x_45527 = x_45525 & x_45526;
assign x_45528 = x_14239 & x_14240;
assign x_45529 = x_14241 & x_14242;
assign x_45530 = x_45528 & x_45529;
assign x_45531 = x_45527 & x_45530;
assign x_45532 = x_45524 & x_45531;
assign x_45533 = x_45517 & x_45532;
assign x_45534 = x_45503 & x_45533;
assign x_45535 = x_14244 & x_14245;
assign x_45536 = x_14243 & x_45535;
assign x_45537 = x_14246 & x_14247;
assign x_45538 = x_14248 & x_14249;
assign x_45539 = x_45537 & x_45538;
assign x_45540 = x_45536 & x_45539;
assign x_45541 = x_14250 & x_14251;
assign x_45542 = x_14252 & x_14253;
assign x_45543 = x_45541 & x_45542;
assign x_45544 = x_14254 & x_14255;
assign x_45545 = x_14256 & x_14257;
assign x_45546 = x_45544 & x_45545;
assign x_45547 = x_45543 & x_45546;
assign x_45548 = x_45540 & x_45547;
assign x_45549 = x_14259 & x_14260;
assign x_45550 = x_14258 & x_45549;
assign x_45551 = x_14261 & x_14262;
assign x_45552 = x_14263 & x_14264;
assign x_45553 = x_45551 & x_45552;
assign x_45554 = x_45550 & x_45553;
assign x_45555 = x_14265 & x_14266;
assign x_45556 = x_14267 & x_14268;
assign x_45557 = x_45555 & x_45556;
assign x_45558 = x_14269 & x_14270;
assign x_45559 = x_14271 & x_14272;
assign x_45560 = x_45558 & x_45559;
assign x_45561 = x_45557 & x_45560;
assign x_45562 = x_45554 & x_45561;
assign x_45563 = x_45548 & x_45562;
assign x_45564 = x_14274 & x_14275;
assign x_45565 = x_14273 & x_45564;
assign x_45566 = x_14276 & x_14277;
assign x_45567 = x_14278 & x_14279;
assign x_45568 = x_45566 & x_45567;
assign x_45569 = x_45565 & x_45568;
assign x_45570 = x_14280 & x_14281;
assign x_45571 = x_14282 & x_14283;
assign x_45572 = x_45570 & x_45571;
assign x_45573 = x_14284 & x_14285;
assign x_45574 = x_14286 & x_14287;
assign x_45575 = x_45573 & x_45574;
assign x_45576 = x_45572 & x_45575;
assign x_45577 = x_45569 & x_45576;
assign x_45578 = x_14288 & x_14289;
assign x_45579 = x_14290 & x_14291;
assign x_45580 = x_45578 & x_45579;
assign x_45581 = x_14292 & x_14293;
assign x_45582 = x_14294 & x_14295;
assign x_45583 = x_45581 & x_45582;
assign x_45584 = x_45580 & x_45583;
assign x_45585 = x_14296 & x_14297;
assign x_45586 = x_14298 & x_14299;
assign x_45587 = x_45585 & x_45586;
assign x_45588 = x_14300 & x_14301;
assign x_45589 = x_14302 & x_14303;
assign x_45590 = x_45588 & x_45589;
assign x_45591 = x_45587 & x_45590;
assign x_45592 = x_45584 & x_45591;
assign x_45593 = x_45577 & x_45592;
assign x_45594 = x_45563 & x_45593;
assign x_45595 = x_45534 & x_45594;
assign x_45596 = x_14305 & x_14306;
assign x_45597 = x_14304 & x_45596;
assign x_45598 = x_14307 & x_14308;
assign x_45599 = x_14309 & x_14310;
assign x_45600 = x_45598 & x_45599;
assign x_45601 = x_45597 & x_45600;
assign x_45602 = x_14311 & x_14312;
assign x_45603 = x_14313 & x_14314;
assign x_45604 = x_45602 & x_45603;
assign x_45605 = x_14315 & x_14316;
assign x_45606 = x_14317 & x_14318;
assign x_45607 = x_45605 & x_45606;
assign x_45608 = x_45604 & x_45607;
assign x_45609 = x_45601 & x_45608;
assign x_45610 = x_14320 & x_14321;
assign x_45611 = x_14319 & x_45610;
assign x_45612 = x_14322 & x_14323;
assign x_45613 = x_14324 & x_14325;
assign x_45614 = x_45612 & x_45613;
assign x_45615 = x_45611 & x_45614;
assign x_45616 = x_14326 & x_14327;
assign x_45617 = x_14328 & x_14329;
assign x_45618 = x_45616 & x_45617;
assign x_45619 = x_14330 & x_14331;
assign x_45620 = x_14332 & x_14333;
assign x_45621 = x_45619 & x_45620;
assign x_45622 = x_45618 & x_45621;
assign x_45623 = x_45615 & x_45622;
assign x_45624 = x_45609 & x_45623;
assign x_45625 = x_14335 & x_14336;
assign x_45626 = x_14334 & x_45625;
assign x_45627 = x_14337 & x_14338;
assign x_45628 = x_14339 & x_14340;
assign x_45629 = x_45627 & x_45628;
assign x_45630 = x_45626 & x_45629;
assign x_45631 = x_14341 & x_14342;
assign x_45632 = x_14343 & x_14344;
assign x_45633 = x_45631 & x_45632;
assign x_45634 = x_14345 & x_14346;
assign x_45635 = x_14347 & x_14348;
assign x_45636 = x_45634 & x_45635;
assign x_45637 = x_45633 & x_45636;
assign x_45638 = x_45630 & x_45637;
assign x_45639 = x_14349 & x_14350;
assign x_45640 = x_14351 & x_14352;
assign x_45641 = x_45639 & x_45640;
assign x_45642 = x_14353 & x_14354;
assign x_45643 = x_14355 & x_14356;
assign x_45644 = x_45642 & x_45643;
assign x_45645 = x_45641 & x_45644;
assign x_45646 = x_14357 & x_14358;
assign x_45647 = x_14359 & x_14360;
assign x_45648 = x_45646 & x_45647;
assign x_45649 = x_14361 & x_14362;
assign x_45650 = x_14363 & x_14364;
assign x_45651 = x_45649 & x_45650;
assign x_45652 = x_45648 & x_45651;
assign x_45653 = x_45645 & x_45652;
assign x_45654 = x_45638 & x_45653;
assign x_45655 = x_45624 & x_45654;
assign x_45656 = x_14366 & x_14367;
assign x_45657 = x_14365 & x_45656;
assign x_45658 = x_14368 & x_14369;
assign x_45659 = x_14370 & x_14371;
assign x_45660 = x_45658 & x_45659;
assign x_45661 = x_45657 & x_45660;
assign x_45662 = x_14372 & x_14373;
assign x_45663 = x_14374 & x_14375;
assign x_45664 = x_45662 & x_45663;
assign x_45665 = x_14376 & x_14377;
assign x_45666 = x_14378 & x_14379;
assign x_45667 = x_45665 & x_45666;
assign x_45668 = x_45664 & x_45667;
assign x_45669 = x_45661 & x_45668;
assign x_45670 = x_14381 & x_14382;
assign x_45671 = x_14380 & x_45670;
assign x_45672 = x_14383 & x_14384;
assign x_45673 = x_14385 & x_14386;
assign x_45674 = x_45672 & x_45673;
assign x_45675 = x_45671 & x_45674;
assign x_45676 = x_14387 & x_14388;
assign x_45677 = x_14389 & x_14390;
assign x_45678 = x_45676 & x_45677;
assign x_45679 = x_14391 & x_14392;
assign x_45680 = x_14393 & x_14394;
assign x_45681 = x_45679 & x_45680;
assign x_45682 = x_45678 & x_45681;
assign x_45683 = x_45675 & x_45682;
assign x_45684 = x_45669 & x_45683;
assign x_45685 = x_14396 & x_14397;
assign x_45686 = x_14395 & x_45685;
assign x_45687 = x_14398 & x_14399;
assign x_45688 = x_14400 & x_14401;
assign x_45689 = x_45687 & x_45688;
assign x_45690 = x_45686 & x_45689;
assign x_45691 = x_14402 & x_14403;
assign x_45692 = x_14404 & x_14405;
assign x_45693 = x_45691 & x_45692;
assign x_45694 = x_14406 & x_14407;
assign x_45695 = x_14408 & x_14409;
assign x_45696 = x_45694 & x_45695;
assign x_45697 = x_45693 & x_45696;
assign x_45698 = x_45690 & x_45697;
assign x_45699 = x_14410 & x_14411;
assign x_45700 = x_14412 & x_14413;
assign x_45701 = x_45699 & x_45700;
assign x_45702 = x_14414 & x_14415;
assign x_45703 = x_14416 & x_14417;
assign x_45704 = x_45702 & x_45703;
assign x_45705 = x_45701 & x_45704;
assign x_45706 = x_14418 & x_14419;
assign x_45707 = x_14420 & x_14421;
assign x_45708 = x_45706 & x_45707;
assign x_45709 = x_14422 & x_14423;
assign x_45710 = x_14424 & x_14425;
assign x_45711 = x_45709 & x_45710;
assign x_45712 = x_45708 & x_45711;
assign x_45713 = x_45705 & x_45712;
assign x_45714 = x_45698 & x_45713;
assign x_45715 = x_45684 & x_45714;
assign x_45716 = x_45655 & x_45715;
assign x_45717 = x_45595 & x_45716;
assign x_45718 = x_14427 & x_14428;
assign x_45719 = x_14426 & x_45718;
assign x_45720 = x_14429 & x_14430;
assign x_45721 = x_14431 & x_14432;
assign x_45722 = x_45720 & x_45721;
assign x_45723 = x_45719 & x_45722;
assign x_45724 = x_14433 & x_14434;
assign x_45725 = x_14435 & x_14436;
assign x_45726 = x_45724 & x_45725;
assign x_45727 = x_14437 & x_14438;
assign x_45728 = x_14439 & x_14440;
assign x_45729 = x_45727 & x_45728;
assign x_45730 = x_45726 & x_45729;
assign x_45731 = x_45723 & x_45730;
assign x_45732 = x_14442 & x_14443;
assign x_45733 = x_14441 & x_45732;
assign x_45734 = x_14444 & x_14445;
assign x_45735 = x_14446 & x_14447;
assign x_45736 = x_45734 & x_45735;
assign x_45737 = x_45733 & x_45736;
assign x_45738 = x_14448 & x_14449;
assign x_45739 = x_14450 & x_14451;
assign x_45740 = x_45738 & x_45739;
assign x_45741 = x_14452 & x_14453;
assign x_45742 = x_14454 & x_14455;
assign x_45743 = x_45741 & x_45742;
assign x_45744 = x_45740 & x_45743;
assign x_45745 = x_45737 & x_45744;
assign x_45746 = x_45731 & x_45745;
assign x_45747 = x_14457 & x_14458;
assign x_45748 = x_14456 & x_45747;
assign x_45749 = x_14459 & x_14460;
assign x_45750 = x_14461 & x_14462;
assign x_45751 = x_45749 & x_45750;
assign x_45752 = x_45748 & x_45751;
assign x_45753 = x_14463 & x_14464;
assign x_45754 = x_14465 & x_14466;
assign x_45755 = x_45753 & x_45754;
assign x_45756 = x_14467 & x_14468;
assign x_45757 = x_14469 & x_14470;
assign x_45758 = x_45756 & x_45757;
assign x_45759 = x_45755 & x_45758;
assign x_45760 = x_45752 & x_45759;
assign x_45761 = x_14471 & x_14472;
assign x_45762 = x_14473 & x_14474;
assign x_45763 = x_45761 & x_45762;
assign x_45764 = x_14475 & x_14476;
assign x_45765 = x_14477 & x_14478;
assign x_45766 = x_45764 & x_45765;
assign x_45767 = x_45763 & x_45766;
assign x_45768 = x_14479 & x_14480;
assign x_45769 = x_14481 & x_14482;
assign x_45770 = x_45768 & x_45769;
assign x_45771 = x_14483 & x_14484;
assign x_45772 = x_14485 & x_14486;
assign x_45773 = x_45771 & x_45772;
assign x_45774 = x_45770 & x_45773;
assign x_45775 = x_45767 & x_45774;
assign x_45776 = x_45760 & x_45775;
assign x_45777 = x_45746 & x_45776;
assign x_45778 = x_14488 & x_14489;
assign x_45779 = x_14487 & x_45778;
assign x_45780 = x_14490 & x_14491;
assign x_45781 = x_14492 & x_14493;
assign x_45782 = x_45780 & x_45781;
assign x_45783 = x_45779 & x_45782;
assign x_45784 = x_14494 & x_14495;
assign x_45785 = x_14496 & x_14497;
assign x_45786 = x_45784 & x_45785;
assign x_45787 = x_14498 & x_14499;
assign x_45788 = x_14500 & x_14501;
assign x_45789 = x_45787 & x_45788;
assign x_45790 = x_45786 & x_45789;
assign x_45791 = x_45783 & x_45790;
assign x_45792 = x_14503 & x_14504;
assign x_45793 = x_14502 & x_45792;
assign x_45794 = x_14505 & x_14506;
assign x_45795 = x_14507 & x_14508;
assign x_45796 = x_45794 & x_45795;
assign x_45797 = x_45793 & x_45796;
assign x_45798 = x_14509 & x_14510;
assign x_45799 = x_14511 & x_14512;
assign x_45800 = x_45798 & x_45799;
assign x_45801 = x_14513 & x_14514;
assign x_45802 = x_14515 & x_14516;
assign x_45803 = x_45801 & x_45802;
assign x_45804 = x_45800 & x_45803;
assign x_45805 = x_45797 & x_45804;
assign x_45806 = x_45791 & x_45805;
assign x_45807 = x_14518 & x_14519;
assign x_45808 = x_14517 & x_45807;
assign x_45809 = x_14520 & x_14521;
assign x_45810 = x_14522 & x_14523;
assign x_45811 = x_45809 & x_45810;
assign x_45812 = x_45808 & x_45811;
assign x_45813 = x_14524 & x_14525;
assign x_45814 = x_14526 & x_14527;
assign x_45815 = x_45813 & x_45814;
assign x_45816 = x_14528 & x_14529;
assign x_45817 = x_14530 & x_14531;
assign x_45818 = x_45816 & x_45817;
assign x_45819 = x_45815 & x_45818;
assign x_45820 = x_45812 & x_45819;
assign x_45821 = x_14532 & x_14533;
assign x_45822 = x_14534 & x_14535;
assign x_45823 = x_45821 & x_45822;
assign x_45824 = x_14536 & x_14537;
assign x_45825 = x_14538 & x_14539;
assign x_45826 = x_45824 & x_45825;
assign x_45827 = x_45823 & x_45826;
assign x_45828 = x_14540 & x_14541;
assign x_45829 = x_14542 & x_14543;
assign x_45830 = x_45828 & x_45829;
assign x_45831 = x_14544 & x_14545;
assign x_45832 = x_14546 & x_14547;
assign x_45833 = x_45831 & x_45832;
assign x_45834 = x_45830 & x_45833;
assign x_45835 = x_45827 & x_45834;
assign x_45836 = x_45820 & x_45835;
assign x_45837 = x_45806 & x_45836;
assign x_45838 = x_45777 & x_45837;
assign x_45839 = x_14549 & x_14550;
assign x_45840 = x_14548 & x_45839;
assign x_45841 = x_14551 & x_14552;
assign x_45842 = x_14553 & x_14554;
assign x_45843 = x_45841 & x_45842;
assign x_45844 = x_45840 & x_45843;
assign x_45845 = x_14555 & x_14556;
assign x_45846 = x_14557 & x_14558;
assign x_45847 = x_45845 & x_45846;
assign x_45848 = x_14559 & x_14560;
assign x_45849 = x_14561 & x_14562;
assign x_45850 = x_45848 & x_45849;
assign x_45851 = x_45847 & x_45850;
assign x_45852 = x_45844 & x_45851;
assign x_45853 = x_14564 & x_14565;
assign x_45854 = x_14563 & x_45853;
assign x_45855 = x_14566 & x_14567;
assign x_45856 = x_14568 & x_14569;
assign x_45857 = x_45855 & x_45856;
assign x_45858 = x_45854 & x_45857;
assign x_45859 = x_14570 & x_14571;
assign x_45860 = x_14572 & x_14573;
assign x_45861 = x_45859 & x_45860;
assign x_45862 = x_14574 & x_14575;
assign x_45863 = x_14576 & x_14577;
assign x_45864 = x_45862 & x_45863;
assign x_45865 = x_45861 & x_45864;
assign x_45866 = x_45858 & x_45865;
assign x_45867 = x_45852 & x_45866;
assign x_45868 = x_14579 & x_14580;
assign x_45869 = x_14578 & x_45868;
assign x_45870 = x_14581 & x_14582;
assign x_45871 = x_14583 & x_14584;
assign x_45872 = x_45870 & x_45871;
assign x_45873 = x_45869 & x_45872;
assign x_45874 = x_14585 & x_14586;
assign x_45875 = x_14587 & x_14588;
assign x_45876 = x_45874 & x_45875;
assign x_45877 = x_14589 & x_14590;
assign x_45878 = x_14591 & x_14592;
assign x_45879 = x_45877 & x_45878;
assign x_45880 = x_45876 & x_45879;
assign x_45881 = x_45873 & x_45880;
assign x_45882 = x_14593 & x_14594;
assign x_45883 = x_14595 & x_14596;
assign x_45884 = x_45882 & x_45883;
assign x_45885 = x_14597 & x_14598;
assign x_45886 = x_14599 & x_14600;
assign x_45887 = x_45885 & x_45886;
assign x_45888 = x_45884 & x_45887;
assign x_45889 = x_14601 & x_14602;
assign x_45890 = x_14603 & x_14604;
assign x_45891 = x_45889 & x_45890;
assign x_45892 = x_14605 & x_14606;
assign x_45893 = x_14607 & x_14608;
assign x_45894 = x_45892 & x_45893;
assign x_45895 = x_45891 & x_45894;
assign x_45896 = x_45888 & x_45895;
assign x_45897 = x_45881 & x_45896;
assign x_45898 = x_45867 & x_45897;
assign x_45899 = x_14610 & x_14611;
assign x_45900 = x_14609 & x_45899;
assign x_45901 = x_14612 & x_14613;
assign x_45902 = x_14614 & x_14615;
assign x_45903 = x_45901 & x_45902;
assign x_45904 = x_45900 & x_45903;
assign x_45905 = x_14616 & x_14617;
assign x_45906 = x_14618 & x_14619;
assign x_45907 = x_45905 & x_45906;
assign x_45908 = x_14620 & x_14621;
assign x_45909 = x_14622 & x_14623;
assign x_45910 = x_45908 & x_45909;
assign x_45911 = x_45907 & x_45910;
assign x_45912 = x_45904 & x_45911;
assign x_45913 = x_14624 & x_14625;
assign x_45914 = x_14626 & x_14627;
assign x_45915 = x_45913 & x_45914;
assign x_45916 = x_14628 & x_14629;
assign x_45917 = x_14630 & x_14631;
assign x_45918 = x_45916 & x_45917;
assign x_45919 = x_45915 & x_45918;
assign x_45920 = x_14632 & x_14633;
assign x_45921 = x_14634 & x_14635;
assign x_45922 = x_45920 & x_45921;
assign x_45923 = x_14636 & x_14637;
assign x_45924 = x_14638 & x_14639;
assign x_45925 = x_45923 & x_45924;
assign x_45926 = x_45922 & x_45925;
assign x_45927 = x_45919 & x_45926;
assign x_45928 = x_45912 & x_45927;
assign x_45929 = x_14641 & x_14642;
assign x_45930 = x_14640 & x_45929;
assign x_45931 = x_14643 & x_14644;
assign x_45932 = x_14645 & x_14646;
assign x_45933 = x_45931 & x_45932;
assign x_45934 = x_45930 & x_45933;
assign x_45935 = x_14647 & x_14648;
assign x_45936 = x_14649 & x_14650;
assign x_45937 = x_45935 & x_45936;
assign x_45938 = x_14651 & x_14652;
assign x_45939 = x_14653 & x_14654;
assign x_45940 = x_45938 & x_45939;
assign x_45941 = x_45937 & x_45940;
assign x_45942 = x_45934 & x_45941;
assign x_45943 = x_14655 & x_14656;
assign x_45944 = x_14657 & x_14658;
assign x_45945 = x_45943 & x_45944;
assign x_45946 = x_14659 & x_14660;
assign x_45947 = x_14661 & x_14662;
assign x_45948 = x_45946 & x_45947;
assign x_45949 = x_45945 & x_45948;
assign x_45950 = x_14663 & x_14664;
assign x_45951 = x_14665 & x_14666;
assign x_45952 = x_45950 & x_45951;
assign x_45953 = x_14667 & x_14668;
assign x_45954 = x_14669 & x_14670;
assign x_45955 = x_45953 & x_45954;
assign x_45956 = x_45952 & x_45955;
assign x_45957 = x_45949 & x_45956;
assign x_45958 = x_45942 & x_45957;
assign x_45959 = x_45928 & x_45958;
assign x_45960 = x_45898 & x_45959;
assign x_45961 = x_45838 & x_45960;
assign x_45962 = x_45717 & x_45961;
assign x_45963 = x_45474 & x_45962;
assign x_45964 = x_14672 & x_14673;
assign x_45965 = x_14671 & x_45964;
assign x_45966 = x_14674 & x_14675;
assign x_45967 = x_14676 & x_14677;
assign x_45968 = x_45966 & x_45967;
assign x_45969 = x_45965 & x_45968;
assign x_45970 = x_14678 & x_14679;
assign x_45971 = x_14680 & x_14681;
assign x_45972 = x_45970 & x_45971;
assign x_45973 = x_14682 & x_14683;
assign x_45974 = x_14684 & x_14685;
assign x_45975 = x_45973 & x_45974;
assign x_45976 = x_45972 & x_45975;
assign x_45977 = x_45969 & x_45976;
assign x_45978 = x_14687 & x_14688;
assign x_45979 = x_14686 & x_45978;
assign x_45980 = x_14689 & x_14690;
assign x_45981 = x_14691 & x_14692;
assign x_45982 = x_45980 & x_45981;
assign x_45983 = x_45979 & x_45982;
assign x_45984 = x_14693 & x_14694;
assign x_45985 = x_14695 & x_14696;
assign x_45986 = x_45984 & x_45985;
assign x_45987 = x_14697 & x_14698;
assign x_45988 = x_14699 & x_14700;
assign x_45989 = x_45987 & x_45988;
assign x_45990 = x_45986 & x_45989;
assign x_45991 = x_45983 & x_45990;
assign x_45992 = x_45977 & x_45991;
assign x_45993 = x_14702 & x_14703;
assign x_45994 = x_14701 & x_45993;
assign x_45995 = x_14704 & x_14705;
assign x_45996 = x_14706 & x_14707;
assign x_45997 = x_45995 & x_45996;
assign x_45998 = x_45994 & x_45997;
assign x_45999 = x_14708 & x_14709;
assign x_46000 = x_14710 & x_14711;
assign x_46001 = x_45999 & x_46000;
assign x_46002 = x_14712 & x_14713;
assign x_46003 = x_14714 & x_14715;
assign x_46004 = x_46002 & x_46003;
assign x_46005 = x_46001 & x_46004;
assign x_46006 = x_45998 & x_46005;
assign x_46007 = x_14716 & x_14717;
assign x_46008 = x_14718 & x_14719;
assign x_46009 = x_46007 & x_46008;
assign x_46010 = x_14720 & x_14721;
assign x_46011 = x_14722 & x_14723;
assign x_46012 = x_46010 & x_46011;
assign x_46013 = x_46009 & x_46012;
assign x_46014 = x_14724 & x_14725;
assign x_46015 = x_14726 & x_14727;
assign x_46016 = x_46014 & x_46015;
assign x_46017 = x_14728 & x_14729;
assign x_46018 = x_14730 & x_14731;
assign x_46019 = x_46017 & x_46018;
assign x_46020 = x_46016 & x_46019;
assign x_46021 = x_46013 & x_46020;
assign x_46022 = x_46006 & x_46021;
assign x_46023 = x_45992 & x_46022;
assign x_46024 = x_14733 & x_14734;
assign x_46025 = x_14732 & x_46024;
assign x_46026 = x_14735 & x_14736;
assign x_46027 = x_14737 & x_14738;
assign x_46028 = x_46026 & x_46027;
assign x_46029 = x_46025 & x_46028;
assign x_46030 = x_14739 & x_14740;
assign x_46031 = x_14741 & x_14742;
assign x_46032 = x_46030 & x_46031;
assign x_46033 = x_14743 & x_14744;
assign x_46034 = x_14745 & x_14746;
assign x_46035 = x_46033 & x_46034;
assign x_46036 = x_46032 & x_46035;
assign x_46037 = x_46029 & x_46036;
assign x_46038 = x_14748 & x_14749;
assign x_46039 = x_14747 & x_46038;
assign x_46040 = x_14750 & x_14751;
assign x_46041 = x_14752 & x_14753;
assign x_46042 = x_46040 & x_46041;
assign x_46043 = x_46039 & x_46042;
assign x_46044 = x_14754 & x_14755;
assign x_46045 = x_14756 & x_14757;
assign x_46046 = x_46044 & x_46045;
assign x_46047 = x_14758 & x_14759;
assign x_46048 = x_14760 & x_14761;
assign x_46049 = x_46047 & x_46048;
assign x_46050 = x_46046 & x_46049;
assign x_46051 = x_46043 & x_46050;
assign x_46052 = x_46037 & x_46051;
assign x_46053 = x_14763 & x_14764;
assign x_46054 = x_14762 & x_46053;
assign x_46055 = x_14765 & x_14766;
assign x_46056 = x_14767 & x_14768;
assign x_46057 = x_46055 & x_46056;
assign x_46058 = x_46054 & x_46057;
assign x_46059 = x_14769 & x_14770;
assign x_46060 = x_14771 & x_14772;
assign x_46061 = x_46059 & x_46060;
assign x_46062 = x_14773 & x_14774;
assign x_46063 = x_14775 & x_14776;
assign x_46064 = x_46062 & x_46063;
assign x_46065 = x_46061 & x_46064;
assign x_46066 = x_46058 & x_46065;
assign x_46067 = x_14777 & x_14778;
assign x_46068 = x_14779 & x_14780;
assign x_46069 = x_46067 & x_46068;
assign x_46070 = x_14781 & x_14782;
assign x_46071 = x_14783 & x_14784;
assign x_46072 = x_46070 & x_46071;
assign x_46073 = x_46069 & x_46072;
assign x_46074 = x_14785 & x_14786;
assign x_46075 = x_14787 & x_14788;
assign x_46076 = x_46074 & x_46075;
assign x_46077 = x_14789 & x_14790;
assign x_46078 = x_14791 & x_14792;
assign x_46079 = x_46077 & x_46078;
assign x_46080 = x_46076 & x_46079;
assign x_46081 = x_46073 & x_46080;
assign x_46082 = x_46066 & x_46081;
assign x_46083 = x_46052 & x_46082;
assign x_46084 = x_46023 & x_46083;
assign x_46085 = x_14794 & x_14795;
assign x_46086 = x_14793 & x_46085;
assign x_46087 = x_14796 & x_14797;
assign x_46088 = x_14798 & x_14799;
assign x_46089 = x_46087 & x_46088;
assign x_46090 = x_46086 & x_46089;
assign x_46091 = x_14800 & x_14801;
assign x_46092 = x_14802 & x_14803;
assign x_46093 = x_46091 & x_46092;
assign x_46094 = x_14804 & x_14805;
assign x_46095 = x_14806 & x_14807;
assign x_46096 = x_46094 & x_46095;
assign x_46097 = x_46093 & x_46096;
assign x_46098 = x_46090 & x_46097;
assign x_46099 = x_14809 & x_14810;
assign x_46100 = x_14808 & x_46099;
assign x_46101 = x_14811 & x_14812;
assign x_46102 = x_14813 & x_14814;
assign x_46103 = x_46101 & x_46102;
assign x_46104 = x_46100 & x_46103;
assign x_46105 = x_14815 & x_14816;
assign x_46106 = x_14817 & x_14818;
assign x_46107 = x_46105 & x_46106;
assign x_46108 = x_14819 & x_14820;
assign x_46109 = x_14821 & x_14822;
assign x_46110 = x_46108 & x_46109;
assign x_46111 = x_46107 & x_46110;
assign x_46112 = x_46104 & x_46111;
assign x_46113 = x_46098 & x_46112;
assign x_46114 = x_14824 & x_14825;
assign x_46115 = x_14823 & x_46114;
assign x_46116 = x_14826 & x_14827;
assign x_46117 = x_14828 & x_14829;
assign x_46118 = x_46116 & x_46117;
assign x_46119 = x_46115 & x_46118;
assign x_46120 = x_14830 & x_14831;
assign x_46121 = x_14832 & x_14833;
assign x_46122 = x_46120 & x_46121;
assign x_46123 = x_14834 & x_14835;
assign x_46124 = x_14836 & x_14837;
assign x_46125 = x_46123 & x_46124;
assign x_46126 = x_46122 & x_46125;
assign x_46127 = x_46119 & x_46126;
assign x_46128 = x_14838 & x_14839;
assign x_46129 = x_14840 & x_14841;
assign x_46130 = x_46128 & x_46129;
assign x_46131 = x_14842 & x_14843;
assign x_46132 = x_14844 & x_14845;
assign x_46133 = x_46131 & x_46132;
assign x_46134 = x_46130 & x_46133;
assign x_46135 = x_14846 & x_14847;
assign x_46136 = x_14848 & x_14849;
assign x_46137 = x_46135 & x_46136;
assign x_46138 = x_14850 & x_14851;
assign x_46139 = x_14852 & x_14853;
assign x_46140 = x_46138 & x_46139;
assign x_46141 = x_46137 & x_46140;
assign x_46142 = x_46134 & x_46141;
assign x_46143 = x_46127 & x_46142;
assign x_46144 = x_46113 & x_46143;
assign x_46145 = x_14855 & x_14856;
assign x_46146 = x_14854 & x_46145;
assign x_46147 = x_14857 & x_14858;
assign x_46148 = x_14859 & x_14860;
assign x_46149 = x_46147 & x_46148;
assign x_46150 = x_46146 & x_46149;
assign x_46151 = x_14861 & x_14862;
assign x_46152 = x_14863 & x_14864;
assign x_46153 = x_46151 & x_46152;
assign x_46154 = x_14865 & x_14866;
assign x_46155 = x_14867 & x_14868;
assign x_46156 = x_46154 & x_46155;
assign x_46157 = x_46153 & x_46156;
assign x_46158 = x_46150 & x_46157;
assign x_46159 = x_14870 & x_14871;
assign x_46160 = x_14869 & x_46159;
assign x_46161 = x_14872 & x_14873;
assign x_46162 = x_14874 & x_14875;
assign x_46163 = x_46161 & x_46162;
assign x_46164 = x_46160 & x_46163;
assign x_46165 = x_14876 & x_14877;
assign x_46166 = x_14878 & x_14879;
assign x_46167 = x_46165 & x_46166;
assign x_46168 = x_14880 & x_14881;
assign x_46169 = x_14882 & x_14883;
assign x_46170 = x_46168 & x_46169;
assign x_46171 = x_46167 & x_46170;
assign x_46172 = x_46164 & x_46171;
assign x_46173 = x_46158 & x_46172;
assign x_46174 = x_14885 & x_14886;
assign x_46175 = x_14884 & x_46174;
assign x_46176 = x_14887 & x_14888;
assign x_46177 = x_14889 & x_14890;
assign x_46178 = x_46176 & x_46177;
assign x_46179 = x_46175 & x_46178;
assign x_46180 = x_14891 & x_14892;
assign x_46181 = x_14893 & x_14894;
assign x_46182 = x_46180 & x_46181;
assign x_46183 = x_14895 & x_14896;
assign x_46184 = x_14897 & x_14898;
assign x_46185 = x_46183 & x_46184;
assign x_46186 = x_46182 & x_46185;
assign x_46187 = x_46179 & x_46186;
assign x_46188 = x_14899 & x_14900;
assign x_46189 = x_14901 & x_14902;
assign x_46190 = x_46188 & x_46189;
assign x_46191 = x_14903 & x_14904;
assign x_46192 = x_14905 & x_14906;
assign x_46193 = x_46191 & x_46192;
assign x_46194 = x_46190 & x_46193;
assign x_46195 = x_14907 & x_14908;
assign x_46196 = x_14909 & x_14910;
assign x_46197 = x_46195 & x_46196;
assign x_46198 = x_14911 & x_14912;
assign x_46199 = x_14913 & x_14914;
assign x_46200 = x_46198 & x_46199;
assign x_46201 = x_46197 & x_46200;
assign x_46202 = x_46194 & x_46201;
assign x_46203 = x_46187 & x_46202;
assign x_46204 = x_46173 & x_46203;
assign x_46205 = x_46144 & x_46204;
assign x_46206 = x_46084 & x_46205;
assign x_46207 = x_14916 & x_14917;
assign x_46208 = x_14915 & x_46207;
assign x_46209 = x_14918 & x_14919;
assign x_46210 = x_14920 & x_14921;
assign x_46211 = x_46209 & x_46210;
assign x_46212 = x_46208 & x_46211;
assign x_46213 = x_14922 & x_14923;
assign x_46214 = x_14924 & x_14925;
assign x_46215 = x_46213 & x_46214;
assign x_46216 = x_14926 & x_14927;
assign x_46217 = x_14928 & x_14929;
assign x_46218 = x_46216 & x_46217;
assign x_46219 = x_46215 & x_46218;
assign x_46220 = x_46212 & x_46219;
assign x_46221 = x_14931 & x_14932;
assign x_46222 = x_14930 & x_46221;
assign x_46223 = x_14933 & x_14934;
assign x_46224 = x_14935 & x_14936;
assign x_46225 = x_46223 & x_46224;
assign x_46226 = x_46222 & x_46225;
assign x_46227 = x_14937 & x_14938;
assign x_46228 = x_14939 & x_14940;
assign x_46229 = x_46227 & x_46228;
assign x_46230 = x_14941 & x_14942;
assign x_46231 = x_14943 & x_14944;
assign x_46232 = x_46230 & x_46231;
assign x_46233 = x_46229 & x_46232;
assign x_46234 = x_46226 & x_46233;
assign x_46235 = x_46220 & x_46234;
assign x_46236 = x_14946 & x_14947;
assign x_46237 = x_14945 & x_46236;
assign x_46238 = x_14948 & x_14949;
assign x_46239 = x_14950 & x_14951;
assign x_46240 = x_46238 & x_46239;
assign x_46241 = x_46237 & x_46240;
assign x_46242 = x_14952 & x_14953;
assign x_46243 = x_14954 & x_14955;
assign x_46244 = x_46242 & x_46243;
assign x_46245 = x_14956 & x_14957;
assign x_46246 = x_14958 & x_14959;
assign x_46247 = x_46245 & x_46246;
assign x_46248 = x_46244 & x_46247;
assign x_46249 = x_46241 & x_46248;
assign x_46250 = x_14960 & x_14961;
assign x_46251 = x_14962 & x_14963;
assign x_46252 = x_46250 & x_46251;
assign x_46253 = x_14964 & x_14965;
assign x_46254 = x_14966 & x_14967;
assign x_46255 = x_46253 & x_46254;
assign x_46256 = x_46252 & x_46255;
assign x_46257 = x_14968 & x_14969;
assign x_46258 = x_14970 & x_14971;
assign x_46259 = x_46257 & x_46258;
assign x_46260 = x_14972 & x_14973;
assign x_46261 = x_14974 & x_14975;
assign x_46262 = x_46260 & x_46261;
assign x_46263 = x_46259 & x_46262;
assign x_46264 = x_46256 & x_46263;
assign x_46265 = x_46249 & x_46264;
assign x_46266 = x_46235 & x_46265;
assign x_46267 = x_14977 & x_14978;
assign x_46268 = x_14976 & x_46267;
assign x_46269 = x_14979 & x_14980;
assign x_46270 = x_14981 & x_14982;
assign x_46271 = x_46269 & x_46270;
assign x_46272 = x_46268 & x_46271;
assign x_46273 = x_14983 & x_14984;
assign x_46274 = x_14985 & x_14986;
assign x_46275 = x_46273 & x_46274;
assign x_46276 = x_14987 & x_14988;
assign x_46277 = x_14989 & x_14990;
assign x_46278 = x_46276 & x_46277;
assign x_46279 = x_46275 & x_46278;
assign x_46280 = x_46272 & x_46279;
assign x_46281 = x_14992 & x_14993;
assign x_46282 = x_14991 & x_46281;
assign x_46283 = x_14994 & x_14995;
assign x_46284 = x_14996 & x_14997;
assign x_46285 = x_46283 & x_46284;
assign x_46286 = x_46282 & x_46285;
assign x_46287 = x_14998 & x_14999;
assign x_46288 = x_15000 & x_15001;
assign x_46289 = x_46287 & x_46288;
assign x_46290 = x_15002 & x_15003;
assign x_46291 = x_15004 & x_15005;
assign x_46292 = x_46290 & x_46291;
assign x_46293 = x_46289 & x_46292;
assign x_46294 = x_46286 & x_46293;
assign x_46295 = x_46280 & x_46294;
assign x_46296 = x_15007 & x_15008;
assign x_46297 = x_15006 & x_46296;
assign x_46298 = x_15009 & x_15010;
assign x_46299 = x_15011 & x_15012;
assign x_46300 = x_46298 & x_46299;
assign x_46301 = x_46297 & x_46300;
assign x_46302 = x_15013 & x_15014;
assign x_46303 = x_15015 & x_15016;
assign x_46304 = x_46302 & x_46303;
assign x_46305 = x_15017 & x_15018;
assign x_46306 = x_15019 & x_15020;
assign x_46307 = x_46305 & x_46306;
assign x_46308 = x_46304 & x_46307;
assign x_46309 = x_46301 & x_46308;
assign x_46310 = x_15021 & x_15022;
assign x_46311 = x_15023 & x_15024;
assign x_46312 = x_46310 & x_46311;
assign x_46313 = x_15025 & x_15026;
assign x_46314 = x_15027 & x_15028;
assign x_46315 = x_46313 & x_46314;
assign x_46316 = x_46312 & x_46315;
assign x_46317 = x_15029 & x_15030;
assign x_46318 = x_15031 & x_15032;
assign x_46319 = x_46317 & x_46318;
assign x_46320 = x_15033 & x_15034;
assign x_46321 = x_15035 & x_15036;
assign x_46322 = x_46320 & x_46321;
assign x_46323 = x_46319 & x_46322;
assign x_46324 = x_46316 & x_46323;
assign x_46325 = x_46309 & x_46324;
assign x_46326 = x_46295 & x_46325;
assign x_46327 = x_46266 & x_46326;
assign x_46328 = x_15038 & x_15039;
assign x_46329 = x_15037 & x_46328;
assign x_46330 = x_15040 & x_15041;
assign x_46331 = x_15042 & x_15043;
assign x_46332 = x_46330 & x_46331;
assign x_46333 = x_46329 & x_46332;
assign x_46334 = x_15044 & x_15045;
assign x_46335 = x_15046 & x_15047;
assign x_46336 = x_46334 & x_46335;
assign x_46337 = x_15048 & x_15049;
assign x_46338 = x_15050 & x_15051;
assign x_46339 = x_46337 & x_46338;
assign x_46340 = x_46336 & x_46339;
assign x_46341 = x_46333 & x_46340;
assign x_46342 = x_15053 & x_15054;
assign x_46343 = x_15052 & x_46342;
assign x_46344 = x_15055 & x_15056;
assign x_46345 = x_15057 & x_15058;
assign x_46346 = x_46344 & x_46345;
assign x_46347 = x_46343 & x_46346;
assign x_46348 = x_15059 & x_15060;
assign x_46349 = x_15061 & x_15062;
assign x_46350 = x_46348 & x_46349;
assign x_46351 = x_15063 & x_15064;
assign x_46352 = x_15065 & x_15066;
assign x_46353 = x_46351 & x_46352;
assign x_46354 = x_46350 & x_46353;
assign x_46355 = x_46347 & x_46354;
assign x_46356 = x_46341 & x_46355;
assign x_46357 = x_15068 & x_15069;
assign x_46358 = x_15067 & x_46357;
assign x_46359 = x_15070 & x_15071;
assign x_46360 = x_15072 & x_15073;
assign x_46361 = x_46359 & x_46360;
assign x_46362 = x_46358 & x_46361;
assign x_46363 = x_15074 & x_15075;
assign x_46364 = x_15076 & x_15077;
assign x_46365 = x_46363 & x_46364;
assign x_46366 = x_15078 & x_15079;
assign x_46367 = x_15080 & x_15081;
assign x_46368 = x_46366 & x_46367;
assign x_46369 = x_46365 & x_46368;
assign x_46370 = x_46362 & x_46369;
assign x_46371 = x_15082 & x_15083;
assign x_46372 = x_15084 & x_15085;
assign x_46373 = x_46371 & x_46372;
assign x_46374 = x_15086 & x_15087;
assign x_46375 = x_15088 & x_15089;
assign x_46376 = x_46374 & x_46375;
assign x_46377 = x_46373 & x_46376;
assign x_46378 = x_15090 & x_15091;
assign x_46379 = x_15092 & x_15093;
assign x_46380 = x_46378 & x_46379;
assign x_46381 = x_15094 & x_15095;
assign x_46382 = x_15096 & x_15097;
assign x_46383 = x_46381 & x_46382;
assign x_46384 = x_46380 & x_46383;
assign x_46385 = x_46377 & x_46384;
assign x_46386 = x_46370 & x_46385;
assign x_46387 = x_46356 & x_46386;
assign x_46388 = x_15099 & x_15100;
assign x_46389 = x_15098 & x_46388;
assign x_46390 = x_15101 & x_15102;
assign x_46391 = x_15103 & x_15104;
assign x_46392 = x_46390 & x_46391;
assign x_46393 = x_46389 & x_46392;
assign x_46394 = x_15105 & x_15106;
assign x_46395 = x_15107 & x_15108;
assign x_46396 = x_46394 & x_46395;
assign x_46397 = x_15109 & x_15110;
assign x_46398 = x_15111 & x_15112;
assign x_46399 = x_46397 & x_46398;
assign x_46400 = x_46396 & x_46399;
assign x_46401 = x_46393 & x_46400;
assign x_46402 = x_15113 & x_15114;
assign x_46403 = x_15115 & x_15116;
assign x_46404 = x_46402 & x_46403;
assign x_46405 = x_15117 & x_15118;
assign x_46406 = x_15119 & x_15120;
assign x_46407 = x_46405 & x_46406;
assign x_46408 = x_46404 & x_46407;
assign x_46409 = x_15121 & x_15122;
assign x_46410 = x_15123 & x_15124;
assign x_46411 = x_46409 & x_46410;
assign x_46412 = x_15125 & x_15126;
assign x_46413 = x_15127 & x_15128;
assign x_46414 = x_46412 & x_46413;
assign x_46415 = x_46411 & x_46414;
assign x_46416 = x_46408 & x_46415;
assign x_46417 = x_46401 & x_46416;
assign x_46418 = x_15130 & x_15131;
assign x_46419 = x_15129 & x_46418;
assign x_46420 = x_15132 & x_15133;
assign x_46421 = x_15134 & x_15135;
assign x_46422 = x_46420 & x_46421;
assign x_46423 = x_46419 & x_46422;
assign x_46424 = x_15136 & x_15137;
assign x_46425 = x_15138 & x_15139;
assign x_46426 = x_46424 & x_46425;
assign x_46427 = x_15140 & x_15141;
assign x_46428 = x_15142 & x_15143;
assign x_46429 = x_46427 & x_46428;
assign x_46430 = x_46426 & x_46429;
assign x_46431 = x_46423 & x_46430;
assign x_46432 = x_15144 & x_15145;
assign x_46433 = x_15146 & x_15147;
assign x_46434 = x_46432 & x_46433;
assign x_46435 = x_15148 & x_15149;
assign x_46436 = x_15150 & x_15151;
assign x_46437 = x_46435 & x_46436;
assign x_46438 = x_46434 & x_46437;
assign x_46439 = x_15152 & x_15153;
assign x_46440 = x_15154 & x_15155;
assign x_46441 = x_46439 & x_46440;
assign x_46442 = x_15156 & x_15157;
assign x_46443 = x_15158 & x_15159;
assign x_46444 = x_46442 & x_46443;
assign x_46445 = x_46441 & x_46444;
assign x_46446 = x_46438 & x_46445;
assign x_46447 = x_46431 & x_46446;
assign x_46448 = x_46417 & x_46447;
assign x_46449 = x_46387 & x_46448;
assign x_46450 = x_46327 & x_46449;
assign x_46451 = x_46206 & x_46450;
assign x_46452 = x_15161 & x_15162;
assign x_46453 = x_15160 & x_46452;
assign x_46454 = x_15163 & x_15164;
assign x_46455 = x_15165 & x_15166;
assign x_46456 = x_46454 & x_46455;
assign x_46457 = x_46453 & x_46456;
assign x_46458 = x_15167 & x_15168;
assign x_46459 = x_15169 & x_15170;
assign x_46460 = x_46458 & x_46459;
assign x_46461 = x_15171 & x_15172;
assign x_46462 = x_15173 & x_15174;
assign x_46463 = x_46461 & x_46462;
assign x_46464 = x_46460 & x_46463;
assign x_46465 = x_46457 & x_46464;
assign x_46466 = x_15176 & x_15177;
assign x_46467 = x_15175 & x_46466;
assign x_46468 = x_15178 & x_15179;
assign x_46469 = x_15180 & x_15181;
assign x_46470 = x_46468 & x_46469;
assign x_46471 = x_46467 & x_46470;
assign x_46472 = x_15182 & x_15183;
assign x_46473 = x_15184 & x_15185;
assign x_46474 = x_46472 & x_46473;
assign x_46475 = x_15186 & x_15187;
assign x_46476 = x_15188 & x_15189;
assign x_46477 = x_46475 & x_46476;
assign x_46478 = x_46474 & x_46477;
assign x_46479 = x_46471 & x_46478;
assign x_46480 = x_46465 & x_46479;
assign x_46481 = x_15191 & x_15192;
assign x_46482 = x_15190 & x_46481;
assign x_46483 = x_15193 & x_15194;
assign x_46484 = x_15195 & x_15196;
assign x_46485 = x_46483 & x_46484;
assign x_46486 = x_46482 & x_46485;
assign x_46487 = x_15197 & x_15198;
assign x_46488 = x_15199 & x_15200;
assign x_46489 = x_46487 & x_46488;
assign x_46490 = x_15201 & x_15202;
assign x_46491 = x_15203 & x_15204;
assign x_46492 = x_46490 & x_46491;
assign x_46493 = x_46489 & x_46492;
assign x_46494 = x_46486 & x_46493;
assign x_46495 = x_15205 & x_15206;
assign x_46496 = x_15207 & x_15208;
assign x_46497 = x_46495 & x_46496;
assign x_46498 = x_15209 & x_15210;
assign x_46499 = x_15211 & x_15212;
assign x_46500 = x_46498 & x_46499;
assign x_46501 = x_46497 & x_46500;
assign x_46502 = x_15213 & x_15214;
assign x_46503 = x_15215 & x_15216;
assign x_46504 = x_46502 & x_46503;
assign x_46505 = x_15217 & x_15218;
assign x_46506 = x_15219 & x_15220;
assign x_46507 = x_46505 & x_46506;
assign x_46508 = x_46504 & x_46507;
assign x_46509 = x_46501 & x_46508;
assign x_46510 = x_46494 & x_46509;
assign x_46511 = x_46480 & x_46510;
assign x_46512 = x_15222 & x_15223;
assign x_46513 = x_15221 & x_46512;
assign x_46514 = x_15224 & x_15225;
assign x_46515 = x_15226 & x_15227;
assign x_46516 = x_46514 & x_46515;
assign x_46517 = x_46513 & x_46516;
assign x_46518 = x_15228 & x_15229;
assign x_46519 = x_15230 & x_15231;
assign x_46520 = x_46518 & x_46519;
assign x_46521 = x_15232 & x_15233;
assign x_46522 = x_15234 & x_15235;
assign x_46523 = x_46521 & x_46522;
assign x_46524 = x_46520 & x_46523;
assign x_46525 = x_46517 & x_46524;
assign x_46526 = x_15237 & x_15238;
assign x_46527 = x_15236 & x_46526;
assign x_46528 = x_15239 & x_15240;
assign x_46529 = x_15241 & x_15242;
assign x_46530 = x_46528 & x_46529;
assign x_46531 = x_46527 & x_46530;
assign x_46532 = x_15243 & x_15244;
assign x_46533 = x_15245 & x_15246;
assign x_46534 = x_46532 & x_46533;
assign x_46535 = x_15247 & x_15248;
assign x_46536 = x_15249 & x_15250;
assign x_46537 = x_46535 & x_46536;
assign x_46538 = x_46534 & x_46537;
assign x_46539 = x_46531 & x_46538;
assign x_46540 = x_46525 & x_46539;
assign x_46541 = x_15252 & x_15253;
assign x_46542 = x_15251 & x_46541;
assign x_46543 = x_15254 & x_15255;
assign x_46544 = x_15256 & x_15257;
assign x_46545 = x_46543 & x_46544;
assign x_46546 = x_46542 & x_46545;
assign x_46547 = x_15258 & x_15259;
assign x_46548 = x_15260 & x_15261;
assign x_46549 = x_46547 & x_46548;
assign x_46550 = x_15262 & x_15263;
assign x_46551 = x_15264 & x_15265;
assign x_46552 = x_46550 & x_46551;
assign x_46553 = x_46549 & x_46552;
assign x_46554 = x_46546 & x_46553;
assign x_46555 = x_15266 & x_15267;
assign x_46556 = x_15268 & x_15269;
assign x_46557 = x_46555 & x_46556;
assign x_46558 = x_15270 & x_15271;
assign x_46559 = x_15272 & x_15273;
assign x_46560 = x_46558 & x_46559;
assign x_46561 = x_46557 & x_46560;
assign x_46562 = x_15274 & x_15275;
assign x_46563 = x_15276 & x_15277;
assign x_46564 = x_46562 & x_46563;
assign x_46565 = x_15278 & x_15279;
assign x_46566 = x_15280 & x_15281;
assign x_46567 = x_46565 & x_46566;
assign x_46568 = x_46564 & x_46567;
assign x_46569 = x_46561 & x_46568;
assign x_46570 = x_46554 & x_46569;
assign x_46571 = x_46540 & x_46570;
assign x_46572 = x_46511 & x_46571;
assign x_46573 = x_15283 & x_15284;
assign x_46574 = x_15282 & x_46573;
assign x_46575 = x_15285 & x_15286;
assign x_46576 = x_15287 & x_15288;
assign x_46577 = x_46575 & x_46576;
assign x_46578 = x_46574 & x_46577;
assign x_46579 = x_15289 & x_15290;
assign x_46580 = x_15291 & x_15292;
assign x_46581 = x_46579 & x_46580;
assign x_46582 = x_15293 & x_15294;
assign x_46583 = x_15295 & x_15296;
assign x_46584 = x_46582 & x_46583;
assign x_46585 = x_46581 & x_46584;
assign x_46586 = x_46578 & x_46585;
assign x_46587 = x_15298 & x_15299;
assign x_46588 = x_15297 & x_46587;
assign x_46589 = x_15300 & x_15301;
assign x_46590 = x_15302 & x_15303;
assign x_46591 = x_46589 & x_46590;
assign x_46592 = x_46588 & x_46591;
assign x_46593 = x_15304 & x_15305;
assign x_46594 = x_15306 & x_15307;
assign x_46595 = x_46593 & x_46594;
assign x_46596 = x_15308 & x_15309;
assign x_46597 = x_15310 & x_15311;
assign x_46598 = x_46596 & x_46597;
assign x_46599 = x_46595 & x_46598;
assign x_46600 = x_46592 & x_46599;
assign x_46601 = x_46586 & x_46600;
assign x_46602 = x_15313 & x_15314;
assign x_46603 = x_15312 & x_46602;
assign x_46604 = x_15315 & x_15316;
assign x_46605 = x_15317 & x_15318;
assign x_46606 = x_46604 & x_46605;
assign x_46607 = x_46603 & x_46606;
assign x_46608 = x_15319 & x_15320;
assign x_46609 = x_15321 & x_15322;
assign x_46610 = x_46608 & x_46609;
assign x_46611 = x_15323 & x_15324;
assign x_46612 = x_15325 & x_15326;
assign x_46613 = x_46611 & x_46612;
assign x_46614 = x_46610 & x_46613;
assign x_46615 = x_46607 & x_46614;
assign x_46616 = x_15327 & x_15328;
assign x_46617 = x_15329 & x_15330;
assign x_46618 = x_46616 & x_46617;
assign x_46619 = x_15331 & x_15332;
assign x_46620 = x_15333 & x_15334;
assign x_46621 = x_46619 & x_46620;
assign x_46622 = x_46618 & x_46621;
assign x_46623 = x_15335 & x_15336;
assign x_46624 = x_15337 & x_15338;
assign x_46625 = x_46623 & x_46624;
assign x_46626 = x_15339 & x_15340;
assign x_46627 = x_15341 & x_15342;
assign x_46628 = x_46626 & x_46627;
assign x_46629 = x_46625 & x_46628;
assign x_46630 = x_46622 & x_46629;
assign x_46631 = x_46615 & x_46630;
assign x_46632 = x_46601 & x_46631;
assign x_46633 = x_15344 & x_15345;
assign x_46634 = x_15343 & x_46633;
assign x_46635 = x_15346 & x_15347;
assign x_46636 = x_15348 & x_15349;
assign x_46637 = x_46635 & x_46636;
assign x_46638 = x_46634 & x_46637;
assign x_46639 = x_15350 & x_15351;
assign x_46640 = x_15352 & x_15353;
assign x_46641 = x_46639 & x_46640;
assign x_46642 = x_15354 & x_15355;
assign x_46643 = x_15356 & x_15357;
assign x_46644 = x_46642 & x_46643;
assign x_46645 = x_46641 & x_46644;
assign x_46646 = x_46638 & x_46645;
assign x_46647 = x_15359 & x_15360;
assign x_46648 = x_15358 & x_46647;
assign x_46649 = x_15361 & x_15362;
assign x_46650 = x_15363 & x_15364;
assign x_46651 = x_46649 & x_46650;
assign x_46652 = x_46648 & x_46651;
assign x_46653 = x_15365 & x_15366;
assign x_46654 = x_15367 & x_15368;
assign x_46655 = x_46653 & x_46654;
assign x_46656 = x_15369 & x_15370;
assign x_46657 = x_15371 & x_15372;
assign x_46658 = x_46656 & x_46657;
assign x_46659 = x_46655 & x_46658;
assign x_46660 = x_46652 & x_46659;
assign x_46661 = x_46646 & x_46660;
assign x_46662 = x_15374 & x_15375;
assign x_46663 = x_15373 & x_46662;
assign x_46664 = x_15376 & x_15377;
assign x_46665 = x_15378 & x_15379;
assign x_46666 = x_46664 & x_46665;
assign x_46667 = x_46663 & x_46666;
assign x_46668 = x_15380 & x_15381;
assign x_46669 = x_15382 & x_15383;
assign x_46670 = x_46668 & x_46669;
assign x_46671 = x_15384 & x_15385;
assign x_46672 = x_15386 & x_15387;
assign x_46673 = x_46671 & x_46672;
assign x_46674 = x_46670 & x_46673;
assign x_46675 = x_46667 & x_46674;
assign x_46676 = x_15388 & x_15389;
assign x_46677 = x_15390 & x_15391;
assign x_46678 = x_46676 & x_46677;
assign x_46679 = x_15392 & x_15393;
assign x_46680 = x_15394 & x_15395;
assign x_46681 = x_46679 & x_46680;
assign x_46682 = x_46678 & x_46681;
assign x_46683 = x_15396 & x_15397;
assign x_46684 = x_15398 & x_15399;
assign x_46685 = x_46683 & x_46684;
assign x_46686 = x_15400 & x_15401;
assign x_46687 = x_15402 & x_15403;
assign x_46688 = x_46686 & x_46687;
assign x_46689 = x_46685 & x_46688;
assign x_46690 = x_46682 & x_46689;
assign x_46691 = x_46675 & x_46690;
assign x_46692 = x_46661 & x_46691;
assign x_46693 = x_46632 & x_46692;
assign x_46694 = x_46572 & x_46693;
assign x_46695 = x_15405 & x_15406;
assign x_46696 = x_15404 & x_46695;
assign x_46697 = x_15407 & x_15408;
assign x_46698 = x_15409 & x_15410;
assign x_46699 = x_46697 & x_46698;
assign x_46700 = x_46696 & x_46699;
assign x_46701 = x_15411 & x_15412;
assign x_46702 = x_15413 & x_15414;
assign x_46703 = x_46701 & x_46702;
assign x_46704 = x_15415 & x_15416;
assign x_46705 = x_15417 & x_15418;
assign x_46706 = x_46704 & x_46705;
assign x_46707 = x_46703 & x_46706;
assign x_46708 = x_46700 & x_46707;
assign x_46709 = x_15420 & x_15421;
assign x_46710 = x_15419 & x_46709;
assign x_46711 = x_15422 & x_15423;
assign x_46712 = x_15424 & x_15425;
assign x_46713 = x_46711 & x_46712;
assign x_46714 = x_46710 & x_46713;
assign x_46715 = x_15426 & x_15427;
assign x_46716 = x_15428 & x_15429;
assign x_46717 = x_46715 & x_46716;
assign x_46718 = x_15430 & x_15431;
assign x_46719 = x_15432 & x_15433;
assign x_46720 = x_46718 & x_46719;
assign x_46721 = x_46717 & x_46720;
assign x_46722 = x_46714 & x_46721;
assign x_46723 = x_46708 & x_46722;
assign x_46724 = x_15435 & x_15436;
assign x_46725 = x_15434 & x_46724;
assign x_46726 = x_15437 & x_15438;
assign x_46727 = x_15439 & x_15440;
assign x_46728 = x_46726 & x_46727;
assign x_46729 = x_46725 & x_46728;
assign x_46730 = x_15441 & x_15442;
assign x_46731 = x_15443 & x_15444;
assign x_46732 = x_46730 & x_46731;
assign x_46733 = x_15445 & x_15446;
assign x_46734 = x_15447 & x_15448;
assign x_46735 = x_46733 & x_46734;
assign x_46736 = x_46732 & x_46735;
assign x_46737 = x_46729 & x_46736;
assign x_46738 = x_15449 & x_15450;
assign x_46739 = x_15451 & x_15452;
assign x_46740 = x_46738 & x_46739;
assign x_46741 = x_15453 & x_15454;
assign x_46742 = x_15455 & x_15456;
assign x_46743 = x_46741 & x_46742;
assign x_46744 = x_46740 & x_46743;
assign x_46745 = x_15457 & x_15458;
assign x_46746 = x_15459 & x_15460;
assign x_46747 = x_46745 & x_46746;
assign x_46748 = x_15461 & x_15462;
assign x_46749 = x_15463 & x_15464;
assign x_46750 = x_46748 & x_46749;
assign x_46751 = x_46747 & x_46750;
assign x_46752 = x_46744 & x_46751;
assign x_46753 = x_46737 & x_46752;
assign x_46754 = x_46723 & x_46753;
assign x_46755 = x_15466 & x_15467;
assign x_46756 = x_15465 & x_46755;
assign x_46757 = x_15468 & x_15469;
assign x_46758 = x_15470 & x_15471;
assign x_46759 = x_46757 & x_46758;
assign x_46760 = x_46756 & x_46759;
assign x_46761 = x_15472 & x_15473;
assign x_46762 = x_15474 & x_15475;
assign x_46763 = x_46761 & x_46762;
assign x_46764 = x_15476 & x_15477;
assign x_46765 = x_15478 & x_15479;
assign x_46766 = x_46764 & x_46765;
assign x_46767 = x_46763 & x_46766;
assign x_46768 = x_46760 & x_46767;
assign x_46769 = x_15481 & x_15482;
assign x_46770 = x_15480 & x_46769;
assign x_46771 = x_15483 & x_15484;
assign x_46772 = x_15485 & x_15486;
assign x_46773 = x_46771 & x_46772;
assign x_46774 = x_46770 & x_46773;
assign x_46775 = x_15487 & x_15488;
assign x_46776 = x_15489 & x_15490;
assign x_46777 = x_46775 & x_46776;
assign x_46778 = x_15491 & x_15492;
assign x_46779 = x_15493 & x_15494;
assign x_46780 = x_46778 & x_46779;
assign x_46781 = x_46777 & x_46780;
assign x_46782 = x_46774 & x_46781;
assign x_46783 = x_46768 & x_46782;
assign x_46784 = x_15496 & x_15497;
assign x_46785 = x_15495 & x_46784;
assign x_46786 = x_15498 & x_15499;
assign x_46787 = x_15500 & x_15501;
assign x_46788 = x_46786 & x_46787;
assign x_46789 = x_46785 & x_46788;
assign x_46790 = x_15502 & x_15503;
assign x_46791 = x_15504 & x_15505;
assign x_46792 = x_46790 & x_46791;
assign x_46793 = x_15506 & x_15507;
assign x_46794 = x_15508 & x_15509;
assign x_46795 = x_46793 & x_46794;
assign x_46796 = x_46792 & x_46795;
assign x_46797 = x_46789 & x_46796;
assign x_46798 = x_15510 & x_15511;
assign x_46799 = x_15512 & x_15513;
assign x_46800 = x_46798 & x_46799;
assign x_46801 = x_15514 & x_15515;
assign x_46802 = x_15516 & x_15517;
assign x_46803 = x_46801 & x_46802;
assign x_46804 = x_46800 & x_46803;
assign x_46805 = x_15518 & x_15519;
assign x_46806 = x_15520 & x_15521;
assign x_46807 = x_46805 & x_46806;
assign x_46808 = x_15522 & x_15523;
assign x_46809 = x_15524 & x_15525;
assign x_46810 = x_46808 & x_46809;
assign x_46811 = x_46807 & x_46810;
assign x_46812 = x_46804 & x_46811;
assign x_46813 = x_46797 & x_46812;
assign x_46814 = x_46783 & x_46813;
assign x_46815 = x_46754 & x_46814;
assign x_46816 = x_15527 & x_15528;
assign x_46817 = x_15526 & x_46816;
assign x_46818 = x_15529 & x_15530;
assign x_46819 = x_15531 & x_15532;
assign x_46820 = x_46818 & x_46819;
assign x_46821 = x_46817 & x_46820;
assign x_46822 = x_15533 & x_15534;
assign x_46823 = x_15535 & x_15536;
assign x_46824 = x_46822 & x_46823;
assign x_46825 = x_15537 & x_15538;
assign x_46826 = x_15539 & x_15540;
assign x_46827 = x_46825 & x_46826;
assign x_46828 = x_46824 & x_46827;
assign x_46829 = x_46821 & x_46828;
assign x_46830 = x_15542 & x_15543;
assign x_46831 = x_15541 & x_46830;
assign x_46832 = x_15544 & x_15545;
assign x_46833 = x_15546 & x_15547;
assign x_46834 = x_46832 & x_46833;
assign x_46835 = x_46831 & x_46834;
assign x_46836 = x_15548 & x_15549;
assign x_46837 = x_15550 & x_15551;
assign x_46838 = x_46836 & x_46837;
assign x_46839 = x_15552 & x_15553;
assign x_46840 = x_15554 & x_15555;
assign x_46841 = x_46839 & x_46840;
assign x_46842 = x_46838 & x_46841;
assign x_46843 = x_46835 & x_46842;
assign x_46844 = x_46829 & x_46843;
assign x_46845 = x_15557 & x_15558;
assign x_46846 = x_15556 & x_46845;
assign x_46847 = x_15559 & x_15560;
assign x_46848 = x_15561 & x_15562;
assign x_46849 = x_46847 & x_46848;
assign x_46850 = x_46846 & x_46849;
assign x_46851 = x_15563 & x_15564;
assign x_46852 = x_15565 & x_15566;
assign x_46853 = x_46851 & x_46852;
assign x_46854 = x_15567 & x_15568;
assign x_46855 = x_15569 & x_15570;
assign x_46856 = x_46854 & x_46855;
assign x_46857 = x_46853 & x_46856;
assign x_46858 = x_46850 & x_46857;
assign x_46859 = x_15571 & x_15572;
assign x_46860 = x_15573 & x_15574;
assign x_46861 = x_46859 & x_46860;
assign x_46862 = x_15575 & x_15576;
assign x_46863 = x_15577 & x_15578;
assign x_46864 = x_46862 & x_46863;
assign x_46865 = x_46861 & x_46864;
assign x_46866 = x_15579 & x_15580;
assign x_46867 = x_15581 & x_15582;
assign x_46868 = x_46866 & x_46867;
assign x_46869 = x_15583 & x_15584;
assign x_46870 = x_15585 & x_15586;
assign x_46871 = x_46869 & x_46870;
assign x_46872 = x_46868 & x_46871;
assign x_46873 = x_46865 & x_46872;
assign x_46874 = x_46858 & x_46873;
assign x_46875 = x_46844 & x_46874;
assign x_46876 = x_15588 & x_15589;
assign x_46877 = x_15587 & x_46876;
assign x_46878 = x_15590 & x_15591;
assign x_46879 = x_15592 & x_15593;
assign x_46880 = x_46878 & x_46879;
assign x_46881 = x_46877 & x_46880;
assign x_46882 = x_15594 & x_15595;
assign x_46883 = x_15596 & x_15597;
assign x_46884 = x_46882 & x_46883;
assign x_46885 = x_15598 & x_15599;
assign x_46886 = x_15600 & x_15601;
assign x_46887 = x_46885 & x_46886;
assign x_46888 = x_46884 & x_46887;
assign x_46889 = x_46881 & x_46888;
assign x_46890 = x_15602 & x_15603;
assign x_46891 = x_15604 & x_15605;
assign x_46892 = x_46890 & x_46891;
assign x_46893 = x_15606 & x_15607;
assign x_46894 = x_15608 & x_15609;
assign x_46895 = x_46893 & x_46894;
assign x_46896 = x_46892 & x_46895;
assign x_46897 = x_15610 & x_15611;
assign x_46898 = x_15612 & x_15613;
assign x_46899 = x_46897 & x_46898;
assign x_46900 = x_15614 & x_15615;
assign x_46901 = x_15616 & x_15617;
assign x_46902 = x_46900 & x_46901;
assign x_46903 = x_46899 & x_46902;
assign x_46904 = x_46896 & x_46903;
assign x_46905 = x_46889 & x_46904;
assign x_46906 = x_15619 & x_15620;
assign x_46907 = x_15618 & x_46906;
assign x_46908 = x_15621 & x_15622;
assign x_46909 = x_15623 & x_15624;
assign x_46910 = x_46908 & x_46909;
assign x_46911 = x_46907 & x_46910;
assign x_46912 = x_15625 & x_15626;
assign x_46913 = x_15627 & x_15628;
assign x_46914 = x_46912 & x_46913;
assign x_46915 = x_15629 & x_15630;
assign x_46916 = x_15631 & x_15632;
assign x_46917 = x_46915 & x_46916;
assign x_46918 = x_46914 & x_46917;
assign x_46919 = x_46911 & x_46918;
assign x_46920 = x_15633 & x_15634;
assign x_46921 = x_15635 & x_15636;
assign x_46922 = x_46920 & x_46921;
assign x_46923 = x_15637 & x_15638;
assign x_46924 = x_15639 & x_15640;
assign x_46925 = x_46923 & x_46924;
assign x_46926 = x_46922 & x_46925;
assign x_46927 = x_15641 & x_15642;
assign x_46928 = x_15643 & x_15644;
assign x_46929 = x_46927 & x_46928;
assign x_46930 = x_15645 & x_15646;
assign x_46931 = x_15647 & x_15648;
assign x_46932 = x_46930 & x_46931;
assign x_46933 = x_46929 & x_46932;
assign x_46934 = x_46926 & x_46933;
assign x_46935 = x_46919 & x_46934;
assign x_46936 = x_46905 & x_46935;
assign x_46937 = x_46875 & x_46936;
assign x_46938 = x_46815 & x_46937;
assign x_46939 = x_46694 & x_46938;
assign x_46940 = x_46451 & x_46939;
assign x_46941 = x_45963 & x_46940;
assign x_46942 = x_44986 & x_46941;
assign x_46943 = x_43031 & x_46942;
assign x_46944 = x_39120 & x_46943;
assign x_46945 = x_15650 & x_15651;
assign x_46946 = x_15649 & x_46945;
assign x_46947 = x_15652 & x_15653;
assign x_46948 = x_15654 & x_15655;
assign x_46949 = x_46947 & x_46948;
assign x_46950 = x_46946 & x_46949;
assign x_46951 = x_15656 & x_15657;
assign x_46952 = x_15658 & x_15659;
assign x_46953 = x_46951 & x_46952;
assign x_46954 = x_15660 & x_15661;
assign x_46955 = x_15662 & x_15663;
assign x_46956 = x_46954 & x_46955;
assign x_46957 = x_46953 & x_46956;
assign x_46958 = x_46950 & x_46957;
assign x_46959 = x_15665 & x_15666;
assign x_46960 = x_15664 & x_46959;
assign x_46961 = x_15667 & x_15668;
assign x_46962 = x_15669 & x_15670;
assign x_46963 = x_46961 & x_46962;
assign x_46964 = x_46960 & x_46963;
assign x_46965 = x_15671 & x_15672;
assign x_46966 = x_15673 & x_15674;
assign x_46967 = x_46965 & x_46966;
assign x_46968 = x_15675 & x_15676;
assign x_46969 = x_15677 & x_15678;
assign x_46970 = x_46968 & x_46969;
assign x_46971 = x_46967 & x_46970;
assign x_46972 = x_46964 & x_46971;
assign x_46973 = x_46958 & x_46972;
assign x_46974 = x_15680 & x_15681;
assign x_46975 = x_15679 & x_46974;
assign x_46976 = x_15682 & x_15683;
assign x_46977 = x_15684 & x_15685;
assign x_46978 = x_46976 & x_46977;
assign x_46979 = x_46975 & x_46978;
assign x_46980 = x_15686 & x_15687;
assign x_46981 = x_15688 & x_15689;
assign x_46982 = x_46980 & x_46981;
assign x_46983 = x_15690 & x_15691;
assign x_46984 = x_15692 & x_15693;
assign x_46985 = x_46983 & x_46984;
assign x_46986 = x_46982 & x_46985;
assign x_46987 = x_46979 & x_46986;
assign x_46988 = x_15694 & x_15695;
assign x_46989 = x_15696 & x_15697;
assign x_46990 = x_46988 & x_46989;
assign x_46991 = x_15698 & x_15699;
assign x_46992 = x_15700 & x_15701;
assign x_46993 = x_46991 & x_46992;
assign x_46994 = x_46990 & x_46993;
assign x_46995 = x_15702 & x_15703;
assign x_46996 = x_15704 & x_15705;
assign x_46997 = x_46995 & x_46996;
assign x_46998 = x_15706 & x_15707;
assign x_46999 = x_15708 & x_15709;
assign x_47000 = x_46998 & x_46999;
assign x_47001 = x_46997 & x_47000;
assign x_47002 = x_46994 & x_47001;
assign x_47003 = x_46987 & x_47002;
assign x_47004 = x_46973 & x_47003;
assign x_47005 = x_15711 & x_15712;
assign x_47006 = x_15710 & x_47005;
assign x_47007 = x_15713 & x_15714;
assign x_47008 = x_15715 & x_15716;
assign x_47009 = x_47007 & x_47008;
assign x_47010 = x_47006 & x_47009;
assign x_47011 = x_15717 & x_15718;
assign x_47012 = x_15719 & x_15720;
assign x_47013 = x_47011 & x_47012;
assign x_47014 = x_15721 & x_15722;
assign x_47015 = x_15723 & x_15724;
assign x_47016 = x_47014 & x_47015;
assign x_47017 = x_47013 & x_47016;
assign x_47018 = x_47010 & x_47017;
assign x_47019 = x_15726 & x_15727;
assign x_47020 = x_15725 & x_47019;
assign x_47021 = x_15728 & x_15729;
assign x_47022 = x_15730 & x_15731;
assign x_47023 = x_47021 & x_47022;
assign x_47024 = x_47020 & x_47023;
assign x_47025 = x_15732 & x_15733;
assign x_47026 = x_15734 & x_15735;
assign x_47027 = x_47025 & x_47026;
assign x_47028 = x_15736 & x_15737;
assign x_47029 = x_15738 & x_15739;
assign x_47030 = x_47028 & x_47029;
assign x_47031 = x_47027 & x_47030;
assign x_47032 = x_47024 & x_47031;
assign x_47033 = x_47018 & x_47032;
assign x_47034 = x_15741 & x_15742;
assign x_47035 = x_15740 & x_47034;
assign x_47036 = x_15743 & x_15744;
assign x_47037 = x_15745 & x_15746;
assign x_47038 = x_47036 & x_47037;
assign x_47039 = x_47035 & x_47038;
assign x_47040 = x_15747 & x_15748;
assign x_47041 = x_15749 & x_15750;
assign x_47042 = x_47040 & x_47041;
assign x_47043 = x_15751 & x_15752;
assign x_47044 = x_15753 & x_15754;
assign x_47045 = x_47043 & x_47044;
assign x_47046 = x_47042 & x_47045;
assign x_47047 = x_47039 & x_47046;
assign x_47048 = x_15755 & x_15756;
assign x_47049 = x_15757 & x_15758;
assign x_47050 = x_47048 & x_47049;
assign x_47051 = x_15759 & x_15760;
assign x_47052 = x_15761 & x_15762;
assign x_47053 = x_47051 & x_47052;
assign x_47054 = x_47050 & x_47053;
assign x_47055 = x_15763 & x_15764;
assign x_47056 = x_15765 & x_15766;
assign x_47057 = x_47055 & x_47056;
assign x_47058 = x_15767 & x_15768;
assign x_47059 = x_15769 & x_15770;
assign x_47060 = x_47058 & x_47059;
assign x_47061 = x_47057 & x_47060;
assign x_47062 = x_47054 & x_47061;
assign x_47063 = x_47047 & x_47062;
assign x_47064 = x_47033 & x_47063;
assign x_47065 = x_47004 & x_47064;
assign x_47066 = x_15772 & x_15773;
assign x_47067 = x_15771 & x_47066;
assign x_47068 = x_15774 & x_15775;
assign x_47069 = x_15776 & x_15777;
assign x_47070 = x_47068 & x_47069;
assign x_47071 = x_47067 & x_47070;
assign x_47072 = x_15778 & x_15779;
assign x_47073 = x_15780 & x_15781;
assign x_47074 = x_47072 & x_47073;
assign x_47075 = x_15782 & x_15783;
assign x_47076 = x_15784 & x_15785;
assign x_47077 = x_47075 & x_47076;
assign x_47078 = x_47074 & x_47077;
assign x_47079 = x_47071 & x_47078;
assign x_47080 = x_15787 & x_15788;
assign x_47081 = x_15786 & x_47080;
assign x_47082 = x_15789 & x_15790;
assign x_47083 = x_15791 & x_15792;
assign x_47084 = x_47082 & x_47083;
assign x_47085 = x_47081 & x_47084;
assign x_47086 = x_15793 & x_15794;
assign x_47087 = x_15795 & x_15796;
assign x_47088 = x_47086 & x_47087;
assign x_47089 = x_15797 & x_15798;
assign x_47090 = x_15799 & x_15800;
assign x_47091 = x_47089 & x_47090;
assign x_47092 = x_47088 & x_47091;
assign x_47093 = x_47085 & x_47092;
assign x_47094 = x_47079 & x_47093;
assign x_47095 = x_15802 & x_15803;
assign x_47096 = x_15801 & x_47095;
assign x_47097 = x_15804 & x_15805;
assign x_47098 = x_15806 & x_15807;
assign x_47099 = x_47097 & x_47098;
assign x_47100 = x_47096 & x_47099;
assign x_47101 = x_15808 & x_15809;
assign x_47102 = x_15810 & x_15811;
assign x_47103 = x_47101 & x_47102;
assign x_47104 = x_15812 & x_15813;
assign x_47105 = x_15814 & x_15815;
assign x_47106 = x_47104 & x_47105;
assign x_47107 = x_47103 & x_47106;
assign x_47108 = x_47100 & x_47107;
assign x_47109 = x_15816 & x_15817;
assign x_47110 = x_15818 & x_15819;
assign x_47111 = x_47109 & x_47110;
assign x_47112 = x_15820 & x_15821;
assign x_47113 = x_15822 & x_15823;
assign x_47114 = x_47112 & x_47113;
assign x_47115 = x_47111 & x_47114;
assign x_47116 = x_15824 & x_15825;
assign x_47117 = x_15826 & x_15827;
assign x_47118 = x_47116 & x_47117;
assign x_47119 = x_15828 & x_15829;
assign x_47120 = x_15830 & x_15831;
assign x_47121 = x_47119 & x_47120;
assign x_47122 = x_47118 & x_47121;
assign x_47123 = x_47115 & x_47122;
assign x_47124 = x_47108 & x_47123;
assign x_47125 = x_47094 & x_47124;
assign x_47126 = x_15833 & x_15834;
assign x_47127 = x_15832 & x_47126;
assign x_47128 = x_15835 & x_15836;
assign x_47129 = x_15837 & x_15838;
assign x_47130 = x_47128 & x_47129;
assign x_47131 = x_47127 & x_47130;
assign x_47132 = x_15839 & x_15840;
assign x_47133 = x_15841 & x_15842;
assign x_47134 = x_47132 & x_47133;
assign x_47135 = x_15843 & x_15844;
assign x_47136 = x_15845 & x_15846;
assign x_47137 = x_47135 & x_47136;
assign x_47138 = x_47134 & x_47137;
assign x_47139 = x_47131 & x_47138;
assign x_47140 = x_15848 & x_15849;
assign x_47141 = x_15847 & x_47140;
assign x_47142 = x_15850 & x_15851;
assign x_47143 = x_15852 & x_15853;
assign x_47144 = x_47142 & x_47143;
assign x_47145 = x_47141 & x_47144;
assign x_47146 = x_15854 & x_15855;
assign x_47147 = x_15856 & x_15857;
assign x_47148 = x_47146 & x_47147;
assign x_47149 = x_15858 & x_15859;
assign x_47150 = x_15860 & x_15861;
assign x_47151 = x_47149 & x_47150;
assign x_47152 = x_47148 & x_47151;
assign x_47153 = x_47145 & x_47152;
assign x_47154 = x_47139 & x_47153;
assign x_47155 = x_15863 & x_15864;
assign x_47156 = x_15862 & x_47155;
assign x_47157 = x_15865 & x_15866;
assign x_47158 = x_15867 & x_15868;
assign x_47159 = x_47157 & x_47158;
assign x_47160 = x_47156 & x_47159;
assign x_47161 = x_15869 & x_15870;
assign x_47162 = x_15871 & x_15872;
assign x_47163 = x_47161 & x_47162;
assign x_47164 = x_15873 & x_15874;
assign x_47165 = x_15875 & x_15876;
assign x_47166 = x_47164 & x_47165;
assign x_47167 = x_47163 & x_47166;
assign x_47168 = x_47160 & x_47167;
assign x_47169 = x_15877 & x_15878;
assign x_47170 = x_15879 & x_15880;
assign x_47171 = x_47169 & x_47170;
assign x_47172 = x_15881 & x_15882;
assign x_47173 = x_15883 & x_15884;
assign x_47174 = x_47172 & x_47173;
assign x_47175 = x_47171 & x_47174;
assign x_47176 = x_15885 & x_15886;
assign x_47177 = x_15887 & x_15888;
assign x_47178 = x_47176 & x_47177;
assign x_47179 = x_15889 & x_15890;
assign x_47180 = x_15891 & x_15892;
assign x_47181 = x_47179 & x_47180;
assign x_47182 = x_47178 & x_47181;
assign x_47183 = x_47175 & x_47182;
assign x_47184 = x_47168 & x_47183;
assign x_47185 = x_47154 & x_47184;
assign x_47186 = x_47125 & x_47185;
assign x_47187 = x_47065 & x_47186;
assign x_47188 = x_15894 & x_15895;
assign x_47189 = x_15893 & x_47188;
assign x_47190 = x_15896 & x_15897;
assign x_47191 = x_15898 & x_15899;
assign x_47192 = x_47190 & x_47191;
assign x_47193 = x_47189 & x_47192;
assign x_47194 = x_15900 & x_15901;
assign x_47195 = x_15902 & x_15903;
assign x_47196 = x_47194 & x_47195;
assign x_47197 = x_15904 & x_15905;
assign x_47198 = x_15906 & x_15907;
assign x_47199 = x_47197 & x_47198;
assign x_47200 = x_47196 & x_47199;
assign x_47201 = x_47193 & x_47200;
assign x_47202 = x_15909 & x_15910;
assign x_47203 = x_15908 & x_47202;
assign x_47204 = x_15911 & x_15912;
assign x_47205 = x_15913 & x_15914;
assign x_47206 = x_47204 & x_47205;
assign x_47207 = x_47203 & x_47206;
assign x_47208 = x_15915 & x_15916;
assign x_47209 = x_15917 & x_15918;
assign x_47210 = x_47208 & x_47209;
assign x_47211 = x_15919 & x_15920;
assign x_47212 = x_15921 & x_15922;
assign x_47213 = x_47211 & x_47212;
assign x_47214 = x_47210 & x_47213;
assign x_47215 = x_47207 & x_47214;
assign x_47216 = x_47201 & x_47215;
assign x_47217 = x_15924 & x_15925;
assign x_47218 = x_15923 & x_47217;
assign x_47219 = x_15926 & x_15927;
assign x_47220 = x_15928 & x_15929;
assign x_47221 = x_47219 & x_47220;
assign x_47222 = x_47218 & x_47221;
assign x_47223 = x_15930 & x_15931;
assign x_47224 = x_15932 & x_15933;
assign x_47225 = x_47223 & x_47224;
assign x_47226 = x_15934 & x_15935;
assign x_47227 = x_15936 & x_15937;
assign x_47228 = x_47226 & x_47227;
assign x_47229 = x_47225 & x_47228;
assign x_47230 = x_47222 & x_47229;
assign x_47231 = x_15938 & x_15939;
assign x_47232 = x_15940 & x_15941;
assign x_47233 = x_47231 & x_47232;
assign x_47234 = x_15942 & x_15943;
assign x_47235 = x_15944 & x_15945;
assign x_47236 = x_47234 & x_47235;
assign x_47237 = x_47233 & x_47236;
assign x_47238 = x_15946 & x_15947;
assign x_47239 = x_15948 & x_15949;
assign x_47240 = x_47238 & x_47239;
assign x_47241 = x_15950 & x_15951;
assign x_47242 = x_15952 & x_15953;
assign x_47243 = x_47241 & x_47242;
assign x_47244 = x_47240 & x_47243;
assign x_47245 = x_47237 & x_47244;
assign x_47246 = x_47230 & x_47245;
assign x_47247 = x_47216 & x_47246;
assign x_47248 = x_15955 & x_15956;
assign x_47249 = x_15954 & x_47248;
assign x_47250 = x_15957 & x_15958;
assign x_47251 = x_15959 & x_15960;
assign x_47252 = x_47250 & x_47251;
assign x_47253 = x_47249 & x_47252;
assign x_47254 = x_15961 & x_15962;
assign x_47255 = x_15963 & x_15964;
assign x_47256 = x_47254 & x_47255;
assign x_47257 = x_15965 & x_15966;
assign x_47258 = x_15967 & x_15968;
assign x_47259 = x_47257 & x_47258;
assign x_47260 = x_47256 & x_47259;
assign x_47261 = x_47253 & x_47260;
assign x_47262 = x_15970 & x_15971;
assign x_47263 = x_15969 & x_47262;
assign x_47264 = x_15972 & x_15973;
assign x_47265 = x_15974 & x_15975;
assign x_47266 = x_47264 & x_47265;
assign x_47267 = x_47263 & x_47266;
assign x_47268 = x_15976 & x_15977;
assign x_47269 = x_15978 & x_15979;
assign x_47270 = x_47268 & x_47269;
assign x_47271 = x_15980 & x_15981;
assign x_47272 = x_15982 & x_15983;
assign x_47273 = x_47271 & x_47272;
assign x_47274 = x_47270 & x_47273;
assign x_47275 = x_47267 & x_47274;
assign x_47276 = x_47261 & x_47275;
assign x_47277 = x_15985 & x_15986;
assign x_47278 = x_15984 & x_47277;
assign x_47279 = x_15987 & x_15988;
assign x_47280 = x_15989 & x_15990;
assign x_47281 = x_47279 & x_47280;
assign x_47282 = x_47278 & x_47281;
assign x_47283 = x_15991 & x_15992;
assign x_47284 = x_15993 & x_15994;
assign x_47285 = x_47283 & x_47284;
assign x_47286 = x_15995 & x_15996;
assign x_47287 = x_15997 & x_15998;
assign x_47288 = x_47286 & x_47287;
assign x_47289 = x_47285 & x_47288;
assign x_47290 = x_47282 & x_47289;
assign x_47291 = x_15999 & x_16000;
assign x_47292 = x_16001 & x_16002;
assign x_47293 = x_47291 & x_47292;
assign x_47294 = x_16003 & x_16004;
assign x_47295 = x_16005 & x_16006;
assign x_47296 = x_47294 & x_47295;
assign x_47297 = x_47293 & x_47296;
assign x_47298 = x_16007 & x_16008;
assign x_47299 = x_16009 & x_16010;
assign x_47300 = x_47298 & x_47299;
assign x_47301 = x_16011 & x_16012;
assign x_47302 = x_16013 & x_16014;
assign x_47303 = x_47301 & x_47302;
assign x_47304 = x_47300 & x_47303;
assign x_47305 = x_47297 & x_47304;
assign x_47306 = x_47290 & x_47305;
assign x_47307 = x_47276 & x_47306;
assign x_47308 = x_47247 & x_47307;
assign x_47309 = x_16016 & x_16017;
assign x_47310 = x_16015 & x_47309;
assign x_47311 = x_16018 & x_16019;
assign x_47312 = x_16020 & x_16021;
assign x_47313 = x_47311 & x_47312;
assign x_47314 = x_47310 & x_47313;
assign x_47315 = x_16022 & x_16023;
assign x_47316 = x_16024 & x_16025;
assign x_47317 = x_47315 & x_47316;
assign x_47318 = x_16026 & x_16027;
assign x_47319 = x_16028 & x_16029;
assign x_47320 = x_47318 & x_47319;
assign x_47321 = x_47317 & x_47320;
assign x_47322 = x_47314 & x_47321;
assign x_47323 = x_16031 & x_16032;
assign x_47324 = x_16030 & x_47323;
assign x_47325 = x_16033 & x_16034;
assign x_47326 = x_16035 & x_16036;
assign x_47327 = x_47325 & x_47326;
assign x_47328 = x_47324 & x_47327;
assign x_47329 = x_16037 & x_16038;
assign x_47330 = x_16039 & x_16040;
assign x_47331 = x_47329 & x_47330;
assign x_47332 = x_16041 & x_16042;
assign x_47333 = x_16043 & x_16044;
assign x_47334 = x_47332 & x_47333;
assign x_47335 = x_47331 & x_47334;
assign x_47336 = x_47328 & x_47335;
assign x_47337 = x_47322 & x_47336;
assign x_47338 = x_16046 & x_16047;
assign x_47339 = x_16045 & x_47338;
assign x_47340 = x_16048 & x_16049;
assign x_47341 = x_16050 & x_16051;
assign x_47342 = x_47340 & x_47341;
assign x_47343 = x_47339 & x_47342;
assign x_47344 = x_16052 & x_16053;
assign x_47345 = x_16054 & x_16055;
assign x_47346 = x_47344 & x_47345;
assign x_47347 = x_16056 & x_16057;
assign x_47348 = x_16058 & x_16059;
assign x_47349 = x_47347 & x_47348;
assign x_47350 = x_47346 & x_47349;
assign x_47351 = x_47343 & x_47350;
assign x_47352 = x_16060 & x_16061;
assign x_47353 = x_16062 & x_16063;
assign x_47354 = x_47352 & x_47353;
assign x_47355 = x_16064 & x_16065;
assign x_47356 = x_16066 & x_16067;
assign x_47357 = x_47355 & x_47356;
assign x_47358 = x_47354 & x_47357;
assign x_47359 = x_16068 & x_16069;
assign x_47360 = x_16070 & x_16071;
assign x_47361 = x_47359 & x_47360;
assign x_47362 = x_16072 & x_16073;
assign x_47363 = x_16074 & x_16075;
assign x_47364 = x_47362 & x_47363;
assign x_47365 = x_47361 & x_47364;
assign x_47366 = x_47358 & x_47365;
assign x_47367 = x_47351 & x_47366;
assign x_47368 = x_47337 & x_47367;
assign x_47369 = x_16077 & x_16078;
assign x_47370 = x_16076 & x_47369;
assign x_47371 = x_16079 & x_16080;
assign x_47372 = x_16081 & x_16082;
assign x_47373 = x_47371 & x_47372;
assign x_47374 = x_47370 & x_47373;
assign x_47375 = x_16083 & x_16084;
assign x_47376 = x_16085 & x_16086;
assign x_47377 = x_47375 & x_47376;
assign x_47378 = x_16087 & x_16088;
assign x_47379 = x_16089 & x_16090;
assign x_47380 = x_47378 & x_47379;
assign x_47381 = x_47377 & x_47380;
assign x_47382 = x_47374 & x_47381;
assign x_47383 = x_16091 & x_16092;
assign x_47384 = x_16093 & x_16094;
assign x_47385 = x_47383 & x_47384;
assign x_47386 = x_16095 & x_16096;
assign x_47387 = x_16097 & x_16098;
assign x_47388 = x_47386 & x_47387;
assign x_47389 = x_47385 & x_47388;
assign x_47390 = x_16099 & x_16100;
assign x_47391 = x_16101 & x_16102;
assign x_47392 = x_47390 & x_47391;
assign x_47393 = x_16103 & x_16104;
assign x_47394 = x_16105 & x_16106;
assign x_47395 = x_47393 & x_47394;
assign x_47396 = x_47392 & x_47395;
assign x_47397 = x_47389 & x_47396;
assign x_47398 = x_47382 & x_47397;
assign x_47399 = x_16108 & x_16109;
assign x_47400 = x_16107 & x_47399;
assign x_47401 = x_16110 & x_16111;
assign x_47402 = x_16112 & x_16113;
assign x_47403 = x_47401 & x_47402;
assign x_47404 = x_47400 & x_47403;
assign x_47405 = x_16114 & x_16115;
assign x_47406 = x_16116 & x_16117;
assign x_47407 = x_47405 & x_47406;
assign x_47408 = x_16118 & x_16119;
assign x_47409 = x_16120 & x_16121;
assign x_47410 = x_47408 & x_47409;
assign x_47411 = x_47407 & x_47410;
assign x_47412 = x_47404 & x_47411;
assign x_47413 = x_16122 & x_16123;
assign x_47414 = x_16124 & x_16125;
assign x_47415 = x_47413 & x_47414;
assign x_47416 = x_16126 & x_16127;
assign x_47417 = x_16128 & x_16129;
assign x_47418 = x_47416 & x_47417;
assign x_47419 = x_47415 & x_47418;
assign x_47420 = x_16130 & x_16131;
assign x_47421 = x_16132 & x_16133;
assign x_47422 = x_47420 & x_47421;
assign x_47423 = x_16134 & x_16135;
assign x_47424 = x_16136 & x_16137;
assign x_47425 = x_47423 & x_47424;
assign x_47426 = x_47422 & x_47425;
assign x_47427 = x_47419 & x_47426;
assign x_47428 = x_47412 & x_47427;
assign x_47429 = x_47398 & x_47428;
assign x_47430 = x_47368 & x_47429;
assign x_47431 = x_47308 & x_47430;
assign x_47432 = x_47187 & x_47431;
assign x_47433 = x_16139 & x_16140;
assign x_47434 = x_16138 & x_47433;
assign x_47435 = x_16141 & x_16142;
assign x_47436 = x_16143 & x_16144;
assign x_47437 = x_47435 & x_47436;
assign x_47438 = x_47434 & x_47437;
assign x_47439 = x_16145 & x_16146;
assign x_47440 = x_16147 & x_16148;
assign x_47441 = x_47439 & x_47440;
assign x_47442 = x_16149 & x_16150;
assign x_47443 = x_16151 & x_16152;
assign x_47444 = x_47442 & x_47443;
assign x_47445 = x_47441 & x_47444;
assign x_47446 = x_47438 & x_47445;
assign x_47447 = x_16154 & x_16155;
assign x_47448 = x_16153 & x_47447;
assign x_47449 = x_16156 & x_16157;
assign x_47450 = x_16158 & x_16159;
assign x_47451 = x_47449 & x_47450;
assign x_47452 = x_47448 & x_47451;
assign x_47453 = x_16160 & x_16161;
assign x_47454 = x_16162 & x_16163;
assign x_47455 = x_47453 & x_47454;
assign x_47456 = x_16164 & x_16165;
assign x_47457 = x_16166 & x_16167;
assign x_47458 = x_47456 & x_47457;
assign x_47459 = x_47455 & x_47458;
assign x_47460 = x_47452 & x_47459;
assign x_47461 = x_47446 & x_47460;
assign x_47462 = x_16169 & x_16170;
assign x_47463 = x_16168 & x_47462;
assign x_47464 = x_16171 & x_16172;
assign x_47465 = x_16173 & x_16174;
assign x_47466 = x_47464 & x_47465;
assign x_47467 = x_47463 & x_47466;
assign x_47468 = x_16175 & x_16176;
assign x_47469 = x_16177 & x_16178;
assign x_47470 = x_47468 & x_47469;
assign x_47471 = x_16179 & x_16180;
assign x_47472 = x_16181 & x_16182;
assign x_47473 = x_47471 & x_47472;
assign x_47474 = x_47470 & x_47473;
assign x_47475 = x_47467 & x_47474;
assign x_47476 = x_16183 & x_16184;
assign x_47477 = x_16185 & x_16186;
assign x_47478 = x_47476 & x_47477;
assign x_47479 = x_16187 & x_16188;
assign x_47480 = x_16189 & x_16190;
assign x_47481 = x_47479 & x_47480;
assign x_47482 = x_47478 & x_47481;
assign x_47483 = x_16191 & x_16192;
assign x_47484 = x_16193 & x_16194;
assign x_47485 = x_47483 & x_47484;
assign x_47486 = x_16195 & x_16196;
assign x_47487 = x_16197 & x_16198;
assign x_47488 = x_47486 & x_47487;
assign x_47489 = x_47485 & x_47488;
assign x_47490 = x_47482 & x_47489;
assign x_47491 = x_47475 & x_47490;
assign x_47492 = x_47461 & x_47491;
assign x_47493 = x_16200 & x_16201;
assign x_47494 = x_16199 & x_47493;
assign x_47495 = x_16202 & x_16203;
assign x_47496 = x_16204 & x_16205;
assign x_47497 = x_47495 & x_47496;
assign x_47498 = x_47494 & x_47497;
assign x_47499 = x_16206 & x_16207;
assign x_47500 = x_16208 & x_16209;
assign x_47501 = x_47499 & x_47500;
assign x_47502 = x_16210 & x_16211;
assign x_47503 = x_16212 & x_16213;
assign x_47504 = x_47502 & x_47503;
assign x_47505 = x_47501 & x_47504;
assign x_47506 = x_47498 & x_47505;
assign x_47507 = x_16215 & x_16216;
assign x_47508 = x_16214 & x_47507;
assign x_47509 = x_16217 & x_16218;
assign x_47510 = x_16219 & x_16220;
assign x_47511 = x_47509 & x_47510;
assign x_47512 = x_47508 & x_47511;
assign x_47513 = x_16221 & x_16222;
assign x_47514 = x_16223 & x_16224;
assign x_47515 = x_47513 & x_47514;
assign x_47516 = x_16225 & x_16226;
assign x_47517 = x_16227 & x_16228;
assign x_47518 = x_47516 & x_47517;
assign x_47519 = x_47515 & x_47518;
assign x_47520 = x_47512 & x_47519;
assign x_47521 = x_47506 & x_47520;
assign x_47522 = x_16230 & x_16231;
assign x_47523 = x_16229 & x_47522;
assign x_47524 = x_16232 & x_16233;
assign x_47525 = x_16234 & x_16235;
assign x_47526 = x_47524 & x_47525;
assign x_47527 = x_47523 & x_47526;
assign x_47528 = x_16236 & x_16237;
assign x_47529 = x_16238 & x_16239;
assign x_47530 = x_47528 & x_47529;
assign x_47531 = x_16240 & x_16241;
assign x_47532 = x_16242 & x_16243;
assign x_47533 = x_47531 & x_47532;
assign x_47534 = x_47530 & x_47533;
assign x_47535 = x_47527 & x_47534;
assign x_47536 = x_16244 & x_16245;
assign x_47537 = x_16246 & x_16247;
assign x_47538 = x_47536 & x_47537;
assign x_47539 = x_16248 & x_16249;
assign x_47540 = x_16250 & x_16251;
assign x_47541 = x_47539 & x_47540;
assign x_47542 = x_47538 & x_47541;
assign x_47543 = x_16252 & x_16253;
assign x_47544 = x_16254 & x_16255;
assign x_47545 = x_47543 & x_47544;
assign x_47546 = x_16256 & x_16257;
assign x_47547 = x_16258 & x_16259;
assign x_47548 = x_47546 & x_47547;
assign x_47549 = x_47545 & x_47548;
assign x_47550 = x_47542 & x_47549;
assign x_47551 = x_47535 & x_47550;
assign x_47552 = x_47521 & x_47551;
assign x_47553 = x_47492 & x_47552;
assign x_47554 = x_16261 & x_16262;
assign x_47555 = x_16260 & x_47554;
assign x_47556 = x_16263 & x_16264;
assign x_47557 = x_16265 & x_16266;
assign x_47558 = x_47556 & x_47557;
assign x_47559 = x_47555 & x_47558;
assign x_47560 = x_16267 & x_16268;
assign x_47561 = x_16269 & x_16270;
assign x_47562 = x_47560 & x_47561;
assign x_47563 = x_16271 & x_16272;
assign x_47564 = x_16273 & x_16274;
assign x_47565 = x_47563 & x_47564;
assign x_47566 = x_47562 & x_47565;
assign x_47567 = x_47559 & x_47566;
assign x_47568 = x_16276 & x_16277;
assign x_47569 = x_16275 & x_47568;
assign x_47570 = x_16278 & x_16279;
assign x_47571 = x_16280 & x_16281;
assign x_47572 = x_47570 & x_47571;
assign x_47573 = x_47569 & x_47572;
assign x_47574 = x_16282 & x_16283;
assign x_47575 = x_16284 & x_16285;
assign x_47576 = x_47574 & x_47575;
assign x_47577 = x_16286 & x_16287;
assign x_47578 = x_16288 & x_16289;
assign x_47579 = x_47577 & x_47578;
assign x_47580 = x_47576 & x_47579;
assign x_47581 = x_47573 & x_47580;
assign x_47582 = x_47567 & x_47581;
assign x_47583 = x_16291 & x_16292;
assign x_47584 = x_16290 & x_47583;
assign x_47585 = x_16293 & x_16294;
assign x_47586 = x_16295 & x_16296;
assign x_47587 = x_47585 & x_47586;
assign x_47588 = x_47584 & x_47587;
assign x_47589 = x_16297 & x_16298;
assign x_47590 = x_16299 & x_16300;
assign x_47591 = x_47589 & x_47590;
assign x_47592 = x_16301 & x_16302;
assign x_47593 = x_16303 & x_16304;
assign x_47594 = x_47592 & x_47593;
assign x_47595 = x_47591 & x_47594;
assign x_47596 = x_47588 & x_47595;
assign x_47597 = x_16305 & x_16306;
assign x_47598 = x_16307 & x_16308;
assign x_47599 = x_47597 & x_47598;
assign x_47600 = x_16309 & x_16310;
assign x_47601 = x_16311 & x_16312;
assign x_47602 = x_47600 & x_47601;
assign x_47603 = x_47599 & x_47602;
assign x_47604 = x_16313 & x_16314;
assign x_47605 = x_16315 & x_16316;
assign x_47606 = x_47604 & x_47605;
assign x_47607 = x_16317 & x_16318;
assign x_47608 = x_16319 & x_16320;
assign x_47609 = x_47607 & x_47608;
assign x_47610 = x_47606 & x_47609;
assign x_47611 = x_47603 & x_47610;
assign x_47612 = x_47596 & x_47611;
assign x_47613 = x_47582 & x_47612;
assign x_47614 = x_16322 & x_16323;
assign x_47615 = x_16321 & x_47614;
assign x_47616 = x_16324 & x_16325;
assign x_47617 = x_16326 & x_16327;
assign x_47618 = x_47616 & x_47617;
assign x_47619 = x_47615 & x_47618;
assign x_47620 = x_16328 & x_16329;
assign x_47621 = x_16330 & x_16331;
assign x_47622 = x_47620 & x_47621;
assign x_47623 = x_16332 & x_16333;
assign x_47624 = x_16334 & x_16335;
assign x_47625 = x_47623 & x_47624;
assign x_47626 = x_47622 & x_47625;
assign x_47627 = x_47619 & x_47626;
assign x_47628 = x_16337 & x_16338;
assign x_47629 = x_16336 & x_47628;
assign x_47630 = x_16339 & x_16340;
assign x_47631 = x_16341 & x_16342;
assign x_47632 = x_47630 & x_47631;
assign x_47633 = x_47629 & x_47632;
assign x_47634 = x_16343 & x_16344;
assign x_47635 = x_16345 & x_16346;
assign x_47636 = x_47634 & x_47635;
assign x_47637 = x_16347 & x_16348;
assign x_47638 = x_16349 & x_16350;
assign x_47639 = x_47637 & x_47638;
assign x_47640 = x_47636 & x_47639;
assign x_47641 = x_47633 & x_47640;
assign x_47642 = x_47627 & x_47641;
assign x_47643 = x_16352 & x_16353;
assign x_47644 = x_16351 & x_47643;
assign x_47645 = x_16354 & x_16355;
assign x_47646 = x_16356 & x_16357;
assign x_47647 = x_47645 & x_47646;
assign x_47648 = x_47644 & x_47647;
assign x_47649 = x_16358 & x_16359;
assign x_47650 = x_16360 & x_16361;
assign x_47651 = x_47649 & x_47650;
assign x_47652 = x_16362 & x_16363;
assign x_47653 = x_16364 & x_16365;
assign x_47654 = x_47652 & x_47653;
assign x_47655 = x_47651 & x_47654;
assign x_47656 = x_47648 & x_47655;
assign x_47657 = x_16366 & x_16367;
assign x_47658 = x_16368 & x_16369;
assign x_47659 = x_47657 & x_47658;
assign x_47660 = x_16370 & x_16371;
assign x_47661 = x_16372 & x_16373;
assign x_47662 = x_47660 & x_47661;
assign x_47663 = x_47659 & x_47662;
assign x_47664 = x_16374 & x_16375;
assign x_47665 = x_16376 & x_16377;
assign x_47666 = x_47664 & x_47665;
assign x_47667 = x_16378 & x_16379;
assign x_47668 = x_16380 & x_16381;
assign x_47669 = x_47667 & x_47668;
assign x_47670 = x_47666 & x_47669;
assign x_47671 = x_47663 & x_47670;
assign x_47672 = x_47656 & x_47671;
assign x_47673 = x_47642 & x_47672;
assign x_47674 = x_47613 & x_47673;
assign x_47675 = x_47553 & x_47674;
assign x_47676 = x_16383 & x_16384;
assign x_47677 = x_16382 & x_47676;
assign x_47678 = x_16385 & x_16386;
assign x_47679 = x_16387 & x_16388;
assign x_47680 = x_47678 & x_47679;
assign x_47681 = x_47677 & x_47680;
assign x_47682 = x_16389 & x_16390;
assign x_47683 = x_16391 & x_16392;
assign x_47684 = x_47682 & x_47683;
assign x_47685 = x_16393 & x_16394;
assign x_47686 = x_16395 & x_16396;
assign x_47687 = x_47685 & x_47686;
assign x_47688 = x_47684 & x_47687;
assign x_47689 = x_47681 & x_47688;
assign x_47690 = x_16398 & x_16399;
assign x_47691 = x_16397 & x_47690;
assign x_47692 = x_16400 & x_16401;
assign x_47693 = x_16402 & x_16403;
assign x_47694 = x_47692 & x_47693;
assign x_47695 = x_47691 & x_47694;
assign x_47696 = x_16404 & x_16405;
assign x_47697 = x_16406 & x_16407;
assign x_47698 = x_47696 & x_47697;
assign x_47699 = x_16408 & x_16409;
assign x_47700 = x_16410 & x_16411;
assign x_47701 = x_47699 & x_47700;
assign x_47702 = x_47698 & x_47701;
assign x_47703 = x_47695 & x_47702;
assign x_47704 = x_47689 & x_47703;
assign x_47705 = x_16413 & x_16414;
assign x_47706 = x_16412 & x_47705;
assign x_47707 = x_16415 & x_16416;
assign x_47708 = x_16417 & x_16418;
assign x_47709 = x_47707 & x_47708;
assign x_47710 = x_47706 & x_47709;
assign x_47711 = x_16419 & x_16420;
assign x_47712 = x_16421 & x_16422;
assign x_47713 = x_47711 & x_47712;
assign x_47714 = x_16423 & x_16424;
assign x_47715 = x_16425 & x_16426;
assign x_47716 = x_47714 & x_47715;
assign x_47717 = x_47713 & x_47716;
assign x_47718 = x_47710 & x_47717;
assign x_47719 = x_16427 & x_16428;
assign x_47720 = x_16429 & x_16430;
assign x_47721 = x_47719 & x_47720;
assign x_47722 = x_16431 & x_16432;
assign x_47723 = x_16433 & x_16434;
assign x_47724 = x_47722 & x_47723;
assign x_47725 = x_47721 & x_47724;
assign x_47726 = x_16435 & x_16436;
assign x_47727 = x_16437 & x_16438;
assign x_47728 = x_47726 & x_47727;
assign x_47729 = x_16439 & x_16440;
assign x_47730 = x_16441 & x_16442;
assign x_47731 = x_47729 & x_47730;
assign x_47732 = x_47728 & x_47731;
assign x_47733 = x_47725 & x_47732;
assign x_47734 = x_47718 & x_47733;
assign x_47735 = x_47704 & x_47734;
assign x_47736 = x_16444 & x_16445;
assign x_47737 = x_16443 & x_47736;
assign x_47738 = x_16446 & x_16447;
assign x_47739 = x_16448 & x_16449;
assign x_47740 = x_47738 & x_47739;
assign x_47741 = x_47737 & x_47740;
assign x_47742 = x_16450 & x_16451;
assign x_47743 = x_16452 & x_16453;
assign x_47744 = x_47742 & x_47743;
assign x_47745 = x_16454 & x_16455;
assign x_47746 = x_16456 & x_16457;
assign x_47747 = x_47745 & x_47746;
assign x_47748 = x_47744 & x_47747;
assign x_47749 = x_47741 & x_47748;
assign x_47750 = x_16459 & x_16460;
assign x_47751 = x_16458 & x_47750;
assign x_47752 = x_16461 & x_16462;
assign x_47753 = x_16463 & x_16464;
assign x_47754 = x_47752 & x_47753;
assign x_47755 = x_47751 & x_47754;
assign x_47756 = x_16465 & x_16466;
assign x_47757 = x_16467 & x_16468;
assign x_47758 = x_47756 & x_47757;
assign x_47759 = x_16469 & x_16470;
assign x_47760 = x_16471 & x_16472;
assign x_47761 = x_47759 & x_47760;
assign x_47762 = x_47758 & x_47761;
assign x_47763 = x_47755 & x_47762;
assign x_47764 = x_47749 & x_47763;
assign x_47765 = x_16474 & x_16475;
assign x_47766 = x_16473 & x_47765;
assign x_47767 = x_16476 & x_16477;
assign x_47768 = x_16478 & x_16479;
assign x_47769 = x_47767 & x_47768;
assign x_47770 = x_47766 & x_47769;
assign x_47771 = x_16480 & x_16481;
assign x_47772 = x_16482 & x_16483;
assign x_47773 = x_47771 & x_47772;
assign x_47774 = x_16484 & x_16485;
assign x_47775 = x_16486 & x_16487;
assign x_47776 = x_47774 & x_47775;
assign x_47777 = x_47773 & x_47776;
assign x_47778 = x_47770 & x_47777;
assign x_47779 = x_16488 & x_16489;
assign x_47780 = x_16490 & x_16491;
assign x_47781 = x_47779 & x_47780;
assign x_47782 = x_16492 & x_16493;
assign x_47783 = x_16494 & x_16495;
assign x_47784 = x_47782 & x_47783;
assign x_47785 = x_47781 & x_47784;
assign x_47786 = x_16496 & x_16497;
assign x_47787 = x_16498 & x_16499;
assign x_47788 = x_47786 & x_47787;
assign x_47789 = x_16500 & x_16501;
assign x_47790 = x_16502 & x_16503;
assign x_47791 = x_47789 & x_47790;
assign x_47792 = x_47788 & x_47791;
assign x_47793 = x_47785 & x_47792;
assign x_47794 = x_47778 & x_47793;
assign x_47795 = x_47764 & x_47794;
assign x_47796 = x_47735 & x_47795;
assign x_47797 = x_16505 & x_16506;
assign x_47798 = x_16504 & x_47797;
assign x_47799 = x_16507 & x_16508;
assign x_47800 = x_16509 & x_16510;
assign x_47801 = x_47799 & x_47800;
assign x_47802 = x_47798 & x_47801;
assign x_47803 = x_16511 & x_16512;
assign x_47804 = x_16513 & x_16514;
assign x_47805 = x_47803 & x_47804;
assign x_47806 = x_16515 & x_16516;
assign x_47807 = x_16517 & x_16518;
assign x_47808 = x_47806 & x_47807;
assign x_47809 = x_47805 & x_47808;
assign x_47810 = x_47802 & x_47809;
assign x_47811 = x_16520 & x_16521;
assign x_47812 = x_16519 & x_47811;
assign x_47813 = x_16522 & x_16523;
assign x_47814 = x_16524 & x_16525;
assign x_47815 = x_47813 & x_47814;
assign x_47816 = x_47812 & x_47815;
assign x_47817 = x_16526 & x_16527;
assign x_47818 = x_16528 & x_16529;
assign x_47819 = x_47817 & x_47818;
assign x_47820 = x_16530 & x_16531;
assign x_47821 = x_16532 & x_16533;
assign x_47822 = x_47820 & x_47821;
assign x_47823 = x_47819 & x_47822;
assign x_47824 = x_47816 & x_47823;
assign x_47825 = x_47810 & x_47824;
assign x_47826 = x_16535 & x_16536;
assign x_47827 = x_16534 & x_47826;
assign x_47828 = x_16537 & x_16538;
assign x_47829 = x_16539 & x_16540;
assign x_47830 = x_47828 & x_47829;
assign x_47831 = x_47827 & x_47830;
assign x_47832 = x_16541 & x_16542;
assign x_47833 = x_16543 & x_16544;
assign x_47834 = x_47832 & x_47833;
assign x_47835 = x_16545 & x_16546;
assign x_47836 = x_16547 & x_16548;
assign x_47837 = x_47835 & x_47836;
assign x_47838 = x_47834 & x_47837;
assign x_47839 = x_47831 & x_47838;
assign x_47840 = x_16549 & x_16550;
assign x_47841 = x_16551 & x_16552;
assign x_47842 = x_47840 & x_47841;
assign x_47843 = x_16553 & x_16554;
assign x_47844 = x_16555 & x_16556;
assign x_47845 = x_47843 & x_47844;
assign x_47846 = x_47842 & x_47845;
assign x_47847 = x_16557 & x_16558;
assign x_47848 = x_16559 & x_16560;
assign x_47849 = x_47847 & x_47848;
assign x_47850 = x_16561 & x_16562;
assign x_47851 = x_16563 & x_16564;
assign x_47852 = x_47850 & x_47851;
assign x_47853 = x_47849 & x_47852;
assign x_47854 = x_47846 & x_47853;
assign x_47855 = x_47839 & x_47854;
assign x_47856 = x_47825 & x_47855;
assign x_47857 = x_16566 & x_16567;
assign x_47858 = x_16565 & x_47857;
assign x_47859 = x_16568 & x_16569;
assign x_47860 = x_16570 & x_16571;
assign x_47861 = x_47859 & x_47860;
assign x_47862 = x_47858 & x_47861;
assign x_47863 = x_16572 & x_16573;
assign x_47864 = x_16574 & x_16575;
assign x_47865 = x_47863 & x_47864;
assign x_47866 = x_16576 & x_16577;
assign x_47867 = x_16578 & x_16579;
assign x_47868 = x_47866 & x_47867;
assign x_47869 = x_47865 & x_47868;
assign x_47870 = x_47862 & x_47869;
assign x_47871 = x_16580 & x_16581;
assign x_47872 = x_16582 & x_16583;
assign x_47873 = x_47871 & x_47872;
assign x_47874 = x_16584 & x_16585;
assign x_47875 = x_16586 & x_16587;
assign x_47876 = x_47874 & x_47875;
assign x_47877 = x_47873 & x_47876;
assign x_47878 = x_16588 & x_16589;
assign x_47879 = x_16590 & x_16591;
assign x_47880 = x_47878 & x_47879;
assign x_47881 = x_16592 & x_16593;
assign x_47882 = x_16594 & x_16595;
assign x_47883 = x_47881 & x_47882;
assign x_47884 = x_47880 & x_47883;
assign x_47885 = x_47877 & x_47884;
assign x_47886 = x_47870 & x_47885;
assign x_47887 = x_16597 & x_16598;
assign x_47888 = x_16596 & x_47887;
assign x_47889 = x_16599 & x_16600;
assign x_47890 = x_16601 & x_16602;
assign x_47891 = x_47889 & x_47890;
assign x_47892 = x_47888 & x_47891;
assign x_47893 = x_16603 & x_16604;
assign x_47894 = x_16605 & x_16606;
assign x_47895 = x_47893 & x_47894;
assign x_47896 = x_16607 & x_16608;
assign x_47897 = x_16609 & x_16610;
assign x_47898 = x_47896 & x_47897;
assign x_47899 = x_47895 & x_47898;
assign x_47900 = x_47892 & x_47899;
assign x_47901 = x_16611 & x_16612;
assign x_47902 = x_16613 & x_16614;
assign x_47903 = x_47901 & x_47902;
assign x_47904 = x_16615 & x_16616;
assign x_47905 = x_16617 & x_16618;
assign x_47906 = x_47904 & x_47905;
assign x_47907 = x_47903 & x_47906;
assign x_47908 = x_16619 & x_16620;
assign x_47909 = x_16621 & x_16622;
assign x_47910 = x_47908 & x_47909;
assign x_47911 = x_16623 & x_16624;
assign x_47912 = x_16625 & x_16626;
assign x_47913 = x_47911 & x_47912;
assign x_47914 = x_47910 & x_47913;
assign x_47915 = x_47907 & x_47914;
assign x_47916 = x_47900 & x_47915;
assign x_47917 = x_47886 & x_47916;
assign x_47918 = x_47856 & x_47917;
assign x_47919 = x_47796 & x_47918;
assign x_47920 = x_47675 & x_47919;
assign x_47921 = x_47432 & x_47920;
assign x_47922 = x_16628 & x_16629;
assign x_47923 = x_16627 & x_47922;
assign x_47924 = x_16630 & x_16631;
assign x_47925 = x_16632 & x_16633;
assign x_47926 = x_47924 & x_47925;
assign x_47927 = x_47923 & x_47926;
assign x_47928 = x_16634 & x_16635;
assign x_47929 = x_16636 & x_16637;
assign x_47930 = x_47928 & x_47929;
assign x_47931 = x_16638 & x_16639;
assign x_47932 = x_16640 & x_16641;
assign x_47933 = x_47931 & x_47932;
assign x_47934 = x_47930 & x_47933;
assign x_47935 = x_47927 & x_47934;
assign x_47936 = x_16643 & x_16644;
assign x_47937 = x_16642 & x_47936;
assign x_47938 = x_16645 & x_16646;
assign x_47939 = x_16647 & x_16648;
assign x_47940 = x_47938 & x_47939;
assign x_47941 = x_47937 & x_47940;
assign x_47942 = x_16649 & x_16650;
assign x_47943 = x_16651 & x_16652;
assign x_47944 = x_47942 & x_47943;
assign x_47945 = x_16653 & x_16654;
assign x_47946 = x_16655 & x_16656;
assign x_47947 = x_47945 & x_47946;
assign x_47948 = x_47944 & x_47947;
assign x_47949 = x_47941 & x_47948;
assign x_47950 = x_47935 & x_47949;
assign x_47951 = x_16658 & x_16659;
assign x_47952 = x_16657 & x_47951;
assign x_47953 = x_16660 & x_16661;
assign x_47954 = x_16662 & x_16663;
assign x_47955 = x_47953 & x_47954;
assign x_47956 = x_47952 & x_47955;
assign x_47957 = x_16664 & x_16665;
assign x_47958 = x_16666 & x_16667;
assign x_47959 = x_47957 & x_47958;
assign x_47960 = x_16668 & x_16669;
assign x_47961 = x_16670 & x_16671;
assign x_47962 = x_47960 & x_47961;
assign x_47963 = x_47959 & x_47962;
assign x_47964 = x_47956 & x_47963;
assign x_47965 = x_16672 & x_16673;
assign x_47966 = x_16674 & x_16675;
assign x_47967 = x_47965 & x_47966;
assign x_47968 = x_16676 & x_16677;
assign x_47969 = x_16678 & x_16679;
assign x_47970 = x_47968 & x_47969;
assign x_47971 = x_47967 & x_47970;
assign x_47972 = x_16680 & x_16681;
assign x_47973 = x_16682 & x_16683;
assign x_47974 = x_47972 & x_47973;
assign x_47975 = x_16684 & x_16685;
assign x_47976 = x_16686 & x_16687;
assign x_47977 = x_47975 & x_47976;
assign x_47978 = x_47974 & x_47977;
assign x_47979 = x_47971 & x_47978;
assign x_47980 = x_47964 & x_47979;
assign x_47981 = x_47950 & x_47980;
assign x_47982 = x_16689 & x_16690;
assign x_47983 = x_16688 & x_47982;
assign x_47984 = x_16691 & x_16692;
assign x_47985 = x_16693 & x_16694;
assign x_47986 = x_47984 & x_47985;
assign x_47987 = x_47983 & x_47986;
assign x_47988 = x_16695 & x_16696;
assign x_47989 = x_16697 & x_16698;
assign x_47990 = x_47988 & x_47989;
assign x_47991 = x_16699 & x_16700;
assign x_47992 = x_16701 & x_16702;
assign x_47993 = x_47991 & x_47992;
assign x_47994 = x_47990 & x_47993;
assign x_47995 = x_47987 & x_47994;
assign x_47996 = x_16704 & x_16705;
assign x_47997 = x_16703 & x_47996;
assign x_47998 = x_16706 & x_16707;
assign x_47999 = x_16708 & x_16709;
assign x_48000 = x_47998 & x_47999;
assign x_48001 = x_47997 & x_48000;
assign x_48002 = x_16710 & x_16711;
assign x_48003 = x_16712 & x_16713;
assign x_48004 = x_48002 & x_48003;
assign x_48005 = x_16714 & x_16715;
assign x_48006 = x_16716 & x_16717;
assign x_48007 = x_48005 & x_48006;
assign x_48008 = x_48004 & x_48007;
assign x_48009 = x_48001 & x_48008;
assign x_48010 = x_47995 & x_48009;
assign x_48011 = x_16719 & x_16720;
assign x_48012 = x_16718 & x_48011;
assign x_48013 = x_16721 & x_16722;
assign x_48014 = x_16723 & x_16724;
assign x_48015 = x_48013 & x_48014;
assign x_48016 = x_48012 & x_48015;
assign x_48017 = x_16725 & x_16726;
assign x_48018 = x_16727 & x_16728;
assign x_48019 = x_48017 & x_48018;
assign x_48020 = x_16729 & x_16730;
assign x_48021 = x_16731 & x_16732;
assign x_48022 = x_48020 & x_48021;
assign x_48023 = x_48019 & x_48022;
assign x_48024 = x_48016 & x_48023;
assign x_48025 = x_16733 & x_16734;
assign x_48026 = x_16735 & x_16736;
assign x_48027 = x_48025 & x_48026;
assign x_48028 = x_16737 & x_16738;
assign x_48029 = x_16739 & x_16740;
assign x_48030 = x_48028 & x_48029;
assign x_48031 = x_48027 & x_48030;
assign x_48032 = x_16741 & x_16742;
assign x_48033 = x_16743 & x_16744;
assign x_48034 = x_48032 & x_48033;
assign x_48035 = x_16745 & x_16746;
assign x_48036 = x_16747 & x_16748;
assign x_48037 = x_48035 & x_48036;
assign x_48038 = x_48034 & x_48037;
assign x_48039 = x_48031 & x_48038;
assign x_48040 = x_48024 & x_48039;
assign x_48041 = x_48010 & x_48040;
assign x_48042 = x_47981 & x_48041;
assign x_48043 = x_16750 & x_16751;
assign x_48044 = x_16749 & x_48043;
assign x_48045 = x_16752 & x_16753;
assign x_48046 = x_16754 & x_16755;
assign x_48047 = x_48045 & x_48046;
assign x_48048 = x_48044 & x_48047;
assign x_48049 = x_16756 & x_16757;
assign x_48050 = x_16758 & x_16759;
assign x_48051 = x_48049 & x_48050;
assign x_48052 = x_16760 & x_16761;
assign x_48053 = x_16762 & x_16763;
assign x_48054 = x_48052 & x_48053;
assign x_48055 = x_48051 & x_48054;
assign x_48056 = x_48048 & x_48055;
assign x_48057 = x_16765 & x_16766;
assign x_48058 = x_16764 & x_48057;
assign x_48059 = x_16767 & x_16768;
assign x_48060 = x_16769 & x_16770;
assign x_48061 = x_48059 & x_48060;
assign x_48062 = x_48058 & x_48061;
assign x_48063 = x_16771 & x_16772;
assign x_48064 = x_16773 & x_16774;
assign x_48065 = x_48063 & x_48064;
assign x_48066 = x_16775 & x_16776;
assign x_48067 = x_16777 & x_16778;
assign x_48068 = x_48066 & x_48067;
assign x_48069 = x_48065 & x_48068;
assign x_48070 = x_48062 & x_48069;
assign x_48071 = x_48056 & x_48070;
assign x_48072 = x_16780 & x_16781;
assign x_48073 = x_16779 & x_48072;
assign x_48074 = x_16782 & x_16783;
assign x_48075 = x_16784 & x_16785;
assign x_48076 = x_48074 & x_48075;
assign x_48077 = x_48073 & x_48076;
assign x_48078 = x_16786 & x_16787;
assign x_48079 = x_16788 & x_16789;
assign x_48080 = x_48078 & x_48079;
assign x_48081 = x_16790 & x_16791;
assign x_48082 = x_16792 & x_16793;
assign x_48083 = x_48081 & x_48082;
assign x_48084 = x_48080 & x_48083;
assign x_48085 = x_48077 & x_48084;
assign x_48086 = x_16794 & x_16795;
assign x_48087 = x_16796 & x_16797;
assign x_48088 = x_48086 & x_48087;
assign x_48089 = x_16798 & x_16799;
assign x_48090 = x_16800 & x_16801;
assign x_48091 = x_48089 & x_48090;
assign x_48092 = x_48088 & x_48091;
assign x_48093 = x_16802 & x_16803;
assign x_48094 = x_16804 & x_16805;
assign x_48095 = x_48093 & x_48094;
assign x_48096 = x_16806 & x_16807;
assign x_48097 = x_16808 & x_16809;
assign x_48098 = x_48096 & x_48097;
assign x_48099 = x_48095 & x_48098;
assign x_48100 = x_48092 & x_48099;
assign x_48101 = x_48085 & x_48100;
assign x_48102 = x_48071 & x_48101;
assign x_48103 = x_16811 & x_16812;
assign x_48104 = x_16810 & x_48103;
assign x_48105 = x_16813 & x_16814;
assign x_48106 = x_16815 & x_16816;
assign x_48107 = x_48105 & x_48106;
assign x_48108 = x_48104 & x_48107;
assign x_48109 = x_16817 & x_16818;
assign x_48110 = x_16819 & x_16820;
assign x_48111 = x_48109 & x_48110;
assign x_48112 = x_16821 & x_16822;
assign x_48113 = x_16823 & x_16824;
assign x_48114 = x_48112 & x_48113;
assign x_48115 = x_48111 & x_48114;
assign x_48116 = x_48108 & x_48115;
assign x_48117 = x_16826 & x_16827;
assign x_48118 = x_16825 & x_48117;
assign x_48119 = x_16828 & x_16829;
assign x_48120 = x_16830 & x_16831;
assign x_48121 = x_48119 & x_48120;
assign x_48122 = x_48118 & x_48121;
assign x_48123 = x_16832 & x_16833;
assign x_48124 = x_16834 & x_16835;
assign x_48125 = x_48123 & x_48124;
assign x_48126 = x_16836 & x_16837;
assign x_48127 = x_16838 & x_16839;
assign x_48128 = x_48126 & x_48127;
assign x_48129 = x_48125 & x_48128;
assign x_48130 = x_48122 & x_48129;
assign x_48131 = x_48116 & x_48130;
assign x_48132 = x_16841 & x_16842;
assign x_48133 = x_16840 & x_48132;
assign x_48134 = x_16843 & x_16844;
assign x_48135 = x_16845 & x_16846;
assign x_48136 = x_48134 & x_48135;
assign x_48137 = x_48133 & x_48136;
assign x_48138 = x_16847 & x_16848;
assign x_48139 = x_16849 & x_16850;
assign x_48140 = x_48138 & x_48139;
assign x_48141 = x_16851 & x_16852;
assign x_48142 = x_16853 & x_16854;
assign x_48143 = x_48141 & x_48142;
assign x_48144 = x_48140 & x_48143;
assign x_48145 = x_48137 & x_48144;
assign x_48146 = x_16855 & x_16856;
assign x_48147 = x_16857 & x_16858;
assign x_48148 = x_48146 & x_48147;
assign x_48149 = x_16859 & x_16860;
assign x_48150 = x_16861 & x_16862;
assign x_48151 = x_48149 & x_48150;
assign x_48152 = x_48148 & x_48151;
assign x_48153 = x_16863 & x_16864;
assign x_48154 = x_16865 & x_16866;
assign x_48155 = x_48153 & x_48154;
assign x_48156 = x_16867 & x_16868;
assign x_48157 = x_16869 & x_16870;
assign x_48158 = x_48156 & x_48157;
assign x_48159 = x_48155 & x_48158;
assign x_48160 = x_48152 & x_48159;
assign x_48161 = x_48145 & x_48160;
assign x_48162 = x_48131 & x_48161;
assign x_48163 = x_48102 & x_48162;
assign x_48164 = x_48042 & x_48163;
assign x_48165 = x_16872 & x_16873;
assign x_48166 = x_16871 & x_48165;
assign x_48167 = x_16874 & x_16875;
assign x_48168 = x_16876 & x_16877;
assign x_48169 = x_48167 & x_48168;
assign x_48170 = x_48166 & x_48169;
assign x_48171 = x_16878 & x_16879;
assign x_48172 = x_16880 & x_16881;
assign x_48173 = x_48171 & x_48172;
assign x_48174 = x_16882 & x_16883;
assign x_48175 = x_16884 & x_16885;
assign x_48176 = x_48174 & x_48175;
assign x_48177 = x_48173 & x_48176;
assign x_48178 = x_48170 & x_48177;
assign x_48179 = x_16887 & x_16888;
assign x_48180 = x_16886 & x_48179;
assign x_48181 = x_16889 & x_16890;
assign x_48182 = x_16891 & x_16892;
assign x_48183 = x_48181 & x_48182;
assign x_48184 = x_48180 & x_48183;
assign x_48185 = x_16893 & x_16894;
assign x_48186 = x_16895 & x_16896;
assign x_48187 = x_48185 & x_48186;
assign x_48188 = x_16897 & x_16898;
assign x_48189 = x_16899 & x_16900;
assign x_48190 = x_48188 & x_48189;
assign x_48191 = x_48187 & x_48190;
assign x_48192 = x_48184 & x_48191;
assign x_48193 = x_48178 & x_48192;
assign x_48194 = x_16902 & x_16903;
assign x_48195 = x_16901 & x_48194;
assign x_48196 = x_16904 & x_16905;
assign x_48197 = x_16906 & x_16907;
assign x_48198 = x_48196 & x_48197;
assign x_48199 = x_48195 & x_48198;
assign x_48200 = x_16908 & x_16909;
assign x_48201 = x_16910 & x_16911;
assign x_48202 = x_48200 & x_48201;
assign x_48203 = x_16912 & x_16913;
assign x_48204 = x_16914 & x_16915;
assign x_48205 = x_48203 & x_48204;
assign x_48206 = x_48202 & x_48205;
assign x_48207 = x_48199 & x_48206;
assign x_48208 = x_16916 & x_16917;
assign x_48209 = x_16918 & x_16919;
assign x_48210 = x_48208 & x_48209;
assign x_48211 = x_16920 & x_16921;
assign x_48212 = x_16922 & x_16923;
assign x_48213 = x_48211 & x_48212;
assign x_48214 = x_48210 & x_48213;
assign x_48215 = x_16924 & x_16925;
assign x_48216 = x_16926 & x_16927;
assign x_48217 = x_48215 & x_48216;
assign x_48218 = x_16928 & x_16929;
assign x_48219 = x_16930 & x_16931;
assign x_48220 = x_48218 & x_48219;
assign x_48221 = x_48217 & x_48220;
assign x_48222 = x_48214 & x_48221;
assign x_48223 = x_48207 & x_48222;
assign x_48224 = x_48193 & x_48223;
assign x_48225 = x_16933 & x_16934;
assign x_48226 = x_16932 & x_48225;
assign x_48227 = x_16935 & x_16936;
assign x_48228 = x_16937 & x_16938;
assign x_48229 = x_48227 & x_48228;
assign x_48230 = x_48226 & x_48229;
assign x_48231 = x_16939 & x_16940;
assign x_48232 = x_16941 & x_16942;
assign x_48233 = x_48231 & x_48232;
assign x_48234 = x_16943 & x_16944;
assign x_48235 = x_16945 & x_16946;
assign x_48236 = x_48234 & x_48235;
assign x_48237 = x_48233 & x_48236;
assign x_48238 = x_48230 & x_48237;
assign x_48239 = x_16948 & x_16949;
assign x_48240 = x_16947 & x_48239;
assign x_48241 = x_16950 & x_16951;
assign x_48242 = x_16952 & x_16953;
assign x_48243 = x_48241 & x_48242;
assign x_48244 = x_48240 & x_48243;
assign x_48245 = x_16954 & x_16955;
assign x_48246 = x_16956 & x_16957;
assign x_48247 = x_48245 & x_48246;
assign x_48248 = x_16958 & x_16959;
assign x_48249 = x_16960 & x_16961;
assign x_48250 = x_48248 & x_48249;
assign x_48251 = x_48247 & x_48250;
assign x_48252 = x_48244 & x_48251;
assign x_48253 = x_48238 & x_48252;
assign x_48254 = x_16963 & x_16964;
assign x_48255 = x_16962 & x_48254;
assign x_48256 = x_16965 & x_16966;
assign x_48257 = x_16967 & x_16968;
assign x_48258 = x_48256 & x_48257;
assign x_48259 = x_48255 & x_48258;
assign x_48260 = x_16969 & x_16970;
assign x_48261 = x_16971 & x_16972;
assign x_48262 = x_48260 & x_48261;
assign x_48263 = x_16973 & x_16974;
assign x_48264 = x_16975 & x_16976;
assign x_48265 = x_48263 & x_48264;
assign x_48266 = x_48262 & x_48265;
assign x_48267 = x_48259 & x_48266;
assign x_48268 = x_16977 & x_16978;
assign x_48269 = x_16979 & x_16980;
assign x_48270 = x_48268 & x_48269;
assign x_48271 = x_16981 & x_16982;
assign x_48272 = x_16983 & x_16984;
assign x_48273 = x_48271 & x_48272;
assign x_48274 = x_48270 & x_48273;
assign x_48275 = x_16985 & x_16986;
assign x_48276 = x_16987 & x_16988;
assign x_48277 = x_48275 & x_48276;
assign x_48278 = x_16989 & x_16990;
assign x_48279 = x_16991 & x_16992;
assign x_48280 = x_48278 & x_48279;
assign x_48281 = x_48277 & x_48280;
assign x_48282 = x_48274 & x_48281;
assign x_48283 = x_48267 & x_48282;
assign x_48284 = x_48253 & x_48283;
assign x_48285 = x_48224 & x_48284;
assign x_48286 = x_16994 & x_16995;
assign x_48287 = x_16993 & x_48286;
assign x_48288 = x_16996 & x_16997;
assign x_48289 = x_16998 & x_16999;
assign x_48290 = x_48288 & x_48289;
assign x_48291 = x_48287 & x_48290;
assign x_48292 = x_17000 & x_17001;
assign x_48293 = x_17002 & x_17003;
assign x_48294 = x_48292 & x_48293;
assign x_48295 = x_17004 & x_17005;
assign x_48296 = x_17006 & x_17007;
assign x_48297 = x_48295 & x_48296;
assign x_48298 = x_48294 & x_48297;
assign x_48299 = x_48291 & x_48298;
assign x_48300 = x_17009 & x_17010;
assign x_48301 = x_17008 & x_48300;
assign x_48302 = x_17011 & x_17012;
assign x_48303 = x_17013 & x_17014;
assign x_48304 = x_48302 & x_48303;
assign x_48305 = x_48301 & x_48304;
assign x_48306 = x_17015 & x_17016;
assign x_48307 = x_17017 & x_17018;
assign x_48308 = x_48306 & x_48307;
assign x_48309 = x_17019 & x_17020;
assign x_48310 = x_17021 & x_17022;
assign x_48311 = x_48309 & x_48310;
assign x_48312 = x_48308 & x_48311;
assign x_48313 = x_48305 & x_48312;
assign x_48314 = x_48299 & x_48313;
assign x_48315 = x_17024 & x_17025;
assign x_48316 = x_17023 & x_48315;
assign x_48317 = x_17026 & x_17027;
assign x_48318 = x_17028 & x_17029;
assign x_48319 = x_48317 & x_48318;
assign x_48320 = x_48316 & x_48319;
assign x_48321 = x_17030 & x_17031;
assign x_48322 = x_17032 & x_17033;
assign x_48323 = x_48321 & x_48322;
assign x_48324 = x_17034 & x_17035;
assign x_48325 = x_17036 & x_17037;
assign x_48326 = x_48324 & x_48325;
assign x_48327 = x_48323 & x_48326;
assign x_48328 = x_48320 & x_48327;
assign x_48329 = x_17038 & x_17039;
assign x_48330 = x_17040 & x_17041;
assign x_48331 = x_48329 & x_48330;
assign x_48332 = x_17042 & x_17043;
assign x_48333 = x_17044 & x_17045;
assign x_48334 = x_48332 & x_48333;
assign x_48335 = x_48331 & x_48334;
assign x_48336 = x_17046 & x_17047;
assign x_48337 = x_17048 & x_17049;
assign x_48338 = x_48336 & x_48337;
assign x_48339 = x_17050 & x_17051;
assign x_48340 = x_17052 & x_17053;
assign x_48341 = x_48339 & x_48340;
assign x_48342 = x_48338 & x_48341;
assign x_48343 = x_48335 & x_48342;
assign x_48344 = x_48328 & x_48343;
assign x_48345 = x_48314 & x_48344;
assign x_48346 = x_17055 & x_17056;
assign x_48347 = x_17054 & x_48346;
assign x_48348 = x_17057 & x_17058;
assign x_48349 = x_17059 & x_17060;
assign x_48350 = x_48348 & x_48349;
assign x_48351 = x_48347 & x_48350;
assign x_48352 = x_17061 & x_17062;
assign x_48353 = x_17063 & x_17064;
assign x_48354 = x_48352 & x_48353;
assign x_48355 = x_17065 & x_17066;
assign x_48356 = x_17067 & x_17068;
assign x_48357 = x_48355 & x_48356;
assign x_48358 = x_48354 & x_48357;
assign x_48359 = x_48351 & x_48358;
assign x_48360 = x_17069 & x_17070;
assign x_48361 = x_17071 & x_17072;
assign x_48362 = x_48360 & x_48361;
assign x_48363 = x_17073 & x_17074;
assign x_48364 = x_17075 & x_17076;
assign x_48365 = x_48363 & x_48364;
assign x_48366 = x_48362 & x_48365;
assign x_48367 = x_17077 & x_17078;
assign x_48368 = x_17079 & x_17080;
assign x_48369 = x_48367 & x_48368;
assign x_48370 = x_17081 & x_17082;
assign x_48371 = x_17083 & x_17084;
assign x_48372 = x_48370 & x_48371;
assign x_48373 = x_48369 & x_48372;
assign x_48374 = x_48366 & x_48373;
assign x_48375 = x_48359 & x_48374;
assign x_48376 = x_17086 & x_17087;
assign x_48377 = x_17085 & x_48376;
assign x_48378 = x_17088 & x_17089;
assign x_48379 = x_17090 & x_17091;
assign x_48380 = x_48378 & x_48379;
assign x_48381 = x_48377 & x_48380;
assign x_48382 = x_17092 & x_17093;
assign x_48383 = x_17094 & x_17095;
assign x_48384 = x_48382 & x_48383;
assign x_48385 = x_17096 & x_17097;
assign x_48386 = x_17098 & x_17099;
assign x_48387 = x_48385 & x_48386;
assign x_48388 = x_48384 & x_48387;
assign x_48389 = x_48381 & x_48388;
assign x_48390 = x_17100 & x_17101;
assign x_48391 = x_17102 & x_17103;
assign x_48392 = x_48390 & x_48391;
assign x_48393 = x_17104 & x_17105;
assign x_48394 = x_17106 & x_17107;
assign x_48395 = x_48393 & x_48394;
assign x_48396 = x_48392 & x_48395;
assign x_48397 = x_17108 & x_17109;
assign x_48398 = x_17110 & x_17111;
assign x_48399 = x_48397 & x_48398;
assign x_48400 = x_17112 & x_17113;
assign x_48401 = x_17114 & x_17115;
assign x_48402 = x_48400 & x_48401;
assign x_48403 = x_48399 & x_48402;
assign x_48404 = x_48396 & x_48403;
assign x_48405 = x_48389 & x_48404;
assign x_48406 = x_48375 & x_48405;
assign x_48407 = x_48345 & x_48406;
assign x_48408 = x_48285 & x_48407;
assign x_48409 = x_48164 & x_48408;
assign x_48410 = x_17117 & x_17118;
assign x_48411 = x_17116 & x_48410;
assign x_48412 = x_17119 & x_17120;
assign x_48413 = x_17121 & x_17122;
assign x_48414 = x_48412 & x_48413;
assign x_48415 = x_48411 & x_48414;
assign x_48416 = x_17123 & x_17124;
assign x_48417 = x_17125 & x_17126;
assign x_48418 = x_48416 & x_48417;
assign x_48419 = x_17127 & x_17128;
assign x_48420 = x_17129 & x_17130;
assign x_48421 = x_48419 & x_48420;
assign x_48422 = x_48418 & x_48421;
assign x_48423 = x_48415 & x_48422;
assign x_48424 = x_17132 & x_17133;
assign x_48425 = x_17131 & x_48424;
assign x_48426 = x_17134 & x_17135;
assign x_48427 = x_17136 & x_17137;
assign x_48428 = x_48426 & x_48427;
assign x_48429 = x_48425 & x_48428;
assign x_48430 = x_17138 & x_17139;
assign x_48431 = x_17140 & x_17141;
assign x_48432 = x_48430 & x_48431;
assign x_48433 = x_17142 & x_17143;
assign x_48434 = x_17144 & x_17145;
assign x_48435 = x_48433 & x_48434;
assign x_48436 = x_48432 & x_48435;
assign x_48437 = x_48429 & x_48436;
assign x_48438 = x_48423 & x_48437;
assign x_48439 = x_17147 & x_17148;
assign x_48440 = x_17146 & x_48439;
assign x_48441 = x_17149 & x_17150;
assign x_48442 = x_17151 & x_17152;
assign x_48443 = x_48441 & x_48442;
assign x_48444 = x_48440 & x_48443;
assign x_48445 = x_17153 & x_17154;
assign x_48446 = x_17155 & x_17156;
assign x_48447 = x_48445 & x_48446;
assign x_48448 = x_17157 & x_17158;
assign x_48449 = x_17159 & x_17160;
assign x_48450 = x_48448 & x_48449;
assign x_48451 = x_48447 & x_48450;
assign x_48452 = x_48444 & x_48451;
assign x_48453 = x_17161 & x_17162;
assign x_48454 = x_17163 & x_17164;
assign x_48455 = x_48453 & x_48454;
assign x_48456 = x_17165 & x_17166;
assign x_48457 = x_17167 & x_17168;
assign x_48458 = x_48456 & x_48457;
assign x_48459 = x_48455 & x_48458;
assign x_48460 = x_17169 & x_17170;
assign x_48461 = x_17171 & x_17172;
assign x_48462 = x_48460 & x_48461;
assign x_48463 = x_17173 & x_17174;
assign x_48464 = x_17175 & x_17176;
assign x_48465 = x_48463 & x_48464;
assign x_48466 = x_48462 & x_48465;
assign x_48467 = x_48459 & x_48466;
assign x_48468 = x_48452 & x_48467;
assign x_48469 = x_48438 & x_48468;
assign x_48470 = x_17178 & x_17179;
assign x_48471 = x_17177 & x_48470;
assign x_48472 = x_17180 & x_17181;
assign x_48473 = x_17182 & x_17183;
assign x_48474 = x_48472 & x_48473;
assign x_48475 = x_48471 & x_48474;
assign x_48476 = x_17184 & x_17185;
assign x_48477 = x_17186 & x_17187;
assign x_48478 = x_48476 & x_48477;
assign x_48479 = x_17188 & x_17189;
assign x_48480 = x_17190 & x_17191;
assign x_48481 = x_48479 & x_48480;
assign x_48482 = x_48478 & x_48481;
assign x_48483 = x_48475 & x_48482;
assign x_48484 = x_17193 & x_17194;
assign x_48485 = x_17192 & x_48484;
assign x_48486 = x_17195 & x_17196;
assign x_48487 = x_17197 & x_17198;
assign x_48488 = x_48486 & x_48487;
assign x_48489 = x_48485 & x_48488;
assign x_48490 = x_17199 & x_17200;
assign x_48491 = x_17201 & x_17202;
assign x_48492 = x_48490 & x_48491;
assign x_48493 = x_17203 & x_17204;
assign x_48494 = x_17205 & x_17206;
assign x_48495 = x_48493 & x_48494;
assign x_48496 = x_48492 & x_48495;
assign x_48497 = x_48489 & x_48496;
assign x_48498 = x_48483 & x_48497;
assign x_48499 = x_17208 & x_17209;
assign x_48500 = x_17207 & x_48499;
assign x_48501 = x_17210 & x_17211;
assign x_48502 = x_17212 & x_17213;
assign x_48503 = x_48501 & x_48502;
assign x_48504 = x_48500 & x_48503;
assign x_48505 = x_17214 & x_17215;
assign x_48506 = x_17216 & x_17217;
assign x_48507 = x_48505 & x_48506;
assign x_48508 = x_17218 & x_17219;
assign x_48509 = x_17220 & x_17221;
assign x_48510 = x_48508 & x_48509;
assign x_48511 = x_48507 & x_48510;
assign x_48512 = x_48504 & x_48511;
assign x_48513 = x_17222 & x_17223;
assign x_48514 = x_17224 & x_17225;
assign x_48515 = x_48513 & x_48514;
assign x_48516 = x_17226 & x_17227;
assign x_48517 = x_17228 & x_17229;
assign x_48518 = x_48516 & x_48517;
assign x_48519 = x_48515 & x_48518;
assign x_48520 = x_17230 & x_17231;
assign x_48521 = x_17232 & x_17233;
assign x_48522 = x_48520 & x_48521;
assign x_48523 = x_17234 & x_17235;
assign x_48524 = x_17236 & x_17237;
assign x_48525 = x_48523 & x_48524;
assign x_48526 = x_48522 & x_48525;
assign x_48527 = x_48519 & x_48526;
assign x_48528 = x_48512 & x_48527;
assign x_48529 = x_48498 & x_48528;
assign x_48530 = x_48469 & x_48529;
assign x_48531 = x_17239 & x_17240;
assign x_48532 = x_17238 & x_48531;
assign x_48533 = x_17241 & x_17242;
assign x_48534 = x_17243 & x_17244;
assign x_48535 = x_48533 & x_48534;
assign x_48536 = x_48532 & x_48535;
assign x_48537 = x_17245 & x_17246;
assign x_48538 = x_17247 & x_17248;
assign x_48539 = x_48537 & x_48538;
assign x_48540 = x_17249 & x_17250;
assign x_48541 = x_17251 & x_17252;
assign x_48542 = x_48540 & x_48541;
assign x_48543 = x_48539 & x_48542;
assign x_48544 = x_48536 & x_48543;
assign x_48545 = x_17254 & x_17255;
assign x_48546 = x_17253 & x_48545;
assign x_48547 = x_17256 & x_17257;
assign x_48548 = x_17258 & x_17259;
assign x_48549 = x_48547 & x_48548;
assign x_48550 = x_48546 & x_48549;
assign x_48551 = x_17260 & x_17261;
assign x_48552 = x_17262 & x_17263;
assign x_48553 = x_48551 & x_48552;
assign x_48554 = x_17264 & x_17265;
assign x_48555 = x_17266 & x_17267;
assign x_48556 = x_48554 & x_48555;
assign x_48557 = x_48553 & x_48556;
assign x_48558 = x_48550 & x_48557;
assign x_48559 = x_48544 & x_48558;
assign x_48560 = x_17269 & x_17270;
assign x_48561 = x_17268 & x_48560;
assign x_48562 = x_17271 & x_17272;
assign x_48563 = x_17273 & x_17274;
assign x_48564 = x_48562 & x_48563;
assign x_48565 = x_48561 & x_48564;
assign x_48566 = x_17275 & x_17276;
assign x_48567 = x_17277 & x_17278;
assign x_48568 = x_48566 & x_48567;
assign x_48569 = x_17279 & x_17280;
assign x_48570 = x_17281 & x_17282;
assign x_48571 = x_48569 & x_48570;
assign x_48572 = x_48568 & x_48571;
assign x_48573 = x_48565 & x_48572;
assign x_48574 = x_17283 & x_17284;
assign x_48575 = x_17285 & x_17286;
assign x_48576 = x_48574 & x_48575;
assign x_48577 = x_17287 & x_17288;
assign x_48578 = x_17289 & x_17290;
assign x_48579 = x_48577 & x_48578;
assign x_48580 = x_48576 & x_48579;
assign x_48581 = x_17291 & x_17292;
assign x_48582 = x_17293 & x_17294;
assign x_48583 = x_48581 & x_48582;
assign x_48584 = x_17295 & x_17296;
assign x_48585 = x_17297 & x_17298;
assign x_48586 = x_48584 & x_48585;
assign x_48587 = x_48583 & x_48586;
assign x_48588 = x_48580 & x_48587;
assign x_48589 = x_48573 & x_48588;
assign x_48590 = x_48559 & x_48589;
assign x_48591 = x_17300 & x_17301;
assign x_48592 = x_17299 & x_48591;
assign x_48593 = x_17302 & x_17303;
assign x_48594 = x_17304 & x_17305;
assign x_48595 = x_48593 & x_48594;
assign x_48596 = x_48592 & x_48595;
assign x_48597 = x_17306 & x_17307;
assign x_48598 = x_17308 & x_17309;
assign x_48599 = x_48597 & x_48598;
assign x_48600 = x_17310 & x_17311;
assign x_48601 = x_17312 & x_17313;
assign x_48602 = x_48600 & x_48601;
assign x_48603 = x_48599 & x_48602;
assign x_48604 = x_48596 & x_48603;
assign x_48605 = x_17315 & x_17316;
assign x_48606 = x_17314 & x_48605;
assign x_48607 = x_17317 & x_17318;
assign x_48608 = x_17319 & x_17320;
assign x_48609 = x_48607 & x_48608;
assign x_48610 = x_48606 & x_48609;
assign x_48611 = x_17321 & x_17322;
assign x_48612 = x_17323 & x_17324;
assign x_48613 = x_48611 & x_48612;
assign x_48614 = x_17325 & x_17326;
assign x_48615 = x_17327 & x_17328;
assign x_48616 = x_48614 & x_48615;
assign x_48617 = x_48613 & x_48616;
assign x_48618 = x_48610 & x_48617;
assign x_48619 = x_48604 & x_48618;
assign x_48620 = x_17330 & x_17331;
assign x_48621 = x_17329 & x_48620;
assign x_48622 = x_17332 & x_17333;
assign x_48623 = x_17334 & x_17335;
assign x_48624 = x_48622 & x_48623;
assign x_48625 = x_48621 & x_48624;
assign x_48626 = x_17336 & x_17337;
assign x_48627 = x_17338 & x_17339;
assign x_48628 = x_48626 & x_48627;
assign x_48629 = x_17340 & x_17341;
assign x_48630 = x_17342 & x_17343;
assign x_48631 = x_48629 & x_48630;
assign x_48632 = x_48628 & x_48631;
assign x_48633 = x_48625 & x_48632;
assign x_48634 = x_17344 & x_17345;
assign x_48635 = x_17346 & x_17347;
assign x_48636 = x_48634 & x_48635;
assign x_48637 = x_17348 & x_17349;
assign x_48638 = x_17350 & x_17351;
assign x_48639 = x_48637 & x_48638;
assign x_48640 = x_48636 & x_48639;
assign x_48641 = x_17352 & x_17353;
assign x_48642 = x_17354 & x_17355;
assign x_48643 = x_48641 & x_48642;
assign x_48644 = x_17356 & x_17357;
assign x_48645 = x_17358 & x_17359;
assign x_48646 = x_48644 & x_48645;
assign x_48647 = x_48643 & x_48646;
assign x_48648 = x_48640 & x_48647;
assign x_48649 = x_48633 & x_48648;
assign x_48650 = x_48619 & x_48649;
assign x_48651 = x_48590 & x_48650;
assign x_48652 = x_48530 & x_48651;
assign x_48653 = x_17361 & x_17362;
assign x_48654 = x_17360 & x_48653;
assign x_48655 = x_17363 & x_17364;
assign x_48656 = x_17365 & x_17366;
assign x_48657 = x_48655 & x_48656;
assign x_48658 = x_48654 & x_48657;
assign x_48659 = x_17367 & x_17368;
assign x_48660 = x_17369 & x_17370;
assign x_48661 = x_48659 & x_48660;
assign x_48662 = x_17371 & x_17372;
assign x_48663 = x_17373 & x_17374;
assign x_48664 = x_48662 & x_48663;
assign x_48665 = x_48661 & x_48664;
assign x_48666 = x_48658 & x_48665;
assign x_48667 = x_17376 & x_17377;
assign x_48668 = x_17375 & x_48667;
assign x_48669 = x_17378 & x_17379;
assign x_48670 = x_17380 & x_17381;
assign x_48671 = x_48669 & x_48670;
assign x_48672 = x_48668 & x_48671;
assign x_48673 = x_17382 & x_17383;
assign x_48674 = x_17384 & x_17385;
assign x_48675 = x_48673 & x_48674;
assign x_48676 = x_17386 & x_17387;
assign x_48677 = x_17388 & x_17389;
assign x_48678 = x_48676 & x_48677;
assign x_48679 = x_48675 & x_48678;
assign x_48680 = x_48672 & x_48679;
assign x_48681 = x_48666 & x_48680;
assign x_48682 = x_17391 & x_17392;
assign x_48683 = x_17390 & x_48682;
assign x_48684 = x_17393 & x_17394;
assign x_48685 = x_17395 & x_17396;
assign x_48686 = x_48684 & x_48685;
assign x_48687 = x_48683 & x_48686;
assign x_48688 = x_17397 & x_17398;
assign x_48689 = x_17399 & x_17400;
assign x_48690 = x_48688 & x_48689;
assign x_48691 = x_17401 & x_17402;
assign x_48692 = x_17403 & x_17404;
assign x_48693 = x_48691 & x_48692;
assign x_48694 = x_48690 & x_48693;
assign x_48695 = x_48687 & x_48694;
assign x_48696 = x_17405 & x_17406;
assign x_48697 = x_17407 & x_17408;
assign x_48698 = x_48696 & x_48697;
assign x_48699 = x_17409 & x_17410;
assign x_48700 = x_17411 & x_17412;
assign x_48701 = x_48699 & x_48700;
assign x_48702 = x_48698 & x_48701;
assign x_48703 = x_17413 & x_17414;
assign x_48704 = x_17415 & x_17416;
assign x_48705 = x_48703 & x_48704;
assign x_48706 = x_17417 & x_17418;
assign x_48707 = x_17419 & x_17420;
assign x_48708 = x_48706 & x_48707;
assign x_48709 = x_48705 & x_48708;
assign x_48710 = x_48702 & x_48709;
assign x_48711 = x_48695 & x_48710;
assign x_48712 = x_48681 & x_48711;
assign x_48713 = x_17422 & x_17423;
assign x_48714 = x_17421 & x_48713;
assign x_48715 = x_17424 & x_17425;
assign x_48716 = x_17426 & x_17427;
assign x_48717 = x_48715 & x_48716;
assign x_48718 = x_48714 & x_48717;
assign x_48719 = x_17428 & x_17429;
assign x_48720 = x_17430 & x_17431;
assign x_48721 = x_48719 & x_48720;
assign x_48722 = x_17432 & x_17433;
assign x_48723 = x_17434 & x_17435;
assign x_48724 = x_48722 & x_48723;
assign x_48725 = x_48721 & x_48724;
assign x_48726 = x_48718 & x_48725;
assign x_48727 = x_17437 & x_17438;
assign x_48728 = x_17436 & x_48727;
assign x_48729 = x_17439 & x_17440;
assign x_48730 = x_17441 & x_17442;
assign x_48731 = x_48729 & x_48730;
assign x_48732 = x_48728 & x_48731;
assign x_48733 = x_17443 & x_17444;
assign x_48734 = x_17445 & x_17446;
assign x_48735 = x_48733 & x_48734;
assign x_48736 = x_17447 & x_17448;
assign x_48737 = x_17449 & x_17450;
assign x_48738 = x_48736 & x_48737;
assign x_48739 = x_48735 & x_48738;
assign x_48740 = x_48732 & x_48739;
assign x_48741 = x_48726 & x_48740;
assign x_48742 = x_17452 & x_17453;
assign x_48743 = x_17451 & x_48742;
assign x_48744 = x_17454 & x_17455;
assign x_48745 = x_17456 & x_17457;
assign x_48746 = x_48744 & x_48745;
assign x_48747 = x_48743 & x_48746;
assign x_48748 = x_17458 & x_17459;
assign x_48749 = x_17460 & x_17461;
assign x_48750 = x_48748 & x_48749;
assign x_48751 = x_17462 & x_17463;
assign x_48752 = x_17464 & x_17465;
assign x_48753 = x_48751 & x_48752;
assign x_48754 = x_48750 & x_48753;
assign x_48755 = x_48747 & x_48754;
assign x_48756 = x_17466 & x_17467;
assign x_48757 = x_17468 & x_17469;
assign x_48758 = x_48756 & x_48757;
assign x_48759 = x_17470 & x_17471;
assign x_48760 = x_17472 & x_17473;
assign x_48761 = x_48759 & x_48760;
assign x_48762 = x_48758 & x_48761;
assign x_48763 = x_17474 & x_17475;
assign x_48764 = x_17476 & x_17477;
assign x_48765 = x_48763 & x_48764;
assign x_48766 = x_17478 & x_17479;
assign x_48767 = x_17480 & x_17481;
assign x_48768 = x_48766 & x_48767;
assign x_48769 = x_48765 & x_48768;
assign x_48770 = x_48762 & x_48769;
assign x_48771 = x_48755 & x_48770;
assign x_48772 = x_48741 & x_48771;
assign x_48773 = x_48712 & x_48772;
assign x_48774 = x_17483 & x_17484;
assign x_48775 = x_17482 & x_48774;
assign x_48776 = x_17485 & x_17486;
assign x_48777 = x_17487 & x_17488;
assign x_48778 = x_48776 & x_48777;
assign x_48779 = x_48775 & x_48778;
assign x_48780 = x_17489 & x_17490;
assign x_48781 = x_17491 & x_17492;
assign x_48782 = x_48780 & x_48781;
assign x_48783 = x_17493 & x_17494;
assign x_48784 = x_17495 & x_17496;
assign x_48785 = x_48783 & x_48784;
assign x_48786 = x_48782 & x_48785;
assign x_48787 = x_48779 & x_48786;
assign x_48788 = x_17498 & x_17499;
assign x_48789 = x_17497 & x_48788;
assign x_48790 = x_17500 & x_17501;
assign x_48791 = x_17502 & x_17503;
assign x_48792 = x_48790 & x_48791;
assign x_48793 = x_48789 & x_48792;
assign x_48794 = x_17504 & x_17505;
assign x_48795 = x_17506 & x_17507;
assign x_48796 = x_48794 & x_48795;
assign x_48797 = x_17508 & x_17509;
assign x_48798 = x_17510 & x_17511;
assign x_48799 = x_48797 & x_48798;
assign x_48800 = x_48796 & x_48799;
assign x_48801 = x_48793 & x_48800;
assign x_48802 = x_48787 & x_48801;
assign x_48803 = x_17513 & x_17514;
assign x_48804 = x_17512 & x_48803;
assign x_48805 = x_17515 & x_17516;
assign x_48806 = x_17517 & x_17518;
assign x_48807 = x_48805 & x_48806;
assign x_48808 = x_48804 & x_48807;
assign x_48809 = x_17519 & x_17520;
assign x_48810 = x_17521 & x_17522;
assign x_48811 = x_48809 & x_48810;
assign x_48812 = x_17523 & x_17524;
assign x_48813 = x_17525 & x_17526;
assign x_48814 = x_48812 & x_48813;
assign x_48815 = x_48811 & x_48814;
assign x_48816 = x_48808 & x_48815;
assign x_48817 = x_17527 & x_17528;
assign x_48818 = x_17529 & x_17530;
assign x_48819 = x_48817 & x_48818;
assign x_48820 = x_17531 & x_17532;
assign x_48821 = x_17533 & x_17534;
assign x_48822 = x_48820 & x_48821;
assign x_48823 = x_48819 & x_48822;
assign x_48824 = x_17535 & x_17536;
assign x_48825 = x_17537 & x_17538;
assign x_48826 = x_48824 & x_48825;
assign x_48827 = x_17539 & x_17540;
assign x_48828 = x_17541 & x_17542;
assign x_48829 = x_48827 & x_48828;
assign x_48830 = x_48826 & x_48829;
assign x_48831 = x_48823 & x_48830;
assign x_48832 = x_48816 & x_48831;
assign x_48833 = x_48802 & x_48832;
assign x_48834 = x_17544 & x_17545;
assign x_48835 = x_17543 & x_48834;
assign x_48836 = x_17546 & x_17547;
assign x_48837 = x_17548 & x_17549;
assign x_48838 = x_48836 & x_48837;
assign x_48839 = x_48835 & x_48838;
assign x_48840 = x_17550 & x_17551;
assign x_48841 = x_17552 & x_17553;
assign x_48842 = x_48840 & x_48841;
assign x_48843 = x_17554 & x_17555;
assign x_48844 = x_17556 & x_17557;
assign x_48845 = x_48843 & x_48844;
assign x_48846 = x_48842 & x_48845;
assign x_48847 = x_48839 & x_48846;
assign x_48848 = x_17558 & x_17559;
assign x_48849 = x_17560 & x_17561;
assign x_48850 = x_48848 & x_48849;
assign x_48851 = x_17562 & x_17563;
assign x_48852 = x_17564 & x_17565;
assign x_48853 = x_48851 & x_48852;
assign x_48854 = x_48850 & x_48853;
assign x_48855 = x_17566 & x_17567;
assign x_48856 = x_17568 & x_17569;
assign x_48857 = x_48855 & x_48856;
assign x_48858 = x_17570 & x_17571;
assign x_48859 = x_17572 & x_17573;
assign x_48860 = x_48858 & x_48859;
assign x_48861 = x_48857 & x_48860;
assign x_48862 = x_48854 & x_48861;
assign x_48863 = x_48847 & x_48862;
assign x_48864 = x_17575 & x_17576;
assign x_48865 = x_17574 & x_48864;
assign x_48866 = x_17577 & x_17578;
assign x_48867 = x_17579 & x_17580;
assign x_48868 = x_48866 & x_48867;
assign x_48869 = x_48865 & x_48868;
assign x_48870 = x_17581 & x_17582;
assign x_48871 = x_17583 & x_17584;
assign x_48872 = x_48870 & x_48871;
assign x_48873 = x_17585 & x_17586;
assign x_48874 = x_17587 & x_17588;
assign x_48875 = x_48873 & x_48874;
assign x_48876 = x_48872 & x_48875;
assign x_48877 = x_48869 & x_48876;
assign x_48878 = x_17589 & x_17590;
assign x_48879 = x_17591 & x_17592;
assign x_48880 = x_48878 & x_48879;
assign x_48881 = x_17593 & x_17594;
assign x_48882 = x_17595 & x_17596;
assign x_48883 = x_48881 & x_48882;
assign x_48884 = x_48880 & x_48883;
assign x_48885 = x_17597 & x_17598;
assign x_48886 = x_17599 & x_17600;
assign x_48887 = x_48885 & x_48886;
assign x_48888 = x_17601 & x_17602;
assign x_48889 = x_17603 & x_17604;
assign x_48890 = x_48888 & x_48889;
assign x_48891 = x_48887 & x_48890;
assign x_48892 = x_48884 & x_48891;
assign x_48893 = x_48877 & x_48892;
assign x_48894 = x_48863 & x_48893;
assign x_48895 = x_48833 & x_48894;
assign x_48896 = x_48773 & x_48895;
assign x_48897 = x_48652 & x_48896;
assign x_48898 = x_48409 & x_48897;
assign x_48899 = x_47921 & x_48898;
assign x_48900 = x_17606 & x_17607;
assign x_48901 = x_17605 & x_48900;
assign x_48902 = x_17608 & x_17609;
assign x_48903 = x_17610 & x_17611;
assign x_48904 = x_48902 & x_48903;
assign x_48905 = x_48901 & x_48904;
assign x_48906 = x_17612 & x_17613;
assign x_48907 = x_17614 & x_17615;
assign x_48908 = x_48906 & x_48907;
assign x_48909 = x_17616 & x_17617;
assign x_48910 = x_17618 & x_17619;
assign x_48911 = x_48909 & x_48910;
assign x_48912 = x_48908 & x_48911;
assign x_48913 = x_48905 & x_48912;
assign x_48914 = x_17621 & x_17622;
assign x_48915 = x_17620 & x_48914;
assign x_48916 = x_17623 & x_17624;
assign x_48917 = x_17625 & x_17626;
assign x_48918 = x_48916 & x_48917;
assign x_48919 = x_48915 & x_48918;
assign x_48920 = x_17627 & x_17628;
assign x_48921 = x_17629 & x_17630;
assign x_48922 = x_48920 & x_48921;
assign x_48923 = x_17631 & x_17632;
assign x_48924 = x_17633 & x_17634;
assign x_48925 = x_48923 & x_48924;
assign x_48926 = x_48922 & x_48925;
assign x_48927 = x_48919 & x_48926;
assign x_48928 = x_48913 & x_48927;
assign x_48929 = x_17636 & x_17637;
assign x_48930 = x_17635 & x_48929;
assign x_48931 = x_17638 & x_17639;
assign x_48932 = x_17640 & x_17641;
assign x_48933 = x_48931 & x_48932;
assign x_48934 = x_48930 & x_48933;
assign x_48935 = x_17642 & x_17643;
assign x_48936 = x_17644 & x_17645;
assign x_48937 = x_48935 & x_48936;
assign x_48938 = x_17646 & x_17647;
assign x_48939 = x_17648 & x_17649;
assign x_48940 = x_48938 & x_48939;
assign x_48941 = x_48937 & x_48940;
assign x_48942 = x_48934 & x_48941;
assign x_48943 = x_17650 & x_17651;
assign x_48944 = x_17652 & x_17653;
assign x_48945 = x_48943 & x_48944;
assign x_48946 = x_17654 & x_17655;
assign x_48947 = x_17656 & x_17657;
assign x_48948 = x_48946 & x_48947;
assign x_48949 = x_48945 & x_48948;
assign x_48950 = x_17658 & x_17659;
assign x_48951 = x_17660 & x_17661;
assign x_48952 = x_48950 & x_48951;
assign x_48953 = x_17662 & x_17663;
assign x_48954 = x_17664 & x_17665;
assign x_48955 = x_48953 & x_48954;
assign x_48956 = x_48952 & x_48955;
assign x_48957 = x_48949 & x_48956;
assign x_48958 = x_48942 & x_48957;
assign x_48959 = x_48928 & x_48958;
assign x_48960 = x_17667 & x_17668;
assign x_48961 = x_17666 & x_48960;
assign x_48962 = x_17669 & x_17670;
assign x_48963 = x_17671 & x_17672;
assign x_48964 = x_48962 & x_48963;
assign x_48965 = x_48961 & x_48964;
assign x_48966 = x_17673 & x_17674;
assign x_48967 = x_17675 & x_17676;
assign x_48968 = x_48966 & x_48967;
assign x_48969 = x_17677 & x_17678;
assign x_48970 = x_17679 & x_17680;
assign x_48971 = x_48969 & x_48970;
assign x_48972 = x_48968 & x_48971;
assign x_48973 = x_48965 & x_48972;
assign x_48974 = x_17682 & x_17683;
assign x_48975 = x_17681 & x_48974;
assign x_48976 = x_17684 & x_17685;
assign x_48977 = x_17686 & x_17687;
assign x_48978 = x_48976 & x_48977;
assign x_48979 = x_48975 & x_48978;
assign x_48980 = x_17688 & x_17689;
assign x_48981 = x_17690 & x_17691;
assign x_48982 = x_48980 & x_48981;
assign x_48983 = x_17692 & x_17693;
assign x_48984 = x_17694 & x_17695;
assign x_48985 = x_48983 & x_48984;
assign x_48986 = x_48982 & x_48985;
assign x_48987 = x_48979 & x_48986;
assign x_48988 = x_48973 & x_48987;
assign x_48989 = x_17697 & x_17698;
assign x_48990 = x_17696 & x_48989;
assign x_48991 = x_17699 & x_17700;
assign x_48992 = x_17701 & x_17702;
assign x_48993 = x_48991 & x_48992;
assign x_48994 = x_48990 & x_48993;
assign x_48995 = x_17703 & x_17704;
assign x_48996 = x_17705 & x_17706;
assign x_48997 = x_48995 & x_48996;
assign x_48998 = x_17707 & x_17708;
assign x_48999 = x_17709 & x_17710;
assign x_49000 = x_48998 & x_48999;
assign x_49001 = x_48997 & x_49000;
assign x_49002 = x_48994 & x_49001;
assign x_49003 = x_17711 & x_17712;
assign x_49004 = x_17713 & x_17714;
assign x_49005 = x_49003 & x_49004;
assign x_49006 = x_17715 & x_17716;
assign x_49007 = x_17717 & x_17718;
assign x_49008 = x_49006 & x_49007;
assign x_49009 = x_49005 & x_49008;
assign x_49010 = x_17719 & x_17720;
assign x_49011 = x_17721 & x_17722;
assign x_49012 = x_49010 & x_49011;
assign x_49013 = x_17723 & x_17724;
assign x_49014 = x_17725 & x_17726;
assign x_49015 = x_49013 & x_49014;
assign x_49016 = x_49012 & x_49015;
assign x_49017 = x_49009 & x_49016;
assign x_49018 = x_49002 & x_49017;
assign x_49019 = x_48988 & x_49018;
assign x_49020 = x_48959 & x_49019;
assign x_49021 = x_17728 & x_17729;
assign x_49022 = x_17727 & x_49021;
assign x_49023 = x_17730 & x_17731;
assign x_49024 = x_17732 & x_17733;
assign x_49025 = x_49023 & x_49024;
assign x_49026 = x_49022 & x_49025;
assign x_49027 = x_17734 & x_17735;
assign x_49028 = x_17736 & x_17737;
assign x_49029 = x_49027 & x_49028;
assign x_49030 = x_17738 & x_17739;
assign x_49031 = x_17740 & x_17741;
assign x_49032 = x_49030 & x_49031;
assign x_49033 = x_49029 & x_49032;
assign x_49034 = x_49026 & x_49033;
assign x_49035 = x_17743 & x_17744;
assign x_49036 = x_17742 & x_49035;
assign x_49037 = x_17745 & x_17746;
assign x_49038 = x_17747 & x_17748;
assign x_49039 = x_49037 & x_49038;
assign x_49040 = x_49036 & x_49039;
assign x_49041 = x_17749 & x_17750;
assign x_49042 = x_17751 & x_17752;
assign x_49043 = x_49041 & x_49042;
assign x_49044 = x_17753 & x_17754;
assign x_49045 = x_17755 & x_17756;
assign x_49046 = x_49044 & x_49045;
assign x_49047 = x_49043 & x_49046;
assign x_49048 = x_49040 & x_49047;
assign x_49049 = x_49034 & x_49048;
assign x_49050 = x_17758 & x_17759;
assign x_49051 = x_17757 & x_49050;
assign x_49052 = x_17760 & x_17761;
assign x_49053 = x_17762 & x_17763;
assign x_49054 = x_49052 & x_49053;
assign x_49055 = x_49051 & x_49054;
assign x_49056 = x_17764 & x_17765;
assign x_49057 = x_17766 & x_17767;
assign x_49058 = x_49056 & x_49057;
assign x_49059 = x_17768 & x_17769;
assign x_49060 = x_17770 & x_17771;
assign x_49061 = x_49059 & x_49060;
assign x_49062 = x_49058 & x_49061;
assign x_49063 = x_49055 & x_49062;
assign x_49064 = x_17772 & x_17773;
assign x_49065 = x_17774 & x_17775;
assign x_49066 = x_49064 & x_49065;
assign x_49067 = x_17776 & x_17777;
assign x_49068 = x_17778 & x_17779;
assign x_49069 = x_49067 & x_49068;
assign x_49070 = x_49066 & x_49069;
assign x_49071 = x_17780 & x_17781;
assign x_49072 = x_17782 & x_17783;
assign x_49073 = x_49071 & x_49072;
assign x_49074 = x_17784 & x_17785;
assign x_49075 = x_17786 & x_17787;
assign x_49076 = x_49074 & x_49075;
assign x_49077 = x_49073 & x_49076;
assign x_49078 = x_49070 & x_49077;
assign x_49079 = x_49063 & x_49078;
assign x_49080 = x_49049 & x_49079;
assign x_49081 = x_17789 & x_17790;
assign x_49082 = x_17788 & x_49081;
assign x_49083 = x_17791 & x_17792;
assign x_49084 = x_17793 & x_17794;
assign x_49085 = x_49083 & x_49084;
assign x_49086 = x_49082 & x_49085;
assign x_49087 = x_17795 & x_17796;
assign x_49088 = x_17797 & x_17798;
assign x_49089 = x_49087 & x_49088;
assign x_49090 = x_17799 & x_17800;
assign x_49091 = x_17801 & x_17802;
assign x_49092 = x_49090 & x_49091;
assign x_49093 = x_49089 & x_49092;
assign x_49094 = x_49086 & x_49093;
assign x_49095 = x_17804 & x_17805;
assign x_49096 = x_17803 & x_49095;
assign x_49097 = x_17806 & x_17807;
assign x_49098 = x_17808 & x_17809;
assign x_49099 = x_49097 & x_49098;
assign x_49100 = x_49096 & x_49099;
assign x_49101 = x_17810 & x_17811;
assign x_49102 = x_17812 & x_17813;
assign x_49103 = x_49101 & x_49102;
assign x_49104 = x_17814 & x_17815;
assign x_49105 = x_17816 & x_17817;
assign x_49106 = x_49104 & x_49105;
assign x_49107 = x_49103 & x_49106;
assign x_49108 = x_49100 & x_49107;
assign x_49109 = x_49094 & x_49108;
assign x_49110 = x_17819 & x_17820;
assign x_49111 = x_17818 & x_49110;
assign x_49112 = x_17821 & x_17822;
assign x_49113 = x_17823 & x_17824;
assign x_49114 = x_49112 & x_49113;
assign x_49115 = x_49111 & x_49114;
assign x_49116 = x_17825 & x_17826;
assign x_49117 = x_17827 & x_17828;
assign x_49118 = x_49116 & x_49117;
assign x_49119 = x_17829 & x_17830;
assign x_49120 = x_17831 & x_17832;
assign x_49121 = x_49119 & x_49120;
assign x_49122 = x_49118 & x_49121;
assign x_49123 = x_49115 & x_49122;
assign x_49124 = x_17833 & x_17834;
assign x_49125 = x_17835 & x_17836;
assign x_49126 = x_49124 & x_49125;
assign x_49127 = x_17837 & x_17838;
assign x_49128 = x_17839 & x_17840;
assign x_49129 = x_49127 & x_49128;
assign x_49130 = x_49126 & x_49129;
assign x_49131 = x_17841 & x_17842;
assign x_49132 = x_17843 & x_17844;
assign x_49133 = x_49131 & x_49132;
assign x_49134 = x_17845 & x_17846;
assign x_49135 = x_17847 & x_17848;
assign x_49136 = x_49134 & x_49135;
assign x_49137 = x_49133 & x_49136;
assign x_49138 = x_49130 & x_49137;
assign x_49139 = x_49123 & x_49138;
assign x_49140 = x_49109 & x_49139;
assign x_49141 = x_49080 & x_49140;
assign x_49142 = x_49020 & x_49141;
assign x_49143 = x_17850 & x_17851;
assign x_49144 = x_17849 & x_49143;
assign x_49145 = x_17852 & x_17853;
assign x_49146 = x_17854 & x_17855;
assign x_49147 = x_49145 & x_49146;
assign x_49148 = x_49144 & x_49147;
assign x_49149 = x_17856 & x_17857;
assign x_49150 = x_17858 & x_17859;
assign x_49151 = x_49149 & x_49150;
assign x_49152 = x_17860 & x_17861;
assign x_49153 = x_17862 & x_17863;
assign x_49154 = x_49152 & x_49153;
assign x_49155 = x_49151 & x_49154;
assign x_49156 = x_49148 & x_49155;
assign x_49157 = x_17865 & x_17866;
assign x_49158 = x_17864 & x_49157;
assign x_49159 = x_17867 & x_17868;
assign x_49160 = x_17869 & x_17870;
assign x_49161 = x_49159 & x_49160;
assign x_49162 = x_49158 & x_49161;
assign x_49163 = x_17871 & x_17872;
assign x_49164 = x_17873 & x_17874;
assign x_49165 = x_49163 & x_49164;
assign x_49166 = x_17875 & x_17876;
assign x_49167 = x_17877 & x_17878;
assign x_49168 = x_49166 & x_49167;
assign x_49169 = x_49165 & x_49168;
assign x_49170 = x_49162 & x_49169;
assign x_49171 = x_49156 & x_49170;
assign x_49172 = x_17880 & x_17881;
assign x_49173 = x_17879 & x_49172;
assign x_49174 = x_17882 & x_17883;
assign x_49175 = x_17884 & x_17885;
assign x_49176 = x_49174 & x_49175;
assign x_49177 = x_49173 & x_49176;
assign x_49178 = x_17886 & x_17887;
assign x_49179 = x_17888 & x_17889;
assign x_49180 = x_49178 & x_49179;
assign x_49181 = x_17890 & x_17891;
assign x_49182 = x_17892 & x_17893;
assign x_49183 = x_49181 & x_49182;
assign x_49184 = x_49180 & x_49183;
assign x_49185 = x_49177 & x_49184;
assign x_49186 = x_17894 & x_17895;
assign x_49187 = x_17896 & x_17897;
assign x_49188 = x_49186 & x_49187;
assign x_49189 = x_17898 & x_17899;
assign x_49190 = x_17900 & x_17901;
assign x_49191 = x_49189 & x_49190;
assign x_49192 = x_49188 & x_49191;
assign x_49193 = x_17902 & x_17903;
assign x_49194 = x_17904 & x_17905;
assign x_49195 = x_49193 & x_49194;
assign x_49196 = x_17906 & x_17907;
assign x_49197 = x_17908 & x_17909;
assign x_49198 = x_49196 & x_49197;
assign x_49199 = x_49195 & x_49198;
assign x_49200 = x_49192 & x_49199;
assign x_49201 = x_49185 & x_49200;
assign x_49202 = x_49171 & x_49201;
assign x_49203 = x_17911 & x_17912;
assign x_49204 = x_17910 & x_49203;
assign x_49205 = x_17913 & x_17914;
assign x_49206 = x_17915 & x_17916;
assign x_49207 = x_49205 & x_49206;
assign x_49208 = x_49204 & x_49207;
assign x_49209 = x_17917 & x_17918;
assign x_49210 = x_17919 & x_17920;
assign x_49211 = x_49209 & x_49210;
assign x_49212 = x_17921 & x_17922;
assign x_49213 = x_17923 & x_17924;
assign x_49214 = x_49212 & x_49213;
assign x_49215 = x_49211 & x_49214;
assign x_49216 = x_49208 & x_49215;
assign x_49217 = x_17926 & x_17927;
assign x_49218 = x_17925 & x_49217;
assign x_49219 = x_17928 & x_17929;
assign x_49220 = x_17930 & x_17931;
assign x_49221 = x_49219 & x_49220;
assign x_49222 = x_49218 & x_49221;
assign x_49223 = x_17932 & x_17933;
assign x_49224 = x_17934 & x_17935;
assign x_49225 = x_49223 & x_49224;
assign x_49226 = x_17936 & x_17937;
assign x_49227 = x_17938 & x_17939;
assign x_49228 = x_49226 & x_49227;
assign x_49229 = x_49225 & x_49228;
assign x_49230 = x_49222 & x_49229;
assign x_49231 = x_49216 & x_49230;
assign x_49232 = x_17941 & x_17942;
assign x_49233 = x_17940 & x_49232;
assign x_49234 = x_17943 & x_17944;
assign x_49235 = x_17945 & x_17946;
assign x_49236 = x_49234 & x_49235;
assign x_49237 = x_49233 & x_49236;
assign x_49238 = x_17947 & x_17948;
assign x_49239 = x_17949 & x_17950;
assign x_49240 = x_49238 & x_49239;
assign x_49241 = x_17951 & x_17952;
assign x_49242 = x_17953 & x_17954;
assign x_49243 = x_49241 & x_49242;
assign x_49244 = x_49240 & x_49243;
assign x_49245 = x_49237 & x_49244;
assign x_49246 = x_17955 & x_17956;
assign x_49247 = x_17957 & x_17958;
assign x_49248 = x_49246 & x_49247;
assign x_49249 = x_17959 & x_17960;
assign x_49250 = x_17961 & x_17962;
assign x_49251 = x_49249 & x_49250;
assign x_49252 = x_49248 & x_49251;
assign x_49253 = x_17963 & x_17964;
assign x_49254 = x_17965 & x_17966;
assign x_49255 = x_49253 & x_49254;
assign x_49256 = x_17967 & x_17968;
assign x_49257 = x_17969 & x_17970;
assign x_49258 = x_49256 & x_49257;
assign x_49259 = x_49255 & x_49258;
assign x_49260 = x_49252 & x_49259;
assign x_49261 = x_49245 & x_49260;
assign x_49262 = x_49231 & x_49261;
assign x_49263 = x_49202 & x_49262;
assign x_49264 = x_17972 & x_17973;
assign x_49265 = x_17971 & x_49264;
assign x_49266 = x_17974 & x_17975;
assign x_49267 = x_17976 & x_17977;
assign x_49268 = x_49266 & x_49267;
assign x_49269 = x_49265 & x_49268;
assign x_49270 = x_17978 & x_17979;
assign x_49271 = x_17980 & x_17981;
assign x_49272 = x_49270 & x_49271;
assign x_49273 = x_17982 & x_17983;
assign x_49274 = x_17984 & x_17985;
assign x_49275 = x_49273 & x_49274;
assign x_49276 = x_49272 & x_49275;
assign x_49277 = x_49269 & x_49276;
assign x_49278 = x_17987 & x_17988;
assign x_49279 = x_17986 & x_49278;
assign x_49280 = x_17989 & x_17990;
assign x_49281 = x_17991 & x_17992;
assign x_49282 = x_49280 & x_49281;
assign x_49283 = x_49279 & x_49282;
assign x_49284 = x_17993 & x_17994;
assign x_49285 = x_17995 & x_17996;
assign x_49286 = x_49284 & x_49285;
assign x_49287 = x_17997 & x_17998;
assign x_49288 = x_17999 & x_18000;
assign x_49289 = x_49287 & x_49288;
assign x_49290 = x_49286 & x_49289;
assign x_49291 = x_49283 & x_49290;
assign x_49292 = x_49277 & x_49291;
assign x_49293 = x_18002 & x_18003;
assign x_49294 = x_18001 & x_49293;
assign x_49295 = x_18004 & x_18005;
assign x_49296 = x_18006 & x_18007;
assign x_49297 = x_49295 & x_49296;
assign x_49298 = x_49294 & x_49297;
assign x_49299 = x_18008 & x_18009;
assign x_49300 = x_18010 & x_18011;
assign x_49301 = x_49299 & x_49300;
assign x_49302 = x_18012 & x_18013;
assign x_49303 = x_18014 & x_18015;
assign x_49304 = x_49302 & x_49303;
assign x_49305 = x_49301 & x_49304;
assign x_49306 = x_49298 & x_49305;
assign x_49307 = x_18016 & x_18017;
assign x_49308 = x_18018 & x_18019;
assign x_49309 = x_49307 & x_49308;
assign x_49310 = x_18020 & x_18021;
assign x_49311 = x_18022 & x_18023;
assign x_49312 = x_49310 & x_49311;
assign x_49313 = x_49309 & x_49312;
assign x_49314 = x_18024 & x_18025;
assign x_49315 = x_18026 & x_18027;
assign x_49316 = x_49314 & x_49315;
assign x_49317 = x_18028 & x_18029;
assign x_49318 = x_18030 & x_18031;
assign x_49319 = x_49317 & x_49318;
assign x_49320 = x_49316 & x_49319;
assign x_49321 = x_49313 & x_49320;
assign x_49322 = x_49306 & x_49321;
assign x_49323 = x_49292 & x_49322;
assign x_49324 = x_18033 & x_18034;
assign x_49325 = x_18032 & x_49324;
assign x_49326 = x_18035 & x_18036;
assign x_49327 = x_18037 & x_18038;
assign x_49328 = x_49326 & x_49327;
assign x_49329 = x_49325 & x_49328;
assign x_49330 = x_18039 & x_18040;
assign x_49331 = x_18041 & x_18042;
assign x_49332 = x_49330 & x_49331;
assign x_49333 = x_18043 & x_18044;
assign x_49334 = x_18045 & x_18046;
assign x_49335 = x_49333 & x_49334;
assign x_49336 = x_49332 & x_49335;
assign x_49337 = x_49329 & x_49336;
assign x_49338 = x_18047 & x_18048;
assign x_49339 = x_18049 & x_18050;
assign x_49340 = x_49338 & x_49339;
assign x_49341 = x_18051 & x_18052;
assign x_49342 = x_18053 & x_18054;
assign x_49343 = x_49341 & x_49342;
assign x_49344 = x_49340 & x_49343;
assign x_49345 = x_18055 & x_18056;
assign x_49346 = x_18057 & x_18058;
assign x_49347 = x_49345 & x_49346;
assign x_49348 = x_18059 & x_18060;
assign x_49349 = x_18061 & x_18062;
assign x_49350 = x_49348 & x_49349;
assign x_49351 = x_49347 & x_49350;
assign x_49352 = x_49344 & x_49351;
assign x_49353 = x_49337 & x_49352;
assign x_49354 = x_18064 & x_18065;
assign x_49355 = x_18063 & x_49354;
assign x_49356 = x_18066 & x_18067;
assign x_49357 = x_18068 & x_18069;
assign x_49358 = x_49356 & x_49357;
assign x_49359 = x_49355 & x_49358;
assign x_49360 = x_18070 & x_18071;
assign x_49361 = x_18072 & x_18073;
assign x_49362 = x_49360 & x_49361;
assign x_49363 = x_18074 & x_18075;
assign x_49364 = x_18076 & x_18077;
assign x_49365 = x_49363 & x_49364;
assign x_49366 = x_49362 & x_49365;
assign x_49367 = x_49359 & x_49366;
assign x_49368 = x_18078 & x_18079;
assign x_49369 = x_18080 & x_18081;
assign x_49370 = x_49368 & x_49369;
assign x_49371 = x_18082 & x_18083;
assign x_49372 = x_18084 & x_18085;
assign x_49373 = x_49371 & x_49372;
assign x_49374 = x_49370 & x_49373;
assign x_49375 = x_18086 & x_18087;
assign x_49376 = x_18088 & x_18089;
assign x_49377 = x_49375 & x_49376;
assign x_49378 = x_18090 & x_18091;
assign x_49379 = x_18092 & x_18093;
assign x_49380 = x_49378 & x_49379;
assign x_49381 = x_49377 & x_49380;
assign x_49382 = x_49374 & x_49381;
assign x_49383 = x_49367 & x_49382;
assign x_49384 = x_49353 & x_49383;
assign x_49385 = x_49323 & x_49384;
assign x_49386 = x_49263 & x_49385;
assign x_49387 = x_49142 & x_49386;
assign x_49388 = x_18095 & x_18096;
assign x_49389 = x_18094 & x_49388;
assign x_49390 = x_18097 & x_18098;
assign x_49391 = x_18099 & x_18100;
assign x_49392 = x_49390 & x_49391;
assign x_49393 = x_49389 & x_49392;
assign x_49394 = x_18101 & x_18102;
assign x_49395 = x_18103 & x_18104;
assign x_49396 = x_49394 & x_49395;
assign x_49397 = x_18105 & x_18106;
assign x_49398 = x_18107 & x_18108;
assign x_49399 = x_49397 & x_49398;
assign x_49400 = x_49396 & x_49399;
assign x_49401 = x_49393 & x_49400;
assign x_49402 = x_18110 & x_18111;
assign x_49403 = x_18109 & x_49402;
assign x_49404 = x_18112 & x_18113;
assign x_49405 = x_18114 & x_18115;
assign x_49406 = x_49404 & x_49405;
assign x_49407 = x_49403 & x_49406;
assign x_49408 = x_18116 & x_18117;
assign x_49409 = x_18118 & x_18119;
assign x_49410 = x_49408 & x_49409;
assign x_49411 = x_18120 & x_18121;
assign x_49412 = x_18122 & x_18123;
assign x_49413 = x_49411 & x_49412;
assign x_49414 = x_49410 & x_49413;
assign x_49415 = x_49407 & x_49414;
assign x_49416 = x_49401 & x_49415;
assign x_49417 = x_18125 & x_18126;
assign x_49418 = x_18124 & x_49417;
assign x_49419 = x_18127 & x_18128;
assign x_49420 = x_18129 & x_18130;
assign x_49421 = x_49419 & x_49420;
assign x_49422 = x_49418 & x_49421;
assign x_49423 = x_18131 & x_18132;
assign x_49424 = x_18133 & x_18134;
assign x_49425 = x_49423 & x_49424;
assign x_49426 = x_18135 & x_18136;
assign x_49427 = x_18137 & x_18138;
assign x_49428 = x_49426 & x_49427;
assign x_49429 = x_49425 & x_49428;
assign x_49430 = x_49422 & x_49429;
assign x_49431 = x_18139 & x_18140;
assign x_49432 = x_18141 & x_18142;
assign x_49433 = x_49431 & x_49432;
assign x_49434 = x_18143 & x_18144;
assign x_49435 = x_18145 & x_18146;
assign x_49436 = x_49434 & x_49435;
assign x_49437 = x_49433 & x_49436;
assign x_49438 = x_18147 & x_18148;
assign x_49439 = x_18149 & x_18150;
assign x_49440 = x_49438 & x_49439;
assign x_49441 = x_18151 & x_18152;
assign x_49442 = x_18153 & x_18154;
assign x_49443 = x_49441 & x_49442;
assign x_49444 = x_49440 & x_49443;
assign x_49445 = x_49437 & x_49444;
assign x_49446 = x_49430 & x_49445;
assign x_49447 = x_49416 & x_49446;
assign x_49448 = x_18156 & x_18157;
assign x_49449 = x_18155 & x_49448;
assign x_49450 = x_18158 & x_18159;
assign x_49451 = x_18160 & x_18161;
assign x_49452 = x_49450 & x_49451;
assign x_49453 = x_49449 & x_49452;
assign x_49454 = x_18162 & x_18163;
assign x_49455 = x_18164 & x_18165;
assign x_49456 = x_49454 & x_49455;
assign x_49457 = x_18166 & x_18167;
assign x_49458 = x_18168 & x_18169;
assign x_49459 = x_49457 & x_49458;
assign x_49460 = x_49456 & x_49459;
assign x_49461 = x_49453 & x_49460;
assign x_49462 = x_18171 & x_18172;
assign x_49463 = x_18170 & x_49462;
assign x_49464 = x_18173 & x_18174;
assign x_49465 = x_18175 & x_18176;
assign x_49466 = x_49464 & x_49465;
assign x_49467 = x_49463 & x_49466;
assign x_49468 = x_18177 & x_18178;
assign x_49469 = x_18179 & x_18180;
assign x_49470 = x_49468 & x_49469;
assign x_49471 = x_18181 & x_18182;
assign x_49472 = x_18183 & x_18184;
assign x_49473 = x_49471 & x_49472;
assign x_49474 = x_49470 & x_49473;
assign x_49475 = x_49467 & x_49474;
assign x_49476 = x_49461 & x_49475;
assign x_49477 = x_18186 & x_18187;
assign x_49478 = x_18185 & x_49477;
assign x_49479 = x_18188 & x_18189;
assign x_49480 = x_18190 & x_18191;
assign x_49481 = x_49479 & x_49480;
assign x_49482 = x_49478 & x_49481;
assign x_49483 = x_18192 & x_18193;
assign x_49484 = x_18194 & x_18195;
assign x_49485 = x_49483 & x_49484;
assign x_49486 = x_18196 & x_18197;
assign x_49487 = x_18198 & x_18199;
assign x_49488 = x_49486 & x_49487;
assign x_49489 = x_49485 & x_49488;
assign x_49490 = x_49482 & x_49489;
assign x_49491 = x_18200 & x_18201;
assign x_49492 = x_18202 & x_18203;
assign x_49493 = x_49491 & x_49492;
assign x_49494 = x_18204 & x_18205;
assign x_49495 = x_18206 & x_18207;
assign x_49496 = x_49494 & x_49495;
assign x_49497 = x_49493 & x_49496;
assign x_49498 = x_18208 & x_18209;
assign x_49499 = x_18210 & x_18211;
assign x_49500 = x_49498 & x_49499;
assign x_49501 = x_18212 & x_18213;
assign x_49502 = x_18214 & x_18215;
assign x_49503 = x_49501 & x_49502;
assign x_49504 = x_49500 & x_49503;
assign x_49505 = x_49497 & x_49504;
assign x_49506 = x_49490 & x_49505;
assign x_49507 = x_49476 & x_49506;
assign x_49508 = x_49447 & x_49507;
assign x_49509 = x_18217 & x_18218;
assign x_49510 = x_18216 & x_49509;
assign x_49511 = x_18219 & x_18220;
assign x_49512 = x_18221 & x_18222;
assign x_49513 = x_49511 & x_49512;
assign x_49514 = x_49510 & x_49513;
assign x_49515 = x_18223 & x_18224;
assign x_49516 = x_18225 & x_18226;
assign x_49517 = x_49515 & x_49516;
assign x_49518 = x_18227 & x_18228;
assign x_49519 = x_18229 & x_18230;
assign x_49520 = x_49518 & x_49519;
assign x_49521 = x_49517 & x_49520;
assign x_49522 = x_49514 & x_49521;
assign x_49523 = x_18232 & x_18233;
assign x_49524 = x_18231 & x_49523;
assign x_49525 = x_18234 & x_18235;
assign x_49526 = x_18236 & x_18237;
assign x_49527 = x_49525 & x_49526;
assign x_49528 = x_49524 & x_49527;
assign x_49529 = x_18238 & x_18239;
assign x_49530 = x_18240 & x_18241;
assign x_49531 = x_49529 & x_49530;
assign x_49532 = x_18242 & x_18243;
assign x_49533 = x_18244 & x_18245;
assign x_49534 = x_49532 & x_49533;
assign x_49535 = x_49531 & x_49534;
assign x_49536 = x_49528 & x_49535;
assign x_49537 = x_49522 & x_49536;
assign x_49538 = x_18247 & x_18248;
assign x_49539 = x_18246 & x_49538;
assign x_49540 = x_18249 & x_18250;
assign x_49541 = x_18251 & x_18252;
assign x_49542 = x_49540 & x_49541;
assign x_49543 = x_49539 & x_49542;
assign x_49544 = x_18253 & x_18254;
assign x_49545 = x_18255 & x_18256;
assign x_49546 = x_49544 & x_49545;
assign x_49547 = x_18257 & x_18258;
assign x_49548 = x_18259 & x_18260;
assign x_49549 = x_49547 & x_49548;
assign x_49550 = x_49546 & x_49549;
assign x_49551 = x_49543 & x_49550;
assign x_49552 = x_18261 & x_18262;
assign x_49553 = x_18263 & x_18264;
assign x_49554 = x_49552 & x_49553;
assign x_49555 = x_18265 & x_18266;
assign x_49556 = x_18267 & x_18268;
assign x_49557 = x_49555 & x_49556;
assign x_49558 = x_49554 & x_49557;
assign x_49559 = x_18269 & x_18270;
assign x_49560 = x_18271 & x_18272;
assign x_49561 = x_49559 & x_49560;
assign x_49562 = x_18273 & x_18274;
assign x_49563 = x_18275 & x_18276;
assign x_49564 = x_49562 & x_49563;
assign x_49565 = x_49561 & x_49564;
assign x_49566 = x_49558 & x_49565;
assign x_49567 = x_49551 & x_49566;
assign x_49568 = x_49537 & x_49567;
assign x_49569 = x_18278 & x_18279;
assign x_49570 = x_18277 & x_49569;
assign x_49571 = x_18280 & x_18281;
assign x_49572 = x_18282 & x_18283;
assign x_49573 = x_49571 & x_49572;
assign x_49574 = x_49570 & x_49573;
assign x_49575 = x_18284 & x_18285;
assign x_49576 = x_18286 & x_18287;
assign x_49577 = x_49575 & x_49576;
assign x_49578 = x_18288 & x_18289;
assign x_49579 = x_18290 & x_18291;
assign x_49580 = x_49578 & x_49579;
assign x_49581 = x_49577 & x_49580;
assign x_49582 = x_49574 & x_49581;
assign x_49583 = x_18293 & x_18294;
assign x_49584 = x_18292 & x_49583;
assign x_49585 = x_18295 & x_18296;
assign x_49586 = x_18297 & x_18298;
assign x_49587 = x_49585 & x_49586;
assign x_49588 = x_49584 & x_49587;
assign x_49589 = x_18299 & x_18300;
assign x_49590 = x_18301 & x_18302;
assign x_49591 = x_49589 & x_49590;
assign x_49592 = x_18303 & x_18304;
assign x_49593 = x_18305 & x_18306;
assign x_49594 = x_49592 & x_49593;
assign x_49595 = x_49591 & x_49594;
assign x_49596 = x_49588 & x_49595;
assign x_49597 = x_49582 & x_49596;
assign x_49598 = x_18308 & x_18309;
assign x_49599 = x_18307 & x_49598;
assign x_49600 = x_18310 & x_18311;
assign x_49601 = x_18312 & x_18313;
assign x_49602 = x_49600 & x_49601;
assign x_49603 = x_49599 & x_49602;
assign x_49604 = x_18314 & x_18315;
assign x_49605 = x_18316 & x_18317;
assign x_49606 = x_49604 & x_49605;
assign x_49607 = x_18318 & x_18319;
assign x_49608 = x_18320 & x_18321;
assign x_49609 = x_49607 & x_49608;
assign x_49610 = x_49606 & x_49609;
assign x_49611 = x_49603 & x_49610;
assign x_49612 = x_18322 & x_18323;
assign x_49613 = x_18324 & x_18325;
assign x_49614 = x_49612 & x_49613;
assign x_49615 = x_18326 & x_18327;
assign x_49616 = x_18328 & x_18329;
assign x_49617 = x_49615 & x_49616;
assign x_49618 = x_49614 & x_49617;
assign x_49619 = x_18330 & x_18331;
assign x_49620 = x_18332 & x_18333;
assign x_49621 = x_49619 & x_49620;
assign x_49622 = x_18334 & x_18335;
assign x_49623 = x_18336 & x_18337;
assign x_49624 = x_49622 & x_49623;
assign x_49625 = x_49621 & x_49624;
assign x_49626 = x_49618 & x_49625;
assign x_49627 = x_49611 & x_49626;
assign x_49628 = x_49597 & x_49627;
assign x_49629 = x_49568 & x_49628;
assign x_49630 = x_49508 & x_49629;
assign x_49631 = x_18339 & x_18340;
assign x_49632 = x_18338 & x_49631;
assign x_49633 = x_18341 & x_18342;
assign x_49634 = x_18343 & x_18344;
assign x_49635 = x_49633 & x_49634;
assign x_49636 = x_49632 & x_49635;
assign x_49637 = x_18345 & x_18346;
assign x_49638 = x_18347 & x_18348;
assign x_49639 = x_49637 & x_49638;
assign x_49640 = x_18349 & x_18350;
assign x_49641 = x_18351 & x_18352;
assign x_49642 = x_49640 & x_49641;
assign x_49643 = x_49639 & x_49642;
assign x_49644 = x_49636 & x_49643;
assign x_49645 = x_18354 & x_18355;
assign x_49646 = x_18353 & x_49645;
assign x_49647 = x_18356 & x_18357;
assign x_49648 = x_18358 & x_18359;
assign x_49649 = x_49647 & x_49648;
assign x_49650 = x_49646 & x_49649;
assign x_49651 = x_18360 & x_18361;
assign x_49652 = x_18362 & x_18363;
assign x_49653 = x_49651 & x_49652;
assign x_49654 = x_18364 & x_18365;
assign x_49655 = x_18366 & x_18367;
assign x_49656 = x_49654 & x_49655;
assign x_49657 = x_49653 & x_49656;
assign x_49658 = x_49650 & x_49657;
assign x_49659 = x_49644 & x_49658;
assign x_49660 = x_18369 & x_18370;
assign x_49661 = x_18368 & x_49660;
assign x_49662 = x_18371 & x_18372;
assign x_49663 = x_18373 & x_18374;
assign x_49664 = x_49662 & x_49663;
assign x_49665 = x_49661 & x_49664;
assign x_49666 = x_18375 & x_18376;
assign x_49667 = x_18377 & x_18378;
assign x_49668 = x_49666 & x_49667;
assign x_49669 = x_18379 & x_18380;
assign x_49670 = x_18381 & x_18382;
assign x_49671 = x_49669 & x_49670;
assign x_49672 = x_49668 & x_49671;
assign x_49673 = x_49665 & x_49672;
assign x_49674 = x_18383 & x_18384;
assign x_49675 = x_18385 & x_18386;
assign x_49676 = x_49674 & x_49675;
assign x_49677 = x_18387 & x_18388;
assign x_49678 = x_18389 & x_18390;
assign x_49679 = x_49677 & x_49678;
assign x_49680 = x_49676 & x_49679;
assign x_49681 = x_18391 & x_18392;
assign x_49682 = x_18393 & x_18394;
assign x_49683 = x_49681 & x_49682;
assign x_49684 = x_18395 & x_18396;
assign x_49685 = x_18397 & x_18398;
assign x_49686 = x_49684 & x_49685;
assign x_49687 = x_49683 & x_49686;
assign x_49688 = x_49680 & x_49687;
assign x_49689 = x_49673 & x_49688;
assign x_49690 = x_49659 & x_49689;
assign x_49691 = x_18400 & x_18401;
assign x_49692 = x_18399 & x_49691;
assign x_49693 = x_18402 & x_18403;
assign x_49694 = x_18404 & x_18405;
assign x_49695 = x_49693 & x_49694;
assign x_49696 = x_49692 & x_49695;
assign x_49697 = x_18406 & x_18407;
assign x_49698 = x_18408 & x_18409;
assign x_49699 = x_49697 & x_49698;
assign x_49700 = x_18410 & x_18411;
assign x_49701 = x_18412 & x_18413;
assign x_49702 = x_49700 & x_49701;
assign x_49703 = x_49699 & x_49702;
assign x_49704 = x_49696 & x_49703;
assign x_49705 = x_18415 & x_18416;
assign x_49706 = x_18414 & x_49705;
assign x_49707 = x_18417 & x_18418;
assign x_49708 = x_18419 & x_18420;
assign x_49709 = x_49707 & x_49708;
assign x_49710 = x_49706 & x_49709;
assign x_49711 = x_18421 & x_18422;
assign x_49712 = x_18423 & x_18424;
assign x_49713 = x_49711 & x_49712;
assign x_49714 = x_18425 & x_18426;
assign x_49715 = x_18427 & x_18428;
assign x_49716 = x_49714 & x_49715;
assign x_49717 = x_49713 & x_49716;
assign x_49718 = x_49710 & x_49717;
assign x_49719 = x_49704 & x_49718;
assign x_49720 = x_18430 & x_18431;
assign x_49721 = x_18429 & x_49720;
assign x_49722 = x_18432 & x_18433;
assign x_49723 = x_18434 & x_18435;
assign x_49724 = x_49722 & x_49723;
assign x_49725 = x_49721 & x_49724;
assign x_49726 = x_18436 & x_18437;
assign x_49727 = x_18438 & x_18439;
assign x_49728 = x_49726 & x_49727;
assign x_49729 = x_18440 & x_18441;
assign x_49730 = x_18442 & x_18443;
assign x_49731 = x_49729 & x_49730;
assign x_49732 = x_49728 & x_49731;
assign x_49733 = x_49725 & x_49732;
assign x_49734 = x_18444 & x_18445;
assign x_49735 = x_18446 & x_18447;
assign x_49736 = x_49734 & x_49735;
assign x_49737 = x_18448 & x_18449;
assign x_49738 = x_18450 & x_18451;
assign x_49739 = x_49737 & x_49738;
assign x_49740 = x_49736 & x_49739;
assign x_49741 = x_18452 & x_18453;
assign x_49742 = x_18454 & x_18455;
assign x_49743 = x_49741 & x_49742;
assign x_49744 = x_18456 & x_18457;
assign x_49745 = x_18458 & x_18459;
assign x_49746 = x_49744 & x_49745;
assign x_49747 = x_49743 & x_49746;
assign x_49748 = x_49740 & x_49747;
assign x_49749 = x_49733 & x_49748;
assign x_49750 = x_49719 & x_49749;
assign x_49751 = x_49690 & x_49750;
assign x_49752 = x_18461 & x_18462;
assign x_49753 = x_18460 & x_49752;
assign x_49754 = x_18463 & x_18464;
assign x_49755 = x_18465 & x_18466;
assign x_49756 = x_49754 & x_49755;
assign x_49757 = x_49753 & x_49756;
assign x_49758 = x_18467 & x_18468;
assign x_49759 = x_18469 & x_18470;
assign x_49760 = x_49758 & x_49759;
assign x_49761 = x_18471 & x_18472;
assign x_49762 = x_18473 & x_18474;
assign x_49763 = x_49761 & x_49762;
assign x_49764 = x_49760 & x_49763;
assign x_49765 = x_49757 & x_49764;
assign x_49766 = x_18476 & x_18477;
assign x_49767 = x_18475 & x_49766;
assign x_49768 = x_18478 & x_18479;
assign x_49769 = x_18480 & x_18481;
assign x_49770 = x_49768 & x_49769;
assign x_49771 = x_49767 & x_49770;
assign x_49772 = x_18482 & x_18483;
assign x_49773 = x_18484 & x_18485;
assign x_49774 = x_49772 & x_49773;
assign x_49775 = x_18486 & x_18487;
assign x_49776 = x_18488 & x_18489;
assign x_49777 = x_49775 & x_49776;
assign x_49778 = x_49774 & x_49777;
assign x_49779 = x_49771 & x_49778;
assign x_49780 = x_49765 & x_49779;
assign x_49781 = x_18491 & x_18492;
assign x_49782 = x_18490 & x_49781;
assign x_49783 = x_18493 & x_18494;
assign x_49784 = x_18495 & x_18496;
assign x_49785 = x_49783 & x_49784;
assign x_49786 = x_49782 & x_49785;
assign x_49787 = x_18497 & x_18498;
assign x_49788 = x_18499 & x_18500;
assign x_49789 = x_49787 & x_49788;
assign x_49790 = x_18501 & x_18502;
assign x_49791 = x_18503 & x_18504;
assign x_49792 = x_49790 & x_49791;
assign x_49793 = x_49789 & x_49792;
assign x_49794 = x_49786 & x_49793;
assign x_49795 = x_18505 & x_18506;
assign x_49796 = x_18507 & x_18508;
assign x_49797 = x_49795 & x_49796;
assign x_49798 = x_18509 & x_18510;
assign x_49799 = x_18511 & x_18512;
assign x_49800 = x_49798 & x_49799;
assign x_49801 = x_49797 & x_49800;
assign x_49802 = x_18513 & x_18514;
assign x_49803 = x_18515 & x_18516;
assign x_49804 = x_49802 & x_49803;
assign x_49805 = x_18517 & x_18518;
assign x_49806 = x_18519 & x_18520;
assign x_49807 = x_49805 & x_49806;
assign x_49808 = x_49804 & x_49807;
assign x_49809 = x_49801 & x_49808;
assign x_49810 = x_49794 & x_49809;
assign x_49811 = x_49780 & x_49810;
assign x_49812 = x_18522 & x_18523;
assign x_49813 = x_18521 & x_49812;
assign x_49814 = x_18524 & x_18525;
assign x_49815 = x_18526 & x_18527;
assign x_49816 = x_49814 & x_49815;
assign x_49817 = x_49813 & x_49816;
assign x_49818 = x_18528 & x_18529;
assign x_49819 = x_18530 & x_18531;
assign x_49820 = x_49818 & x_49819;
assign x_49821 = x_18532 & x_18533;
assign x_49822 = x_18534 & x_18535;
assign x_49823 = x_49821 & x_49822;
assign x_49824 = x_49820 & x_49823;
assign x_49825 = x_49817 & x_49824;
assign x_49826 = x_18536 & x_18537;
assign x_49827 = x_18538 & x_18539;
assign x_49828 = x_49826 & x_49827;
assign x_49829 = x_18540 & x_18541;
assign x_49830 = x_18542 & x_18543;
assign x_49831 = x_49829 & x_49830;
assign x_49832 = x_49828 & x_49831;
assign x_49833 = x_18544 & x_18545;
assign x_49834 = x_18546 & x_18547;
assign x_49835 = x_49833 & x_49834;
assign x_49836 = x_18548 & x_18549;
assign x_49837 = x_18550 & x_18551;
assign x_49838 = x_49836 & x_49837;
assign x_49839 = x_49835 & x_49838;
assign x_49840 = x_49832 & x_49839;
assign x_49841 = x_49825 & x_49840;
assign x_49842 = x_18553 & x_18554;
assign x_49843 = x_18552 & x_49842;
assign x_49844 = x_18555 & x_18556;
assign x_49845 = x_18557 & x_18558;
assign x_49846 = x_49844 & x_49845;
assign x_49847 = x_49843 & x_49846;
assign x_49848 = x_18559 & x_18560;
assign x_49849 = x_18561 & x_18562;
assign x_49850 = x_49848 & x_49849;
assign x_49851 = x_18563 & x_18564;
assign x_49852 = x_18565 & x_18566;
assign x_49853 = x_49851 & x_49852;
assign x_49854 = x_49850 & x_49853;
assign x_49855 = x_49847 & x_49854;
assign x_49856 = x_18567 & x_18568;
assign x_49857 = x_18569 & x_18570;
assign x_49858 = x_49856 & x_49857;
assign x_49859 = x_18571 & x_18572;
assign x_49860 = x_18573 & x_18574;
assign x_49861 = x_49859 & x_49860;
assign x_49862 = x_49858 & x_49861;
assign x_49863 = x_18575 & x_18576;
assign x_49864 = x_18577 & x_18578;
assign x_49865 = x_49863 & x_49864;
assign x_49866 = x_18579 & x_18580;
assign x_49867 = x_18581 & x_18582;
assign x_49868 = x_49866 & x_49867;
assign x_49869 = x_49865 & x_49868;
assign x_49870 = x_49862 & x_49869;
assign x_49871 = x_49855 & x_49870;
assign x_49872 = x_49841 & x_49871;
assign x_49873 = x_49811 & x_49872;
assign x_49874 = x_49751 & x_49873;
assign x_49875 = x_49630 & x_49874;
assign x_49876 = x_49387 & x_49875;
assign x_49877 = x_18584 & x_18585;
assign x_49878 = x_18583 & x_49877;
assign x_49879 = x_18586 & x_18587;
assign x_49880 = x_18588 & x_18589;
assign x_49881 = x_49879 & x_49880;
assign x_49882 = x_49878 & x_49881;
assign x_49883 = x_18590 & x_18591;
assign x_49884 = x_18592 & x_18593;
assign x_49885 = x_49883 & x_49884;
assign x_49886 = x_18594 & x_18595;
assign x_49887 = x_18596 & x_18597;
assign x_49888 = x_49886 & x_49887;
assign x_49889 = x_49885 & x_49888;
assign x_49890 = x_49882 & x_49889;
assign x_49891 = x_18599 & x_18600;
assign x_49892 = x_18598 & x_49891;
assign x_49893 = x_18601 & x_18602;
assign x_49894 = x_18603 & x_18604;
assign x_49895 = x_49893 & x_49894;
assign x_49896 = x_49892 & x_49895;
assign x_49897 = x_18605 & x_18606;
assign x_49898 = x_18607 & x_18608;
assign x_49899 = x_49897 & x_49898;
assign x_49900 = x_18609 & x_18610;
assign x_49901 = x_18611 & x_18612;
assign x_49902 = x_49900 & x_49901;
assign x_49903 = x_49899 & x_49902;
assign x_49904 = x_49896 & x_49903;
assign x_49905 = x_49890 & x_49904;
assign x_49906 = x_18614 & x_18615;
assign x_49907 = x_18613 & x_49906;
assign x_49908 = x_18616 & x_18617;
assign x_49909 = x_18618 & x_18619;
assign x_49910 = x_49908 & x_49909;
assign x_49911 = x_49907 & x_49910;
assign x_49912 = x_18620 & x_18621;
assign x_49913 = x_18622 & x_18623;
assign x_49914 = x_49912 & x_49913;
assign x_49915 = x_18624 & x_18625;
assign x_49916 = x_18626 & x_18627;
assign x_49917 = x_49915 & x_49916;
assign x_49918 = x_49914 & x_49917;
assign x_49919 = x_49911 & x_49918;
assign x_49920 = x_18628 & x_18629;
assign x_49921 = x_18630 & x_18631;
assign x_49922 = x_49920 & x_49921;
assign x_49923 = x_18632 & x_18633;
assign x_49924 = x_18634 & x_18635;
assign x_49925 = x_49923 & x_49924;
assign x_49926 = x_49922 & x_49925;
assign x_49927 = x_18636 & x_18637;
assign x_49928 = x_18638 & x_18639;
assign x_49929 = x_49927 & x_49928;
assign x_49930 = x_18640 & x_18641;
assign x_49931 = x_18642 & x_18643;
assign x_49932 = x_49930 & x_49931;
assign x_49933 = x_49929 & x_49932;
assign x_49934 = x_49926 & x_49933;
assign x_49935 = x_49919 & x_49934;
assign x_49936 = x_49905 & x_49935;
assign x_49937 = x_18645 & x_18646;
assign x_49938 = x_18644 & x_49937;
assign x_49939 = x_18647 & x_18648;
assign x_49940 = x_18649 & x_18650;
assign x_49941 = x_49939 & x_49940;
assign x_49942 = x_49938 & x_49941;
assign x_49943 = x_18651 & x_18652;
assign x_49944 = x_18653 & x_18654;
assign x_49945 = x_49943 & x_49944;
assign x_49946 = x_18655 & x_18656;
assign x_49947 = x_18657 & x_18658;
assign x_49948 = x_49946 & x_49947;
assign x_49949 = x_49945 & x_49948;
assign x_49950 = x_49942 & x_49949;
assign x_49951 = x_18660 & x_18661;
assign x_49952 = x_18659 & x_49951;
assign x_49953 = x_18662 & x_18663;
assign x_49954 = x_18664 & x_18665;
assign x_49955 = x_49953 & x_49954;
assign x_49956 = x_49952 & x_49955;
assign x_49957 = x_18666 & x_18667;
assign x_49958 = x_18668 & x_18669;
assign x_49959 = x_49957 & x_49958;
assign x_49960 = x_18670 & x_18671;
assign x_49961 = x_18672 & x_18673;
assign x_49962 = x_49960 & x_49961;
assign x_49963 = x_49959 & x_49962;
assign x_49964 = x_49956 & x_49963;
assign x_49965 = x_49950 & x_49964;
assign x_49966 = x_18675 & x_18676;
assign x_49967 = x_18674 & x_49966;
assign x_49968 = x_18677 & x_18678;
assign x_49969 = x_18679 & x_18680;
assign x_49970 = x_49968 & x_49969;
assign x_49971 = x_49967 & x_49970;
assign x_49972 = x_18681 & x_18682;
assign x_49973 = x_18683 & x_18684;
assign x_49974 = x_49972 & x_49973;
assign x_49975 = x_18685 & x_18686;
assign x_49976 = x_18687 & x_18688;
assign x_49977 = x_49975 & x_49976;
assign x_49978 = x_49974 & x_49977;
assign x_49979 = x_49971 & x_49978;
assign x_49980 = x_18689 & x_18690;
assign x_49981 = x_18691 & x_18692;
assign x_49982 = x_49980 & x_49981;
assign x_49983 = x_18693 & x_18694;
assign x_49984 = x_18695 & x_18696;
assign x_49985 = x_49983 & x_49984;
assign x_49986 = x_49982 & x_49985;
assign x_49987 = x_18697 & x_18698;
assign x_49988 = x_18699 & x_18700;
assign x_49989 = x_49987 & x_49988;
assign x_49990 = x_18701 & x_18702;
assign x_49991 = x_18703 & x_18704;
assign x_49992 = x_49990 & x_49991;
assign x_49993 = x_49989 & x_49992;
assign x_49994 = x_49986 & x_49993;
assign x_49995 = x_49979 & x_49994;
assign x_49996 = x_49965 & x_49995;
assign x_49997 = x_49936 & x_49996;
assign x_49998 = x_18706 & x_18707;
assign x_49999 = x_18705 & x_49998;
assign x_50000 = x_18708 & x_18709;
assign x_50001 = x_18710 & x_18711;
assign x_50002 = x_50000 & x_50001;
assign x_50003 = x_49999 & x_50002;
assign x_50004 = x_18712 & x_18713;
assign x_50005 = x_18714 & x_18715;
assign x_50006 = x_50004 & x_50005;
assign x_50007 = x_18716 & x_18717;
assign x_50008 = x_18718 & x_18719;
assign x_50009 = x_50007 & x_50008;
assign x_50010 = x_50006 & x_50009;
assign x_50011 = x_50003 & x_50010;
assign x_50012 = x_18721 & x_18722;
assign x_50013 = x_18720 & x_50012;
assign x_50014 = x_18723 & x_18724;
assign x_50015 = x_18725 & x_18726;
assign x_50016 = x_50014 & x_50015;
assign x_50017 = x_50013 & x_50016;
assign x_50018 = x_18727 & x_18728;
assign x_50019 = x_18729 & x_18730;
assign x_50020 = x_50018 & x_50019;
assign x_50021 = x_18731 & x_18732;
assign x_50022 = x_18733 & x_18734;
assign x_50023 = x_50021 & x_50022;
assign x_50024 = x_50020 & x_50023;
assign x_50025 = x_50017 & x_50024;
assign x_50026 = x_50011 & x_50025;
assign x_50027 = x_18736 & x_18737;
assign x_50028 = x_18735 & x_50027;
assign x_50029 = x_18738 & x_18739;
assign x_50030 = x_18740 & x_18741;
assign x_50031 = x_50029 & x_50030;
assign x_50032 = x_50028 & x_50031;
assign x_50033 = x_18742 & x_18743;
assign x_50034 = x_18744 & x_18745;
assign x_50035 = x_50033 & x_50034;
assign x_50036 = x_18746 & x_18747;
assign x_50037 = x_18748 & x_18749;
assign x_50038 = x_50036 & x_50037;
assign x_50039 = x_50035 & x_50038;
assign x_50040 = x_50032 & x_50039;
assign x_50041 = x_18750 & x_18751;
assign x_50042 = x_18752 & x_18753;
assign x_50043 = x_50041 & x_50042;
assign x_50044 = x_18754 & x_18755;
assign x_50045 = x_18756 & x_18757;
assign x_50046 = x_50044 & x_50045;
assign x_50047 = x_50043 & x_50046;
assign x_50048 = x_18758 & x_18759;
assign x_50049 = x_18760 & x_18761;
assign x_50050 = x_50048 & x_50049;
assign x_50051 = x_18762 & x_18763;
assign x_50052 = x_18764 & x_18765;
assign x_50053 = x_50051 & x_50052;
assign x_50054 = x_50050 & x_50053;
assign x_50055 = x_50047 & x_50054;
assign x_50056 = x_50040 & x_50055;
assign x_50057 = x_50026 & x_50056;
assign x_50058 = x_18767 & x_18768;
assign x_50059 = x_18766 & x_50058;
assign x_50060 = x_18769 & x_18770;
assign x_50061 = x_18771 & x_18772;
assign x_50062 = x_50060 & x_50061;
assign x_50063 = x_50059 & x_50062;
assign x_50064 = x_18773 & x_18774;
assign x_50065 = x_18775 & x_18776;
assign x_50066 = x_50064 & x_50065;
assign x_50067 = x_18777 & x_18778;
assign x_50068 = x_18779 & x_18780;
assign x_50069 = x_50067 & x_50068;
assign x_50070 = x_50066 & x_50069;
assign x_50071 = x_50063 & x_50070;
assign x_50072 = x_18782 & x_18783;
assign x_50073 = x_18781 & x_50072;
assign x_50074 = x_18784 & x_18785;
assign x_50075 = x_18786 & x_18787;
assign x_50076 = x_50074 & x_50075;
assign x_50077 = x_50073 & x_50076;
assign x_50078 = x_18788 & x_18789;
assign x_50079 = x_18790 & x_18791;
assign x_50080 = x_50078 & x_50079;
assign x_50081 = x_18792 & x_18793;
assign x_50082 = x_18794 & x_18795;
assign x_50083 = x_50081 & x_50082;
assign x_50084 = x_50080 & x_50083;
assign x_50085 = x_50077 & x_50084;
assign x_50086 = x_50071 & x_50085;
assign x_50087 = x_18797 & x_18798;
assign x_50088 = x_18796 & x_50087;
assign x_50089 = x_18799 & x_18800;
assign x_50090 = x_18801 & x_18802;
assign x_50091 = x_50089 & x_50090;
assign x_50092 = x_50088 & x_50091;
assign x_50093 = x_18803 & x_18804;
assign x_50094 = x_18805 & x_18806;
assign x_50095 = x_50093 & x_50094;
assign x_50096 = x_18807 & x_18808;
assign x_50097 = x_18809 & x_18810;
assign x_50098 = x_50096 & x_50097;
assign x_50099 = x_50095 & x_50098;
assign x_50100 = x_50092 & x_50099;
assign x_50101 = x_18811 & x_18812;
assign x_50102 = x_18813 & x_18814;
assign x_50103 = x_50101 & x_50102;
assign x_50104 = x_18815 & x_18816;
assign x_50105 = x_18817 & x_18818;
assign x_50106 = x_50104 & x_50105;
assign x_50107 = x_50103 & x_50106;
assign x_50108 = x_18819 & x_18820;
assign x_50109 = x_18821 & x_18822;
assign x_50110 = x_50108 & x_50109;
assign x_50111 = x_18823 & x_18824;
assign x_50112 = x_18825 & x_18826;
assign x_50113 = x_50111 & x_50112;
assign x_50114 = x_50110 & x_50113;
assign x_50115 = x_50107 & x_50114;
assign x_50116 = x_50100 & x_50115;
assign x_50117 = x_50086 & x_50116;
assign x_50118 = x_50057 & x_50117;
assign x_50119 = x_49997 & x_50118;
assign x_50120 = x_18828 & x_18829;
assign x_50121 = x_18827 & x_50120;
assign x_50122 = x_18830 & x_18831;
assign x_50123 = x_18832 & x_18833;
assign x_50124 = x_50122 & x_50123;
assign x_50125 = x_50121 & x_50124;
assign x_50126 = x_18834 & x_18835;
assign x_50127 = x_18836 & x_18837;
assign x_50128 = x_50126 & x_50127;
assign x_50129 = x_18838 & x_18839;
assign x_50130 = x_18840 & x_18841;
assign x_50131 = x_50129 & x_50130;
assign x_50132 = x_50128 & x_50131;
assign x_50133 = x_50125 & x_50132;
assign x_50134 = x_18843 & x_18844;
assign x_50135 = x_18842 & x_50134;
assign x_50136 = x_18845 & x_18846;
assign x_50137 = x_18847 & x_18848;
assign x_50138 = x_50136 & x_50137;
assign x_50139 = x_50135 & x_50138;
assign x_50140 = x_18849 & x_18850;
assign x_50141 = x_18851 & x_18852;
assign x_50142 = x_50140 & x_50141;
assign x_50143 = x_18853 & x_18854;
assign x_50144 = x_18855 & x_18856;
assign x_50145 = x_50143 & x_50144;
assign x_50146 = x_50142 & x_50145;
assign x_50147 = x_50139 & x_50146;
assign x_50148 = x_50133 & x_50147;
assign x_50149 = x_18858 & x_18859;
assign x_50150 = x_18857 & x_50149;
assign x_50151 = x_18860 & x_18861;
assign x_50152 = x_18862 & x_18863;
assign x_50153 = x_50151 & x_50152;
assign x_50154 = x_50150 & x_50153;
assign x_50155 = x_18864 & x_18865;
assign x_50156 = x_18866 & x_18867;
assign x_50157 = x_50155 & x_50156;
assign x_50158 = x_18868 & x_18869;
assign x_50159 = x_18870 & x_18871;
assign x_50160 = x_50158 & x_50159;
assign x_50161 = x_50157 & x_50160;
assign x_50162 = x_50154 & x_50161;
assign x_50163 = x_18872 & x_18873;
assign x_50164 = x_18874 & x_18875;
assign x_50165 = x_50163 & x_50164;
assign x_50166 = x_18876 & x_18877;
assign x_50167 = x_18878 & x_18879;
assign x_50168 = x_50166 & x_50167;
assign x_50169 = x_50165 & x_50168;
assign x_50170 = x_18880 & x_18881;
assign x_50171 = x_18882 & x_18883;
assign x_50172 = x_50170 & x_50171;
assign x_50173 = x_18884 & x_18885;
assign x_50174 = x_18886 & x_18887;
assign x_50175 = x_50173 & x_50174;
assign x_50176 = x_50172 & x_50175;
assign x_50177 = x_50169 & x_50176;
assign x_50178 = x_50162 & x_50177;
assign x_50179 = x_50148 & x_50178;
assign x_50180 = x_18889 & x_18890;
assign x_50181 = x_18888 & x_50180;
assign x_50182 = x_18891 & x_18892;
assign x_50183 = x_18893 & x_18894;
assign x_50184 = x_50182 & x_50183;
assign x_50185 = x_50181 & x_50184;
assign x_50186 = x_18895 & x_18896;
assign x_50187 = x_18897 & x_18898;
assign x_50188 = x_50186 & x_50187;
assign x_50189 = x_18899 & x_18900;
assign x_50190 = x_18901 & x_18902;
assign x_50191 = x_50189 & x_50190;
assign x_50192 = x_50188 & x_50191;
assign x_50193 = x_50185 & x_50192;
assign x_50194 = x_18904 & x_18905;
assign x_50195 = x_18903 & x_50194;
assign x_50196 = x_18906 & x_18907;
assign x_50197 = x_18908 & x_18909;
assign x_50198 = x_50196 & x_50197;
assign x_50199 = x_50195 & x_50198;
assign x_50200 = x_18910 & x_18911;
assign x_50201 = x_18912 & x_18913;
assign x_50202 = x_50200 & x_50201;
assign x_50203 = x_18914 & x_18915;
assign x_50204 = x_18916 & x_18917;
assign x_50205 = x_50203 & x_50204;
assign x_50206 = x_50202 & x_50205;
assign x_50207 = x_50199 & x_50206;
assign x_50208 = x_50193 & x_50207;
assign x_50209 = x_18919 & x_18920;
assign x_50210 = x_18918 & x_50209;
assign x_50211 = x_18921 & x_18922;
assign x_50212 = x_18923 & x_18924;
assign x_50213 = x_50211 & x_50212;
assign x_50214 = x_50210 & x_50213;
assign x_50215 = x_18925 & x_18926;
assign x_50216 = x_18927 & x_18928;
assign x_50217 = x_50215 & x_50216;
assign x_50218 = x_18929 & x_18930;
assign x_50219 = x_18931 & x_18932;
assign x_50220 = x_50218 & x_50219;
assign x_50221 = x_50217 & x_50220;
assign x_50222 = x_50214 & x_50221;
assign x_50223 = x_18933 & x_18934;
assign x_50224 = x_18935 & x_18936;
assign x_50225 = x_50223 & x_50224;
assign x_50226 = x_18937 & x_18938;
assign x_50227 = x_18939 & x_18940;
assign x_50228 = x_50226 & x_50227;
assign x_50229 = x_50225 & x_50228;
assign x_50230 = x_18941 & x_18942;
assign x_50231 = x_18943 & x_18944;
assign x_50232 = x_50230 & x_50231;
assign x_50233 = x_18945 & x_18946;
assign x_50234 = x_18947 & x_18948;
assign x_50235 = x_50233 & x_50234;
assign x_50236 = x_50232 & x_50235;
assign x_50237 = x_50229 & x_50236;
assign x_50238 = x_50222 & x_50237;
assign x_50239 = x_50208 & x_50238;
assign x_50240 = x_50179 & x_50239;
assign x_50241 = x_18950 & x_18951;
assign x_50242 = x_18949 & x_50241;
assign x_50243 = x_18952 & x_18953;
assign x_50244 = x_18954 & x_18955;
assign x_50245 = x_50243 & x_50244;
assign x_50246 = x_50242 & x_50245;
assign x_50247 = x_18956 & x_18957;
assign x_50248 = x_18958 & x_18959;
assign x_50249 = x_50247 & x_50248;
assign x_50250 = x_18960 & x_18961;
assign x_50251 = x_18962 & x_18963;
assign x_50252 = x_50250 & x_50251;
assign x_50253 = x_50249 & x_50252;
assign x_50254 = x_50246 & x_50253;
assign x_50255 = x_18965 & x_18966;
assign x_50256 = x_18964 & x_50255;
assign x_50257 = x_18967 & x_18968;
assign x_50258 = x_18969 & x_18970;
assign x_50259 = x_50257 & x_50258;
assign x_50260 = x_50256 & x_50259;
assign x_50261 = x_18971 & x_18972;
assign x_50262 = x_18973 & x_18974;
assign x_50263 = x_50261 & x_50262;
assign x_50264 = x_18975 & x_18976;
assign x_50265 = x_18977 & x_18978;
assign x_50266 = x_50264 & x_50265;
assign x_50267 = x_50263 & x_50266;
assign x_50268 = x_50260 & x_50267;
assign x_50269 = x_50254 & x_50268;
assign x_50270 = x_18980 & x_18981;
assign x_50271 = x_18979 & x_50270;
assign x_50272 = x_18982 & x_18983;
assign x_50273 = x_18984 & x_18985;
assign x_50274 = x_50272 & x_50273;
assign x_50275 = x_50271 & x_50274;
assign x_50276 = x_18986 & x_18987;
assign x_50277 = x_18988 & x_18989;
assign x_50278 = x_50276 & x_50277;
assign x_50279 = x_18990 & x_18991;
assign x_50280 = x_18992 & x_18993;
assign x_50281 = x_50279 & x_50280;
assign x_50282 = x_50278 & x_50281;
assign x_50283 = x_50275 & x_50282;
assign x_50284 = x_18994 & x_18995;
assign x_50285 = x_18996 & x_18997;
assign x_50286 = x_50284 & x_50285;
assign x_50287 = x_18998 & x_18999;
assign x_50288 = x_19000 & x_19001;
assign x_50289 = x_50287 & x_50288;
assign x_50290 = x_50286 & x_50289;
assign x_50291 = x_19002 & x_19003;
assign x_50292 = x_19004 & x_19005;
assign x_50293 = x_50291 & x_50292;
assign x_50294 = x_19006 & x_19007;
assign x_50295 = x_19008 & x_19009;
assign x_50296 = x_50294 & x_50295;
assign x_50297 = x_50293 & x_50296;
assign x_50298 = x_50290 & x_50297;
assign x_50299 = x_50283 & x_50298;
assign x_50300 = x_50269 & x_50299;
assign x_50301 = x_19011 & x_19012;
assign x_50302 = x_19010 & x_50301;
assign x_50303 = x_19013 & x_19014;
assign x_50304 = x_19015 & x_19016;
assign x_50305 = x_50303 & x_50304;
assign x_50306 = x_50302 & x_50305;
assign x_50307 = x_19017 & x_19018;
assign x_50308 = x_19019 & x_19020;
assign x_50309 = x_50307 & x_50308;
assign x_50310 = x_19021 & x_19022;
assign x_50311 = x_19023 & x_19024;
assign x_50312 = x_50310 & x_50311;
assign x_50313 = x_50309 & x_50312;
assign x_50314 = x_50306 & x_50313;
assign x_50315 = x_19025 & x_19026;
assign x_50316 = x_19027 & x_19028;
assign x_50317 = x_50315 & x_50316;
assign x_50318 = x_19029 & x_19030;
assign x_50319 = x_19031 & x_19032;
assign x_50320 = x_50318 & x_50319;
assign x_50321 = x_50317 & x_50320;
assign x_50322 = x_19033 & x_19034;
assign x_50323 = x_19035 & x_19036;
assign x_50324 = x_50322 & x_50323;
assign x_50325 = x_19037 & x_19038;
assign x_50326 = x_19039 & x_19040;
assign x_50327 = x_50325 & x_50326;
assign x_50328 = x_50324 & x_50327;
assign x_50329 = x_50321 & x_50328;
assign x_50330 = x_50314 & x_50329;
assign x_50331 = x_19042 & x_19043;
assign x_50332 = x_19041 & x_50331;
assign x_50333 = x_19044 & x_19045;
assign x_50334 = x_19046 & x_19047;
assign x_50335 = x_50333 & x_50334;
assign x_50336 = x_50332 & x_50335;
assign x_50337 = x_19048 & x_19049;
assign x_50338 = x_19050 & x_19051;
assign x_50339 = x_50337 & x_50338;
assign x_50340 = x_19052 & x_19053;
assign x_50341 = x_19054 & x_19055;
assign x_50342 = x_50340 & x_50341;
assign x_50343 = x_50339 & x_50342;
assign x_50344 = x_50336 & x_50343;
assign x_50345 = x_19056 & x_19057;
assign x_50346 = x_19058 & x_19059;
assign x_50347 = x_50345 & x_50346;
assign x_50348 = x_19060 & x_19061;
assign x_50349 = x_19062 & x_19063;
assign x_50350 = x_50348 & x_50349;
assign x_50351 = x_50347 & x_50350;
assign x_50352 = x_19064 & x_19065;
assign x_50353 = x_19066 & x_19067;
assign x_50354 = x_50352 & x_50353;
assign x_50355 = x_19068 & x_19069;
assign x_50356 = x_19070 & x_19071;
assign x_50357 = x_50355 & x_50356;
assign x_50358 = x_50354 & x_50357;
assign x_50359 = x_50351 & x_50358;
assign x_50360 = x_50344 & x_50359;
assign x_50361 = x_50330 & x_50360;
assign x_50362 = x_50300 & x_50361;
assign x_50363 = x_50240 & x_50362;
assign x_50364 = x_50119 & x_50363;
assign x_50365 = x_19073 & x_19074;
assign x_50366 = x_19072 & x_50365;
assign x_50367 = x_19075 & x_19076;
assign x_50368 = x_19077 & x_19078;
assign x_50369 = x_50367 & x_50368;
assign x_50370 = x_50366 & x_50369;
assign x_50371 = x_19079 & x_19080;
assign x_50372 = x_19081 & x_19082;
assign x_50373 = x_50371 & x_50372;
assign x_50374 = x_19083 & x_19084;
assign x_50375 = x_19085 & x_19086;
assign x_50376 = x_50374 & x_50375;
assign x_50377 = x_50373 & x_50376;
assign x_50378 = x_50370 & x_50377;
assign x_50379 = x_19088 & x_19089;
assign x_50380 = x_19087 & x_50379;
assign x_50381 = x_19090 & x_19091;
assign x_50382 = x_19092 & x_19093;
assign x_50383 = x_50381 & x_50382;
assign x_50384 = x_50380 & x_50383;
assign x_50385 = x_19094 & x_19095;
assign x_50386 = x_19096 & x_19097;
assign x_50387 = x_50385 & x_50386;
assign x_50388 = x_19098 & x_19099;
assign x_50389 = x_19100 & x_19101;
assign x_50390 = x_50388 & x_50389;
assign x_50391 = x_50387 & x_50390;
assign x_50392 = x_50384 & x_50391;
assign x_50393 = x_50378 & x_50392;
assign x_50394 = x_19103 & x_19104;
assign x_50395 = x_19102 & x_50394;
assign x_50396 = x_19105 & x_19106;
assign x_50397 = x_19107 & x_19108;
assign x_50398 = x_50396 & x_50397;
assign x_50399 = x_50395 & x_50398;
assign x_50400 = x_19109 & x_19110;
assign x_50401 = x_19111 & x_19112;
assign x_50402 = x_50400 & x_50401;
assign x_50403 = x_19113 & x_19114;
assign x_50404 = x_19115 & x_19116;
assign x_50405 = x_50403 & x_50404;
assign x_50406 = x_50402 & x_50405;
assign x_50407 = x_50399 & x_50406;
assign x_50408 = x_19117 & x_19118;
assign x_50409 = x_19119 & x_19120;
assign x_50410 = x_50408 & x_50409;
assign x_50411 = x_19121 & x_19122;
assign x_50412 = x_19123 & x_19124;
assign x_50413 = x_50411 & x_50412;
assign x_50414 = x_50410 & x_50413;
assign x_50415 = x_19125 & x_19126;
assign x_50416 = x_19127 & x_19128;
assign x_50417 = x_50415 & x_50416;
assign x_50418 = x_19129 & x_19130;
assign x_50419 = x_19131 & x_19132;
assign x_50420 = x_50418 & x_50419;
assign x_50421 = x_50417 & x_50420;
assign x_50422 = x_50414 & x_50421;
assign x_50423 = x_50407 & x_50422;
assign x_50424 = x_50393 & x_50423;
assign x_50425 = x_19134 & x_19135;
assign x_50426 = x_19133 & x_50425;
assign x_50427 = x_19136 & x_19137;
assign x_50428 = x_19138 & x_19139;
assign x_50429 = x_50427 & x_50428;
assign x_50430 = x_50426 & x_50429;
assign x_50431 = x_19140 & x_19141;
assign x_50432 = x_19142 & x_19143;
assign x_50433 = x_50431 & x_50432;
assign x_50434 = x_19144 & x_19145;
assign x_50435 = x_19146 & x_19147;
assign x_50436 = x_50434 & x_50435;
assign x_50437 = x_50433 & x_50436;
assign x_50438 = x_50430 & x_50437;
assign x_50439 = x_19149 & x_19150;
assign x_50440 = x_19148 & x_50439;
assign x_50441 = x_19151 & x_19152;
assign x_50442 = x_19153 & x_19154;
assign x_50443 = x_50441 & x_50442;
assign x_50444 = x_50440 & x_50443;
assign x_50445 = x_19155 & x_19156;
assign x_50446 = x_19157 & x_19158;
assign x_50447 = x_50445 & x_50446;
assign x_50448 = x_19159 & x_19160;
assign x_50449 = x_19161 & x_19162;
assign x_50450 = x_50448 & x_50449;
assign x_50451 = x_50447 & x_50450;
assign x_50452 = x_50444 & x_50451;
assign x_50453 = x_50438 & x_50452;
assign x_50454 = x_19164 & x_19165;
assign x_50455 = x_19163 & x_50454;
assign x_50456 = x_19166 & x_19167;
assign x_50457 = x_19168 & x_19169;
assign x_50458 = x_50456 & x_50457;
assign x_50459 = x_50455 & x_50458;
assign x_50460 = x_19170 & x_19171;
assign x_50461 = x_19172 & x_19173;
assign x_50462 = x_50460 & x_50461;
assign x_50463 = x_19174 & x_19175;
assign x_50464 = x_19176 & x_19177;
assign x_50465 = x_50463 & x_50464;
assign x_50466 = x_50462 & x_50465;
assign x_50467 = x_50459 & x_50466;
assign x_50468 = x_19178 & x_19179;
assign x_50469 = x_19180 & x_19181;
assign x_50470 = x_50468 & x_50469;
assign x_50471 = x_19182 & x_19183;
assign x_50472 = x_19184 & x_19185;
assign x_50473 = x_50471 & x_50472;
assign x_50474 = x_50470 & x_50473;
assign x_50475 = x_19186 & x_19187;
assign x_50476 = x_19188 & x_19189;
assign x_50477 = x_50475 & x_50476;
assign x_50478 = x_19190 & x_19191;
assign x_50479 = x_19192 & x_19193;
assign x_50480 = x_50478 & x_50479;
assign x_50481 = x_50477 & x_50480;
assign x_50482 = x_50474 & x_50481;
assign x_50483 = x_50467 & x_50482;
assign x_50484 = x_50453 & x_50483;
assign x_50485 = x_50424 & x_50484;
assign x_50486 = x_19195 & x_19196;
assign x_50487 = x_19194 & x_50486;
assign x_50488 = x_19197 & x_19198;
assign x_50489 = x_19199 & x_19200;
assign x_50490 = x_50488 & x_50489;
assign x_50491 = x_50487 & x_50490;
assign x_50492 = x_19201 & x_19202;
assign x_50493 = x_19203 & x_19204;
assign x_50494 = x_50492 & x_50493;
assign x_50495 = x_19205 & x_19206;
assign x_50496 = x_19207 & x_19208;
assign x_50497 = x_50495 & x_50496;
assign x_50498 = x_50494 & x_50497;
assign x_50499 = x_50491 & x_50498;
assign x_50500 = x_19210 & x_19211;
assign x_50501 = x_19209 & x_50500;
assign x_50502 = x_19212 & x_19213;
assign x_50503 = x_19214 & x_19215;
assign x_50504 = x_50502 & x_50503;
assign x_50505 = x_50501 & x_50504;
assign x_50506 = x_19216 & x_19217;
assign x_50507 = x_19218 & x_19219;
assign x_50508 = x_50506 & x_50507;
assign x_50509 = x_19220 & x_19221;
assign x_50510 = x_19222 & x_19223;
assign x_50511 = x_50509 & x_50510;
assign x_50512 = x_50508 & x_50511;
assign x_50513 = x_50505 & x_50512;
assign x_50514 = x_50499 & x_50513;
assign x_50515 = x_19225 & x_19226;
assign x_50516 = x_19224 & x_50515;
assign x_50517 = x_19227 & x_19228;
assign x_50518 = x_19229 & x_19230;
assign x_50519 = x_50517 & x_50518;
assign x_50520 = x_50516 & x_50519;
assign x_50521 = x_19231 & x_19232;
assign x_50522 = x_19233 & x_19234;
assign x_50523 = x_50521 & x_50522;
assign x_50524 = x_19235 & x_19236;
assign x_50525 = x_19237 & x_19238;
assign x_50526 = x_50524 & x_50525;
assign x_50527 = x_50523 & x_50526;
assign x_50528 = x_50520 & x_50527;
assign x_50529 = x_19239 & x_19240;
assign x_50530 = x_19241 & x_19242;
assign x_50531 = x_50529 & x_50530;
assign x_50532 = x_19243 & x_19244;
assign x_50533 = x_19245 & x_19246;
assign x_50534 = x_50532 & x_50533;
assign x_50535 = x_50531 & x_50534;
assign x_50536 = x_19247 & x_19248;
assign x_50537 = x_19249 & x_19250;
assign x_50538 = x_50536 & x_50537;
assign x_50539 = x_19251 & x_19252;
assign x_50540 = x_19253 & x_19254;
assign x_50541 = x_50539 & x_50540;
assign x_50542 = x_50538 & x_50541;
assign x_50543 = x_50535 & x_50542;
assign x_50544 = x_50528 & x_50543;
assign x_50545 = x_50514 & x_50544;
assign x_50546 = x_19256 & x_19257;
assign x_50547 = x_19255 & x_50546;
assign x_50548 = x_19258 & x_19259;
assign x_50549 = x_19260 & x_19261;
assign x_50550 = x_50548 & x_50549;
assign x_50551 = x_50547 & x_50550;
assign x_50552 = x_19262 & x_19263;
assign x_50553 = x_19264 & x_19265;
assign x_50554 = x_50552 & x_50553;
assign x_50555 = x_19266 & x_19267;
assign x_50556 = x_19268 & x_19269;
assign x_50557 = x_50555 & x_50556;
assign x_50558 = x_50554 & x_50557;
assign x_50559 = x_50551 & x_50558;
assign x_50560 = x_19271 & x_19272;
assign x_50561 = x_19270 & x_50560;
assign x_50562 = x_19273 & x_19274;
assign x_50563 = x_19275 & x_19276;
assign x_50564 = x_50562 & x_50563;
assign x_50565 = x_50561 & x_50564;
assign x_50566 = x_19277 & x_19278;
assign x_50567 = x_19279 & x_19280;
assign x_50568 = x_50566 & x_50567;
assign x_50569 = x_19281 & x_19282;
assign x_50570 = x_19283 & x_19284;
assign x_50571 = x_50569 & x_50570;
assign x_50572 = x_50568 & x_50571;
assign x_50573 = x_50565 & x_50572;
assign x_50574 = x_50559 & x_50573;
assign x_50575 = x_19286 & x_19287;
assign x_50576 = x_19285 & x_50575;
assign x_50577 = x_19288 & x_19289;
assign x_50578 = x_19290 & x_19291;
assign x_50579 = x_50577 & x_50578;
assign x_50580 = x_50576 & x_50579;
assign x_50581 = x_19292 & x_19293;
assign x_50582 = x_19294 & x_19295;
assign x_50583 = x_50581 & x_50582;
assign x_50584 = x_19296 & x_19297;
assign x_50585 = x_19298 & x_19299;
assign x_50586 = x_50584 & x_50585;
assign x_50587 = x_50583 & x_50586;
assign x_50588 = x_50580 & x_50587;
assign x_50589 = x_19300 & x_19301;
assign x_50590 = x_19302 & x_19303;
assign x_50591 = x_50589 & x_50590;
assign x_50592 = x_19304 & x_19305;
assign x_50593 = x_19306 & x_19307;
assign x_50594 = x_50592 & x_50593;
assign x_50595 = x_50591 & x_50594;
assign x_50596 = x_19308 & x_19309;
assign x_50597 = x_19310 & x_19311;
assign x_50598 = x_50596 & x_50597;
assign x_50599 = x_19312 & x_19313;
assign x_50600 = x_19314 & x_19315;
assign x_50601 = x_50599 & x_50600;
assign x_50602 = x_50598 & x_50601;
assign x_50603 = x_50595 & x_50602;
assign x_50604 = x_50588 & x_50603;
assign x_50605 = x_50574 & x_50604;
assign x_50606 = x_50545 & x_50605;
assign x_50607 = x_50485 & x_50606;
assign x_50608 = x_19317 & x_19318;
assign x_50609 = x_19316 & x_50608;
assign x_50610 = x_19319 & x_19320;
assign x_50611 = x_19321 & x_19322;
assign x_50612 = x_50610 & x_50611;
assign x_50613 = x_50609 & x_50612;
assign x_50614 = x_19323 & x_19324;
assign x_50615 = x_19325 & x_19326;
assign x_50616 = x_50614 & x_50615;
assign x_50617 = x_19327 & x_19328;
assign x_50618 = x_19329 & x_19330;
assign x_50619 = x_50617 & x_50618;
assign x_50620 = x_50616 & x_50619;
assign x_50621 = x_50613 & x_50620;
assign x_50622 = x_19332 & x_19333;
assign x_50623 = x_19331 & x_50622;
assign x_50624 = x_19334 & x_19335;
assign x_50625 = x_19336 & x_19337;
assign x_50626 = x_50624 & x_50625;
assign x_50627 = x_50623 & x_50626;
assign x_50628 = x_19338 & x_19339;
assign x_50629 = x_19340 & x_19341;
assign x_50630 = x_50628 & x_50629;
assign x_50631 = x_19342 & x_19343;
assign x_50632 = x_19344 & x_19345;
assign x_50633 = x_50631 & x_50632;
assign x_50634 = x_50630 & x_50633;
assign x_50635 = x_50627 & x_50634;
assign x_50636 = x_50621 & x_50635;
assign x_50637 = x_19347 & x_19348;
assign x_50638 = x_19346 & x_50637;
assign x_50639 = x_19349 & x_19350;
assign x_50640 = x_19351 & x_19352;
assign x_50641 = x_50639 & x_50640;
assign x_50642 = x_50638 & x_50641;
assign x_50643 = x_19353 & x_19354;
assign x_50644 = x_19355 & x_19356;
assign x_50645 = x_50643 & x_50644;
assign x_50646 = x_19357 & x_19358;
assign x_50647 = x_19359 & x_19360;
assign x_50648 = x_50646 & x_50647;
assign x_50649 = x_50645 & x_50648;
assign x_50650 = x_50642 & x_50649;
assign x_50651 = x_19361 & x_19362;
assign x_50652 = x_19363 & x_19364;
assign x_50653 = x_50651 & x_50652;
assign x_50654 = x_19365 & x_19366;
assign x_50655 = x_19367 & x_19368;
assign x_50656 = x_50654 & x_50655;
assign x_50657 = x_50653 & x_50656;
assign x_50658 = x_19369 & x_19370;
assign x_50659 = x_19371 & x_19372;
assign x_50660 = x_50658 & x_50659;
assign x_50661 = x_19373 & x_19374;
assign x_50662 = x_19375 & x_19376;
assign x_50663 = x_50661 & x_50662;
assign x_50664 = x_50660 & x_50663;
assign x_50665 = x_50657 & x_50664;
assign x_50666 = x_50650 & x_50665;
assign x_50667 = x_50636 & x_50666;
assign x_50668 = x_19378 & x_19379;
assign x_50669 = x_19377 & x_50668;
assign x_50670 = x_19380 & x_19381;
assign x_50671 = x_19382 & x_19383;
assign x_50672 = x_50670 & x_50671;
assign x_50673 = x_50669 & x_50672;
assign x_50674 = x_19384 & x_19385;
assign x_50675 = x_19386 & x_19387;
assign x_50676 = x_50674 & x_50675;
assign x_50677 = x_19388 & x_19389;
assign x_50678 = x_19390 & x_19391;
assign x_50679 = x_50677 & x_50678;
assign x_50680 = x_50676 & x_50679;
assign x_50681 = x_50673 & x_50680;
assign x_50682 = x_19393 & x_19394;
assign x_50683 = x_19392 & x_50682;
assign x_50684 = x_19395 & x_19396;
assign x_50685 = x_19397 & x_19398;
assign x_50686 = x_50684 & x_50685;
assign x_50687 = x_50683 & x_50686;
assign x_50688 = x_19399 & x_19400;
assign x_50689 = x_19401 & x_19402;
assign x_50690 = x_50688 & x_50689;
assign x_50691 = x_19403 & x_19404;
assign x_50692 = x_19405 & x_19406;
assign x_50693 = x_50691 & x_50692;
assign x_50694 = x_50690 & x_50693;
assign x_50695 = x_50687 & x_50694;
assign x_50696 = x_50681 & x_50695;
assign x_50697 = x_19408 & x_19409;
assign x_50698 = x_19407 & x_50697;
assign x_50699 = x_19410 & x_19411;
assign x_50700 = x_19412 & x_19413;
assign x_50701 = x_50699 & x_50700;
assign x_50702 = x_50698 & x_50701;
assign x_50703 = x_19414 & x_19415;
assign x_50704 = x_19416 & x_19417;
assign x_50705 = x_50703 & x_50704;
assign x_50706 = x_19418 & x_19419;
assign x_50707 = x_19420 & x_19421;
assign x_50708 = x_50706 & x_50707;
assign x_50709 = x_50705 & x_50708;
assign x_50710 = x_50702 & x_50709;
assign x_50711 = x_19422 & x_19423;
assign x_50712 = x_19424 & x_19425;
assign x_50713 = x_50711 & x_50712;
assign x_50714 = x_19426 & x_19427;
assign x_50715 = x_19428 & x_19429;
assign x_50716 = x_50714 & x_50715;
assign x_50717 = x_50713 & x_50716;
assign x_50718 = x_19430 & x_19431;
assign x_50719 = x_19432 & x_19433;
assign x_50720 = x_50718 & x_50719;
assign x_50721 = x_19434 & x_19435;
assign x_50722 = x_19436 & x_19437;
assign x_50723 = x_50721 & x_50722;
assign x_50724 = x_50720 & x_50723;
assign x_50725 = x_50717 & x_50724;
assign x_50726 = x_50710 & x_50725;
assign x_50727 = x_50696 & x_50726;
assign x_50728 = x_50667 & x_50727;
assign x_50729 = x_19439 & x_19440;
assign x_50730 = x_19438 & x_50729;
assign x_50731 = x_19441 & x_19442;
assign x_50732 = x_19443 & x_19444;
assign x_50733 = x_50731 & x_50732;
assign x_50734 = x_50730 & x_50733;
assign x_50735 = x_19445 & x_19446;
assign x_50736 = x_19447 & x_19448;
assign x_50737 = x_50735 & x_50736;
assign x_50738 = x_19449 & x_19450;
assign x_50739 = x_19451 & x_19452;
assign x_50740 = x_50738 & x_50739;
assign x_50741 = x_50737 & x_50740;
assign x_50742 = x_50734 & x_50741;
assign x_50743 = x_19454 & x_19455;
assign x_50744 = x_19453 & x_50743;
assign x_50745 = x_19456 & x_19457;
assign x_50746 = x_19458 & x_19459;
assign x_50747 = x_50745 & x_50746;
assign x_50748 = x_50744 & x_50747;
assign x_50749 = x_19460 & x_19461;
assign x_50750 = x_19462 & x_19463;
assign x_50751 = x_50749 & x_50750;
assign x_50752 = x_19464 & x_19465;
assign x_50753 = x_19466 & x_19467;
assign x_50754 = x_50752 & x_50753;
assign x_50755 = x_50751 & x_50754;
assign x_50756 = x_50748 & x_50755;
assign x_50757 = x_50742 & x_50756;
assign x_50758 = x_19469 & x_19470;
assign x_50759 = x_19468 & x_50758;
assign x_50760 = x_19471 & x_19472;
assign x_50761 = x_19473 & x_19474;
assign x_50762 = x_50760 & x_50761;
assign x_50763 = x_50759 & x_50762;
assign x_50764 = x_19475 & x_19476;
assign x_50765 = x_19477 & x_19478;
assign x_50766 = x_50764 & x_50765;
assign x_50767 = x_19479 & x_19480;
assign x_50768 = x_19481 & x_19482;
assign x_50769 = x_50767 & x_50768;
assign x_50770 = x_50766 & x_50769;
assign x_50771 = x_50763 & x_50770;
assign x_50772 = x_19483 & x_19484;
assign x_50773 = x_19485 & x_19486;
assign x_50774 = x_50772 & x_50773;
assign x_50775 = x_19487 & x_19488;
assign x_50776 = x_19489 & x_19490;
assign x_50777 = x_50775 & x_50776;
assign x_50778 = x_50774 & x_50777;
assign x_50779 = x_19491 & x_19492;
assign x_50780 = x_19493 & x_19494;
assign x_50781 = x_50779 & x_50780;
assign x_50782 = x_19495 & x_19496;
assign x_50783 = x_19497 & x_19498;
assign x_50784 = x_50782 & x_50783;
assign x_50785 = x_50781 & x_50784;
assign x_50786 = x_50778 & x_50785;
assign x_50787 = x_50771 & x_50786;
assign x_50788 = x_50757 & x_50787;
assign x_50789 = x_19500 & x_19501;
assign x_50790 = x_19499 & x_50789;
assign x_50791 = x_19502 & x_19503;
assign x_50792 = x_19504 & x_19505;
assign x_50793 = x_50791 & x_50792;
assign x_50794 = x_50790 & x_50793;
assign x_50795 = x_19506 & x_19507;
assign x_50796 = x_19508 & x_19509;
assign x_50797 = x_50795 & x_50796;
assign x_50798 = x_19510 & x_19511;
assign x_50799 = x_19512 & x_19513;
assign x_50800 = x_50798 & x_50799;
assign x_50801 = x_50797 & x_50800;
assign x_50802 = x_50794 & x_50801;
assign x_50803 = x_19514 & x_19515;
assign x_50804 = x_19516 & x_19517;
assign x_50805 = x_50803 & x_50804;
assign x_50806 = x_19518 & x_19519;
assign x_50807 = x_19520 & x_19521;
assign x_50808 = x_50806 & x_50807;
assign x_50809 = x_50805 & x_50808;
assign x_50810 = x_19522 & x_19523;
assign x_50811 = x_19524 & x_19525;
assign x_50812 = x_50810 & x_50811;
assign x_50813 = x_19526 & x_19527;
assign x_50814 = x_19528 & x_19529;
assign x_50815 = x_50813 & x_50814;
assign x_50816 = x_50812 & x_50815;
assign x_50817 = x_50809 & x_50816;
assign x_50818 = x_50802 & x_50817;
assign x_50819 = x_19531 & x_19532;
assign x_50820 = x_19530 & x_50819;
assign x_50821 = x_19533 & x_19534;
assign x_50822 = x_19535 & x_19536;
assign x_50823 = x_50821 & x_50822;
assign x_50824 = x_50820 & x_50823;
assign x_50825 = x_19537 & x_19538;
assign x_50826 = x_19539 & x_19540;
assign x_50827 = x_50825 & x_50826;
assign x_50828 = x_19541 & x_19542;
assign x_50829 = x_19543 & x_19544;
assign x_50830 = x_50828 & x_50829;
assign x_50831 = x_50827 & x_50830;
assign x_50832 = x_50824 & x_50831;
assign x_50833 = x_19545 & x_19546;
assign x_50834 = x_19547 & x_19548;
assign x_50835 = x_50833 & x_50834;
assign x_50836 = x_19549 & x_19550;
assign x_50837 = x_19551 & x_19552;
assign x_50838 = x_50836 & x_50837;
assign x_50839 = x_50835 & x_50838;
assign x_50840 = x_19553 & x_19554;
assign x_50841 = x_19555 & x_19556;
assign x_50842 = x_50840 & x_50841;
assign x_50843 = x_19557 & x_19558;
assign x_50844 = x_19559 & x_19560;
assign x_50845 = x_50843 & x_50844;
assign x_50846 = x_50842 & x_50845;
assign x_50847 = x_50839 & x_50846;
assign x_50848 = x_50832 & x_50847;
assign x_50849 = x_50818 & x_50848;
assign x_50850 = x_50788 & x_50849;
assign x_50851 = x_50728 & x_50850;
assign x_50852 = x_50607 & x_50851;
assign x_50853 = x_50364 & x_50852;
assign x_50854 = x_49876 & x_50853;
assign x_50855 = x_48899 & x_50854;
assign x_50856 = x_19562 & x_19563;
assign x_50857 = x_19561 & x_50856;
assign x_50858 = x_19564 & x_19565;
assign x_50859 = x_19566 & x_19567;
assign x_50860 = x_50858 & x_50859;
assign x_50861 = x_50857 & x_50860;
assign x_50862 = x_19568 & x_19569;
assign x_50863 = x_19570 & x_19571;
assign x_50864 = x_50862 & x_50863;
assign x_50865 = x_19572 & x_19573;
assign x_50866 = x_19574 & x_19575;
assign x_50867 = x_50865 & x_50866;
assign x_50868 = x_50864 & x_50867;
assign x_50869 = x_50861 & x_50868;
assign x_50870 = x_19577 & x_19578;
assign x_50871 = x_19576 & x_50870;
assign x_50872 = x_19579 & x_19580;
assign x_50873 = x_19581 & x_19582;
assign x_50874 = x_50872 & x_50873;
assign x_50875 = x_50871 & x_50874;
assign x_50876 = x_19583 & x_19584;
assign x_50877 = x_19585 & x_19586;
assign x_50878 = x_50876 & x_50877;
assign x_50879 = x_19587 & x_19588;
assign x_50880 = x_19589 & x_19590;
assign x_50881 = x_50879 & x_50880;
assign x_50882 = x_50878 & x_50881;
assign x_50883 = x_50875 & x_50882;
assign x_50884 = x_50869 & x_50883;
assign x_50885 = x_19592 & x_19593;
assign x_50886 = x_19591 & x_50885;
assign x_50887 = x_19594 & x_19595;
assign x_50888 = x_19596 & x_19597;
assign x_50889 = x_50887 & x_50888;
assign x_50890 = x_50886 & x_50889;
assign x_50891 = x_19598 & x_19599;
assign x_50892 = x_19600 & x_19601;
assign x_50893 = x_50891 & x_50892;
assign x_50894 = x_19602 & x_19603;
assign x_50895 = x_19604 & x_19605;
assign x_50896 = x_50894 & x_50895;
assign x_50897 = x_50893 & x_50896;
assign x_50898 = x_50890 & x_50897;
assign x_50899 = x_19606 & x_19607;
assign x_50900 = x_19608 & x_19609;
assign x_50901 = x_50899 & x_50900;
assign x_50902 = x_19610 & x_19611;
assign x_50903 = x_19612 & x_19613;
assign x_50904 = x_50902 & x_50903;
assign x_50905 = x_50901 & x_50904;
assign x_50906 = x_19614 & x_19615;
assign x_50907 = x_19616 & x_19617;
assign x_50908 = x_50906 & x_50907;
assign x_50909 = x_19618 & x_19619;
assign x_50910 = x_19620 & x_19621;
assign x_50911 = x_50909 & x_50910;
assign x_50912 = x_50908 & x_50911;
assign x_50913 = x_50905 & x_50912;
assign x_50914 = x_50898 & x_50913;
assign x_50915 = x_50884 & x_50914;
assign x_50916 = x_19623 & x_19624;
assign x_50917 = x_19622 & x_50916;
assign x_50918 = x_19625 & x_19626;
assign x_50919 = x_19627 & x_19628;
assign x_50920 = x_50918 & x_50919;
assign x_50921 = x_50917 & x_50920;
assign x_50922 = x_19629 & x_19630;
assign x_50923 = x_19631 & x_19632;
assign x_50924 = x_50922 & x_50923;
assign x_50925 = x_19633 & x_19634;
assign x_50926 = x_19635 & x_19636;
assign x_50927 = x_50925 & x_50926;
assign x_50928 = x_50924 & x_50927;
assign x_50929 = x_50921 & x_50928;
assign x_50930 = x_19638 & x_19639;
assign x_50931 = x_19637 & x_50930;
assign x_50932 = x_19640 & x_19641;
assign x_50933 = x_19642 & x_19643;
assign x_50934 = x_50932 & x_50933;
assign x_50935 = x_50931 & x_50934;
assign x_50936 = x_19644 & x_19645;
assign x_50937 = x_19646 & x_19647;
assign x_50938 = x_50936 & x_50937;
assign x_50939 = x_19648 & x_19649;
assign x_50940 = x_19650 & x_19651;
assign x_50941 = x_50939 & x_50940;
assign x_50942 = x_50938 & x_50941;
assign x_50943 = x_50935 & x_50942;
assign x_50944 = x_50929 & x_50943;
assign x_50945 = x_19653 & x_19654;
assign x_50946 = x_19652 & x_50945;
assign x_50947 = x_19655 & x_19656;
assign x_50948 = x_19657 & x_19658;
assign x_50949 = x_50947 & x_50948;
assign x_50950 = x_50946 & x_50949;
assign x_50951 = x_19659 & x_19660;
assign x_50952 = x_19661 & x_19662;
assign x_50953 = x_50951 & x_50952;
assign x_50954 = x_19663 & x_19664;
assign x_50955 = x_19665 & x_19666;
assign x_50956 = x_50954 & x_50955;
assign x_50957 = x_50953 & x_50956;
assign x_50958 = x_50950 & x_50957;
assign x_50959 = x_19667 & x_19668;
assign x_50960 = x_19669 & x_19670;
assign x_50961 = x_50959 & x_50960;
assign x_50962 = x_19671 & x_19672;
assign x_50963 = x_19673 & x_19674;
assign x_50964 = x_50962 & x_50963;
assign x_50965 = x_50961 & x_50964;
assign x_50966 = x_19675 & x_19676;
assign x_50967 = x_19677 & x_19678;
assign x_50968 = x_50966 & x_50967;
assign x_50969 = x_19679 & x_19680;
assign x_50970 = x_19681 & x_19682;
assign x_50971 = x_50969 & x_50970;
assign x_50972 = x_50968 & x_50971;
assign x_50973 = x_50965 & x_50972;
assign x_50974 = x_50958 & x_50973;
assign x_50975 = x_50944 & x_50974;
assign x_50976 = x_50915 & x_50975;
assign x_50977 = x_19684 & x_19685;
assign x_50978 = x_19683 & x_50977;
assign x_50979 = x_19686 & x_19687;
assign x_50980 = x_19688 & x_19689;
assign x_50981 = x_50979 & x_50980;
assign x_50982 = x_50978 & x_50981;
assign x_50983 = x_19690 & x_19691;
assign x_50984 = x_19692 & x_19693;
assign x_50985 = x_50983 & x_50984;
assign x_50986 = x_19694 & x_19695;
assign x_50987 = x_19696 & x_19697;
assign x_50988 = x_50986 & x_50987;
assign x_50989 = x_50985 & x_50988;
assign x_50990 = x_50982 & x_50989;
assign x_50991 = x_19699 & x_19700;
assign x_50992 = x_19698 & x_50991;
assign x_50993 = x_19701 & x_19702;
assign x_50994 = x_19703 & x_19704;
assign x_50995 = x_50993 & x_50994;
assign x_50996 = x_50992 & x_50995;
assign x_50997 = x_19705 & x_19706;
assign x_50998 = x_19707 & x_19708;
assign x_50999 = x_50997 & x_50998;
assign x_51000 = x_19709 & x_19710;
assign x_51001 = x_19711 & x_19712;
assign x_51002 = x_51000 & x_51001;
assign x_51003 = x_50999 & x_51002;
assign x_51004 = x_50996 & x_51003;
assign x_51005 = x_50990 & x_51004;
assign x_51006 = x_19714 & x_19715;
assign x_51007 = x_19713 & x_51006;
assign x_51008 = x_19716 & x_19717;
assign x_51009 = x_19718 & x_19719;
assign x_51010 = x_51008 & x_51009;
assign x_51011 = x_51007 & x_51010;
assign x_51012 = x_19720 & x_19721;
assign x_51013 = x_19722 & x_19723;
assign x_51014 = x_51012 & x_51013;
assign x_51015 = x_19724 & x_19725;
assign x_51016 = x_19726 & x_19727;
assign x_51017 = x_51015 & x_51016;
assign x_51018 = x_51014 & x_51017;
assign x_51019 = x_51011 & x_51018;
assign x_51020 = x_19728 & x_19729;
assign x_51021 = x_19730 & x_19731;
assign x_51022 = x_51020 & x_51021;
assign x_51023 = x_19732 & x_19733;
assign x_51024 = x_19734 & x_19735;
assign x_51025 = x_51023 & x_51024;
assign x_51026 = x_51022 & x_51025;
assign x_51027 = x_19736 & x_19737;
assign x_51028 = x_19738 & x_19739;
assign x_51029 = x_51027 & x_51028;
assign x_51030 = x_19740 & x_19741;
assign x_51031 = x_19742 & x_19743;
assign x_51032 = x_51030 & x_51031;
assign x_51033 = x_51029 & x_51032;
assign x_51034 = x_51026 & x_51033;
assign x_51035 = x_51019 & x_51034;
assign x_51036 = x_51005 & x_51035;
assign x_51037 = x_19745 & x_19746;
assign x_51038 = x_19744 & x_51037;
assign x_51039 = x_19747 & x_19748;
assign x_51040 = x_19749 & x_19750;
assign x_51041 = x_51039 & x_51040;
assign x_51042 = x_51038 & x_51041;
assign x_51043 = x_19751 & x_19752;
assign x_51044 = x_19753 & x_19754;
assign x_51045 = x_51043 & x_51044;
assign x_51046 = x_19755 & x_19756;
assign x_51047 = x_19757 & x_19758;
assign x_51048 = x_51046 & x_51047;
assign x_51049 = x_51045 & x_51048;
assign x_51050 = x_51042 & x_51049;
assign x_51051 = x_19760 & x_19761;
assign x_51052 = x_19759 & x_51051;
assign x_51053 = x_19762 & x_19763;
assign x_51054 = x_19764 & x_19765;
assign x_51055 = x_51053 & x_51054;
assign x_51056 = x_51052 & x_51055;
assign x_51057 = x_19766 & x_19767;
assign x_51058 = x_19768 & x_19769;
assign x_51059 = x_51057 & x_51058;
assign x_51060 = x_19770 & x_19771;
assign x_51061 = x_19772 & x_19773;
assign x_51062 = x_51060 & x_51061;
assign x_51063 = x_51059 & x_51062;
assign x_51064 = x_51056 & x_51063;
assign x_51065 = x_51050 & x_51064;
assign x_51066 = x_19775 & x_19776;
assign x_51067 = x_19774 & x_51066;
assign x_51068 = x_19777 & x_19778;
assign x_51069 = x_19779 & x_19780;
assign x_51070 = x_51068 & x_51069;
assign x_51071 = x_51067 & x_51070;
assign x_51072 = x_19781 & x_19782;
assign x_51073 = x_19783 & x_19784;
assign x_51074 = x_51072 & x_51073;
assign x_51075 = x_19785 & x_19786;
assign x_51076 = x_19787 & x_19788;
assign x_51077 = x_51075 & x_51076;
assign x_51078 = x_51074 & x_51077;
assign x_51079 = x_51071 & x_51078;
assign x_51080 = x_19789 & x_19790;
assign x_51081 = x_19791 & x_19792;
assign x_51082 = x_51080 & x_51081;
assign x_51083 = x_19793 & x_19794;
assign x_51084 = x_19795 & x_19796;
assign x_51085 = x_51083 & x_51084;
assign x_51086 = x_51082 & x_51085;
assign x_51087 = x_19797 & x_19798;
assign x_51088 = x_19799 & x_19800;
assign x_51089 = x_51087 & x_51088;
assign x_51090 = x_19801 & x_19802;
assign x_51091 = x_19803 & x_19804;
assign x_51092 = x_51090 & x_51091;
assign x_51093 = x_51089 & x_51092;
assign x_51094 = x_51086 & x_51093;
assign x_51095 = x_51079 & x_51094;
assign x_51096 = x_51065 & x_51095;
assign x_51097 = x_51036 & x_51096;
assign x_51098 = x_50976 & x_51097;
assign x_51099 = x_19806 & x_19807;
assign x_51100 = x_19805 & x_51099;
assign x_51101 = x_19808 & x_19809;
assign x_51102 = x_19810 & x_19811;
assign x_51103 = x_51101 & x_51102;
assign x_51104 = x_51100 & x_51103;
assign x_51105 = x_19812 & x_19813;
assign x_51106 = x_19814 & x_19815;
assign x_51107 = x_51105 & x_51106;
assign x_51108 = x_19816 & x_19817;
assign x_51109 = x_19818 & x_19819;
assign x_51110 = x_51108 & x_51109;
assign x_51111 = x_51107 & x_51110;
assign x_51112 = x_51104 & x_51111;
assign x_51113 = x_19821 & x_19822;
assign x_51114 = x_19820 & x_51113;
assign x_51115 = x_19823 & x_19824;
assign x_51116 = x_19825 & x_19826;
assign x_51117 = x_51115 & x_51116;
assign x_51118 = x_51114 & x_51117;
assign x_51119 = x_19827 & x_19828;
assign x_51120 = x_19829 & x_19830;
assign x_51121 = x_51119 & x_51120;
assign x_51122 = x_19831 & x_19832;
assign x_51123 = x_19833 & x_19834;
assign x_51124 = x_51122 & x_51123;
assign x_51125 = x_51121 & x_51124;
assign x_51126 = x_51118 & x_51125;
assign x_51127 = x_51112 & x_51126;
assign x_51128 = x_19836 & x_19837;
assign x_51129 = x_19835 & x_51128;
assign x_51130 = x_19838 & x_19839;
assign x_51131 = x_19840 & x_19841;
assign x_51132 = x_51130 & x_51131;
assign x_51133 = x_51129 & x_51132;
assign x_51134 = x_19842 & x_19843;
assign x_51135 = x_19844 & x_19845;
assign x_51136 = x_51134 & x_51135;
assign x_51137 = x_19846 & x_19847;
assign x_51138 = x_19848 & x_19849;
assign x_51139 = x_51137 & x_51138;
assign x_51140 = x_51136 & x_51139;
assign x_51141 = x_51133 & x_51140;
assign x_51142 = x_19850 & x_19851;
assign x_51143 = x_19852 & x_19853;
assign x_51144 = x_51142 & x_51143;
assign x_51145 = x_19854 & x_19855;
assign x_51146 = x_19856 & x_19857;
assign x_51147 = x_51145 & x_51146;
assign x_51148 = x_51144 & x_51147;
assign x_51149 = x_19858 & x_19859;
assign x_51150 = x_19860 & x_19861;
assign x_51151 = x_51149 & x_51150;
assign x_51152 = x_19862 & x_19863;
assign x_51153 = x_19864 & x_19865;
assign x_51154 = x_51152 & x_51153;
assign x_51155 = x_51151 & x_51154;
assign x_51156 = x_51148 & x_51155;
assign x_51157 = x_51141 & x_51156;
assign x_51158 = x_51127 & x_51157;
assign x_51159 = x_19867 & x_19868;
assign x_51160 = x_19866 & x_51159;
assign x_51161 = x_19869 & x_19870;
assign x_51162 = x_19871 & x_19872;
assign x_51163 = x_51161 & x_51162;
assign x_51164 = x_51160 & x_51163;
assign x_51165 = x_19873 & x_19874;
assign x_51166 = x_19875 & x_19876;
assign x_51167 = x_51165 & x_51166;
assign x_51168 = x_19877 & x_19878;
assign x_51169 = x_19879 & x_19880;
assign x_51170 = x_51168 & x_51169;
assign x_51171 = x_51167 & x_51170;
assign x_51172 = x_51164 & x_51171;
assign x_51173 = x_19882 & x_19883;
assign x_51174 = x_19881 & x_51173;
assign x_51175 = x_19884 & x_19885;
assign x_51176 = x_19886 & x_19887;
assign x_51177 = x_51175 & x_51176;
assign x_51178 = x_51174 & x_51177;
assign x_51179 = x_19888 & x_19889;
assign x_51180 = x_19890 & x_19891;
assign x_51181 = x_51179 & x_51180;
assign x_51182 = x_19892 & x_19893;
assign x_51183 = x_19894 & x_19895;
assign x_51184 = x_51182 & x_51183;
assign x_51185 = x_51181 & x_51184;
assign x_51186 = x_51178 & x_51185;
assign x_51187 = x_51172 & x_51186;
assign x_51188 = x_19897 & x_19898;
assign x_51189 = x_19896 & x_51188;
assign x_51190 = x_19899 & x_19900;
assign x_51191 = x_19901 & x_19902;
assign x_51192 = x_51190 & x_51191;
assign x_51193 = x_51189 & x_51192;
assign x_51194 = x_19903 & x_19904;
assign x_51195 = x_19905 & x_19906;
assign x_51196 = x_51194 & x_51195;
assign x_51197 = x_19907 & x_19908;
assign x_51198 = x_19909 & x_19910;
assign x_51199 = x_51197 & x_51198;
assign x_51200 = x_51196 & x_51199;
assign x_51201 = x_51193 & x_51200;
assign x_51202 = x_19911 & x_19912;
assign x_51203 = x_19913 & x_19914;
assign x_51204 = x_51202 & x_51203;
assign x_51205 = x_19915 & x_19916;
assign x_51206 = x_19917 & x_19918;
assign x_51207 = x_51205 & x_51206;
assign x_51208 = x_51204 & x_51207;
assign x_51209 = x_19919 & x_19920;
assign x_51210 = x_19921 & x_19922;
assign x_51211 = x_51209 & x_51210;
assign x_51212 = x_19923 & x_19924;
assign x_51213 = x_19925 & x_19926;
assign x_51214 = x_51212 & x_51213;
assign x_51215 = x_51211 & x_51214;
assign x_51216 = x_51208 & x_51215;
assign x_51217 = x_51201 & x_51216;
assign x_51218 = x_51187 & x_51217;
assign x_51219 = x_51158 & x_51218;
assign x_51220 = x_19928 & x_19929;
assign x_51221 = x_19927 & x_51220;
assign x_51222 = x_19930 & x_19931;
assign x_51223 = x_19932 & x_19933;
assign x_51224 = x_51222 & x_51223;
assign x_51225 = x_51221 & x_51224;
assign x_51226 = x_19934 & x_19935;
assign x_51227 = x_19936 & x_19937;
assign x_51228 = x_51226 & x_51227;
assign x_51229 = x_19938 & x_19939;
assign x_51230 = x_19940 & x_19941;
assign x_51231 = x_51229 & x_51230;
assign x_51232 = x_51228 & x_51231;
assign x_51233 = x_51225 & x_51232;
assign x_51234 = x_19943 & x_19944;
assign x_51235 = x_19942 & x_51234;
assign x_51236 = x_19945 & x_19946;
assign x_51237 = x_19947 & x_19948;
assign x_51238 = x_51236 & x_51237;
assign x_51239 = x_51235 & x_51238;
assign x_51240 = x_19949 & x_19950;
assign x_51241 = x_19951 & x_19952;
assign x_51242 = x_51240 & x_51241;
assign x_51243 = x_19953 & x_19954;
assign x_51244 = x_19955 & x_19956;
assign x_51245 = x_51243 & x_51244;
assign x_51246 = x_51242 & x_51245;
assign x_51247 = x_51239 & x_51246;
assign x_51248 = x_51233 & x_51247;
assign x_51249 = x_19958 & x_19959;
assign x_51250 = x_19957 & x_51249;
assign x_51251 = x_19960 & x_19961;
assign x_51252 = x_19962 & x_19963;
assign x_51253 = x_51251 & x_51252;
assign x_51254 = x_51250 & x_51253;
assign x_51255 = x_19964 & x_19965;
assign x_51256 = x_19966 & x_19967;
assign x_51257 = x_51255 & x_51256;
assign x_51258 = x_19968 & x_19969;
assign x_51259 = x_19970 & x_19971;
assign x_51260 = x_51258 & x_51259;
assign x_51261 = x_51257 & x_51260;
assign x_51262 = x_51254 & x_51261;
assign x_51263 = x_19972 & x_19973;
assign x_51264 = x_19974 & x_19975;
assign x_51265 = x_51263 & x_51264;
assign x_51266 = x_19976 & x_19977;
assign x_51267 = x_19978 & x_19979;
assign x_51268 = x_51266 & x_51267;
assign x_51269 = x_51265 & x_51268;
assign x_51270 = x_19980 & x_19981;
assign x_51271 = x_19982 & x_19983;
assign x_51272 = x_51270 & x_51271;
assign x_51273 = x_19984 & x_19985;
assign x_51274 = x_19986 & x_19987;
assign x_51275 = x_51273 & x_51274;
assign x_51276 = x_51272 & x_51275;
assign x_51277 = x_51269 & x_51276;
assign x_51278 = x_51262 & x_51277;
assign x_51279 = x_51248 & x_51278;
assign x_51280 = x_19989 & x_19990;
assign x_51281 = x_19988 & x_51280;
assign x_51282 = x_19991 & x_19992;
assign x_51283 = x_19993 & x_19994;
assign x_51284 = x_51282 & x_51283;
assign x_51285 = x_51281 & x_51284;
assign x_51286 = x_19995 & x_19996;
assign x_51287 = x_19997 & x_19998;
assign x_51288 = x_51286 & x_51287;
assign x_51289 = x_19999 & x_20000;
assign x_51290 = x_20001 & x_20002;
assign x_51291 = x_51289 & x_51290;
assign x_51292 = x_51288 & x_51291;
assign x_51293 = x_51285 & x_51292;
assign x_51294 = x_20003 & x_20004;
assign x_51295 = x_20005 & x_20006;
assign x_51296 = x_51294 & x_51295;
assign x_51297 = x_20007 & x_20008;
assign x_51298 = x_20009 & x_20010;
assign x_51299 = x_51297 & x_51298;
assign x_51300 = x_51296 & x_51299;
assign x_51301 = x_20011 & x_20012;
assign x_51302 = x_20013 & x_20014;
assign x_51303 = x_51301 & x_51302;
assign x_51304 = x_20015 & x_20016;
assign x_51305 = x_20017 & x_20018;
assign x_51306 = x_51304 & x_51305;
assign x_51307 = x_51303 & x_51306;
assign x_51308 = x_51300 & x_51307;
assign x_51309 = x_51293 & x_51308;
assign x_51310 = x_20020 & x_20021;
assign x_51311 = x_20019 & x_51310;
assign x_51312 = x_20022 & x_20023;
assign x_51313 = x_20024 & x_20025;
assign x_51314 = x_51312 & x_51313;
assign x_51315 = x_51311 & x_51314;
assign x_51316 = x_20026 & x_20027;
assign x_51317 = x_20028 & x_20029;
assign x_51318 = x_51316 & x_51317;
assign x_51319 = x_20030 & x_20031;
assign x_51320 = x_20032 & x_20033;
assign x_51321 = x_51319 & x_51320;
assign x_51322 = x_51318 & x_51321;
assign x_51323 = x_51315 & x_51322;
assign x_51324 = x_20034 & x_20035;
assign x_51325 = x_20036 & x_20037;
assign x_51326 = x_51324 & x_51325;
assign x_51327 = x_20038 & x_20039;
assign x_51328 = x_20040 & x_20041;
assign x_51329 = x_51327 & x_51328;
assign x_51330 = x_51326 & x_51329;
assign x_51331 = x_20042 & x_20043;
assign x_51332 = x_20044 & x_20045;
assign x_51333 = x_51331 & x_51332;
assign x_51334 = x_20046 & x_20047;
assign x_51335 = x_20048 & x_20049;
assign x_51336 = x_51334 & x_51335;
assign x_51337 = x_51333 & x_51336;
assign x_51338 = x_51330 & x_51337;
assign x_51339 = x_51323 & x_51338;
assign x_51340 = x_51309 & x_51339;
assign x_51341 = x_51279 & x_51340;
assign x_51342 = x_51219 & x_51341;
assign x_51343 = x_51098 & x_51342;
assign x_51344 = x_20051 & x_20052;
assign x_51345 = x_20050 & x_51344;
assign x_51346 = x_20053 & x_20054;
assign x_51347 = x_20055 & x_20056;
assign x_51348 = x_51346 & x_51347;
assign x_51349 = x_51345 & x_51348;
assign x_51350 = x_20057 & x_20058;
assign x_51351 = x_20059 & x_20060;
assign x_51352 = x_51350 & x_51351;
assign x_51353 = x_20061 & x_20062;
assign x_51354 = x_20063 & x_20064;
assign x_51355 = x_51353 & x_51354;
assign x_51356 = x_51352 & x_51355;
assign x_51357 = x_51349 & x_51356;
assign x_51358 = x_20066 & x_20067;
assign x_51359 = x_20065 & x_51358;
assign x_51360 = x_20068 & x_20069;
assign x_51361 = x_20070 & x_20071;
assign x_51362 = x_51360 & x_51361;
assign x_51363 = x_51359 & x_51362;
assign x_51364 = x_20072 & x_20073;
assign x_51365 = x_20074 & x_20075;
assign x_51366 = x_51364 & x_51365;
assign x_51367 = x_20076 & x_20077;
assign x_51368 = x_20078 & x_20079;
assign x_51369 = x_51367 & x_51368;
assign x_51370 = x_51366 & x_51369;
assign x_51371 = x_51363 & x_51370;
assign x_51372 = x_51357 & x_51371;
assign x_51373 = x_20081 & x_20082;
assign x_51374 = x_20080 & x_51373;
assign x_51375 = x_20083 & x_20084;
assign x_51376 = x_20085 & x_20086;
assign x_51377 = x_51375 & x_51376;
assign x_51378 = x_51374 & x_51377;
assign x_51379 = x_20087 & x_20088;
assign x_51380 = x_20089 & x_20090;
assign x_51381 = x_51379 & x_51380;
assign x_51382 = x_20091 & x_20092;
assign x_51383 = x_20093 & x_20094;
assign x_51384 = x_51382 & x_51383;
assign x_51385 = x_51381 & x_51384;
assign x_51386 = x_51378 & x_51385;
assign x_51387 = x_20095 & x_20096;
assign x_51388 = x_20097 & x_20098;
assign x_51389 = x_51387 & x_51388;
assign x_51390 = x_20099 & x_20100;
assign x_51391 = x_20101 & x_20102;
assign x_51392 = x_51390 & x_51391;
assign x_51393 = x_51389 & x_51392;
assign x_51394 = x_20103 & x_20104;
assign x_51395 = x_20105 & x_20106;
assign x_51396 = x_51394 & x_51395;
assign x_51397 = x_20107 & x_20108;
assign x_51398 = x_20109 & x_20110;
assign x_51399 = x_51397 & x_51398;
assign x_51400 = x_51396 & x_51399;
assign x_51401 = x_51393 & x_51400;
assign x_51402 = x_51386 & x_51401;
assign x_51403 = x_51372 & x_51402;
assign x_51404 = x_20112 & x_20113;
assign x_51405 = x_20111 & x_51404;
assign x_51406 = x_20114 & x_20115;
assign x_51407 = x_20116 & x_20117;
assign x_51408 = x_51406 & x_51407;
assign x_51409 = x_51405 & x_51408;
assign x_51410 = x_20118 & x_20119;
assign x_51411 = x_20120 & x_20121;
assign x_51412 = x_51410 & x_51411;
assign x_51413 = x_20122 & x_20123;
assign x_51414 = x_20124 & x_20125;
assign x_51415 = x_51413 & x_51414;
assign x_51416 = x_51412 & x_51415;
assign x_51417 = x_51409 & x_51416;
assign x_51418 = x_20127 & x_20128;
assign x_51419 = x_20126 & x_51418;
assign x_51420 = x_20129 & x_20130;
assign x_51421 = x_20131 & x_20132;
assign x_51422 = x_51420 & x_51421;
assign x_51423 = x_51419 & x_51422;
assign x_51424 = x_20133 & x_20134;
assign x_51425 = x_20135 & x_20136;
assign x_51426 = x_51424 & x_51425;
assign x_51427 = x_20137 & x_20138;
assign x_51428 = x_20139 & x_20140;
assign x_51429 = x_51427 & x_51428;
assign x_51430 = x_51426 & x_51429;
assign x_51431 = x_51423 & x_51430;
assign x_51432 = x_51417 & x_51431;
assign x_51433 = x_20142 & x_20143;
assign x_51434 = x_20141 & x_51433;
assign x_51435 = x_20144 & x_20145;
assign x_51436 = x_20146 & x_20147;
assign x_51437 = x_51435 & x_51436;
assign x_51438 = x_51434 & x_51437;
assign x_51439 = x_20148 & x_20149;
assign x_51440 = x_20150 & x_20151;
assign x_51441 = x_51439 & x_51440;
assign x_51442 = x_20152 & x_20153;
assign x_51443 = x_20154 & x_20155;
assign x_51444 = x_51442 & x_51443;
assign x_51445 = x_51441 & x_51444;
assign x_51446 = x_51438 & x_51445;
assign x_51447 = x_20156 & x_20157;
assign x_51448 = x_20158 & x_20159;
assign x_51449 = x_51447 & x_51448;
assign x_51450 = x_20160 & x_20161;
assign x_51451 = x_20162 & x_20163;
assign x_51452 = x_51450 & x_51451;
assign x_51453 = x_51449 & x_51452;
assign x_51454 = x_20164 & x_20165;
assign x_51455 = x_20166 & x_20167;
assign x_51456 = x_51454 & x_51455;
assign x_51457 = x_20168 & x_20169;
assign x_51458 = x_20170 & x_20171;
assign x_51459 = x_51457 & x_51458;
assign x_51460 = x_51456 & x_51459;
assign x_51461 = x_51453 & x_51460;
assign x_51462 = x_51446 & x_51461;
assign x_51463 = x_51432 & x_51462;
assign x_51464 = x_51403 & x_51463;
assign x_51465 = x_20173 & x_20174;
assign x_51466 = x_20172 & x_51465;
assign x_51467 = x_20175 & x_20176;
assign x_51468 = x_20177 & x_20178;
assign x_51469 = x_51467 & x_51468;
assign x_51470 = x_51466 & x_51469;
assign x_51471 = x_20179 & x_20180;
assign x_51472 = x_20181 & x_20182;
assign x_51473 = x_51471 & x_51472;
assign x_51474 = x_20183 & x_20184;
assign x_51475 = x_20185 & x_20186;
assign x_51476 = x_51474 & x_51475;
assign x_51477 = x_51473 & x_51476;
assign x_51478 = x_51470 & x_51477;
assign x_51479 = x_20188 & x_20189;
assign x_51480 = x_20187 & x_51479;
assign x_51481 = x_20190 & x_20191;
assign x_51482 = x_20192 & x_20193;
assign x_51483 = x_51481 & x_51482;
assign x_51484 = x_51480 & x_51483;
assign x_51485 = x_20194 & x_20195;
assign x_51486 = x_20196 & x_20197;
assign x_51487 = x_51485 & x_51486;
assign x_51488 = x_20198 & x_20199;
assign x_51489 = x_20200 & x_20201;
assign x_51490 = x_51488 & x_51489;
assign x_51491 = x_51487 & x_51490;
assign x_51492 = x_51484 & x_51491;
assign x_51493 = x_51478 & x_51492;
assign x_51494 = x_20203 & x_20204;
assign x_51495 = x_20202 & x_51494;
assign x_51496 = x_20205 & x_20206;
assign x_51497 = x_20207 & x_20208;
assign x_51498 = x_51496 & x_51497;
assign x_51499 = x_51495 & x_51498;
assign x_51500 = x_20209 & x_20210;
assign x_51501 = x_20211 & x_20212;
assign x_51502 = x_51500 & x_51501;
assign x_51503 = x_20213 & x_20214;
assign x_51504 = x_20215 & x_20216;
assign x_51505 = x_51503 & x_51504;
assign x_51506 = x_51502 & x_51505;
assign x_51507 = x_51499 & x_51506;
assign x_51508 = x_20217 & x_20218;
assign x_51509 = x_20219 & x_20220;
assign x_51510 = x_51508 & x_51509;
assign x_51511 = x_20221 & x_20222;
assign x_51512 = x_20223 & x_20224;
assign x_51513 = x_51511 & x_51512;
assign x_51514 = x_51510 & x_51513;
assign x_51515 = x_20225 & x_20226;
assign x_51516 = x_20227 & x_20228;
assign x_51517 = x_51515 & x_51516;
assign x_51518 = x_20229 & x_20230;
assign x_51519 = x_20231 & x_20232;
assign x_51520 = x_51518 & x_51519;
assign x_51521 = x_51517 & x_51520;
assign x_51522 = x_51514 & x_51521;
assign x_51523 = x_51507 & x_51522;
assign x_51524 = x_51493 & x_51523;
assign x_51525 = x_20234 & x_20235;
assign x_51526 = x_20233 & x_51525;
assign x_51527 = x_20236 & x_20237;
assign x_51528 = x_20238 & x_20239;
assign x_51529 = x_51527 & x_51528;
assign x_51530 = x_51526 & x_51529;
assign x_51531 = x_20240 & x_20241;
assign x_51532 = x_20242 & x_20243;
assign x_51533 = x_51531 & x_51532;
assign x_51534 = x_20244 & x_20245;
assign x_51535 = x_20246 & x_20247;
assign x_51536 = x_51534 & x_51535;
assign x_51537 = x_51533 & x_51536;
assign x_51538 = x_51530 & x_51537;
assign x_51539 = x_20249 & x_20250;
assign x_51540 = x_20248 & x_51539;
assign x_51541 = x_20251 & x_20252;
assign x_51542 = x_20253 & x_20254;
assign x_51543 = x_51541 & x_51542;
assign x_51544 = x_51540 & x_51543;
assign x_51545 = x_20255 & x_20256;
assign x_51546 = x_20257 & x_20258;
assign x_51547 = x_51545 & x_51546;
assign x_51548 = x_20259 & x_20260;
assign x_51549 = x_20261 & x_20262;
assign x_51550 = x_51548 & x_51549;
assign x_51551 = x_51547 & x_51550;
assign x_51552 = x_51544 & x_51551;
assign x_51553 = x_51538 & x_51552;
assign x_51554 = x_20264 & x_20265;
assign x_51555 = x_20263 & x_51554;
assign x_51556 = x_20266 & x_20267;
assign x_51557 = x_20268 & x_20269;
assign x_51558 = x_51556 & x_51557;
assign x_51559 = x_51555 & x_51558;
assign x_51560 = x_20270 & x_20271;
assign x_51561 = x_20272 & x_20273;
assign x_51562 = x_51560 & x_51561;
assign x_51563 = x_20274 & x_20275;
assign x_51564 = x_20276 & x_20277;
assign x_51565 = x_51563 & x_51564;
assign x_51566 = x_51562 & x_51565;
assign x_51567 = x_51559 & x_51566;
assign x_51568 = x_20278 & x_20279;
assign x_51569 = x_20280 & x_20281;
assign x_51570 = x_51568 & x_51569;
assign x_51571 = x_20282 & x_20283;
assign x_51572 = x_20284 & x_20285;
assign x_51573 = x_51571 & x_51572;
assign x_51574 = x_51570 & x_51573;
assign x_51575 = x_20286 & x_20287;
assign x_51576 = x_20288 & x_20289;
assign x_51577 = x_51575 & x_51576;
assign x_51578 = x_20290 & x_20291;
assign x_51579 = x_20292 & x_20293;
assign x_51580 = x_51578 & x_51579;
assign x_51581 = x_51577 & x_51580;
assign x_51582 = x_51574 & x_51581;
assign x_51583 = x_51567 & x_51582;
assign x_51584 = x_51553 & x_51583;
assign x_51585 = x_51524 & x_51584;
assign x_51586 = x_51464 & x_51585;
assign x_51587 = x_20295 & x_20296;
assign x_51588 = x_20294 & x_51587;
assign x_51589 = x_20297 & x_20298;
assign x_51590 = x_20299 & x_20300;
assign x_51591 = x_51589 & x_51590;
assign x_51592 = x_51588 & x_51591;
assign x_51593 = x_20301 & x_20302;
assign x_51594 = x_20303 & x_20304;
assign x_51595 = x_51593 & x_51594;
assign x_51596 = x_20305 & x_20306;
assign x_51597 = x_20307 & x_20308;
assign x_51598 = x_51596 & x_51597;
assign x_51599 = x_51595 & x_51598;
assign x_51600 = x_51592 & x_51599;
assign x_51601 = x_20310 & x_20311;
assign x_51602 = x_20309 & x_51601;
assign x_51603 = x_20312 & x_20313;
assign x_51604 = x_20314 & x_20315;
assign x_51605 = x_51603 & x_51604;
assign x_51606 = x_51602 & x_51605;
assign x_51607 = x_20316 & x_20317;
assign x_51608 = x_20318 & x_20319;
assign x_51609 = x_51607 & x_51608;
assign x_51610 = x_20320 & x_20321;
assign x_51611 = x_20322 & x_20323;
assign x_51612 = x_51610 & x_51611;
assign x_51613 = x_51609 & x_51612;
assign x_51614 = x_51606 & x_51613;
assign x_51615 = x_51600 & x_51614;
assign x_51616 = x_20325 & x_20326;
assign x_51617 = x_20324 & x_51616;
assign x_51618 = x_20327 & x_20328;
assign x_51619 = x_20329 & x_20330;
assign x_51620 = x_51618 & x_51619;
assign x_51621 = x_51617 & x_51620;
assign x_51622 = x_20331 & x_20332;
assign x_51623 = x_20333 & x_20334;
assign x_51624 = x_51622 & x_51623;
assign x_51625 = x_20335 & x_20336;
assign x_51626 = x_20337 & x_20338;
assign x_51627 = x_51625 & x_51626;
assign x_51628 = x_51624 & x_51627;
assign x_51629 = x_51621 & x_51628;
assign x_51630 = x_20339 & x_20340;
assign x_51631 = x_20341 & x_20342;
assign x_51632 = x_51630 & x_51631;
assign x_51633 = x_20343 & x_20344;
assign x_51634 = x_20345 & x_20346;
assign x_51635 = x_51633 & x_51634;
assign x_51636 = x_51632 & x_51635;
assign x_51637 = x_20347 & x_20348;
assign x_51638 = x_20349 & x_20350;
assign x_51639 = x_51637 & x_51638;
assign x_51640 = x_20351 & x_20352;
assign x_51641 = x_20353 & x_20354;
assign x_51642 = x_51640 & x_51641;
assign x_51643 = x_51639 & x_51642;
assign x_51644 = x_51636 & x_51643;
assign x_51645 = x_51629 & x_51644;
assign x_51646 = x_51615 & x_51645;
assign x_51647 = x_20356 & x_20357;
assign x_51648 = x_20355 & x_51647;
assign x_51649 = x_20358 & x_20359;
assign x_51650 = x_20360 & x_20361;
assign x_51651 = x_51649 & x_51650;
assign x_51652 = x_51648 & x_51651;
assign x_51653 = x_20362 & x_20363;
assign x_51654 = x_20364 & x_20365;
assign x_51655 = x_51653 & x_51654;
assign x_51656 = x_20366 & x_20367;
assign x_51657 = x_20368 & x_20369;
assign x_51658 = x_51656 & x_51657;
assign x_51659 = x_51655 & x_51658;
assign x_51660 = x_51652 & x_51659;
assign x_51661 = x_20371 & x_20372;
assign x_51662 = x_20370 & x_51661;
assign x_51663 = x_20373 & x_20374;
assign x_51664 = x_20375 & x_20376;
assign x_51665 = x_51663 & x_51664;
assign x_51666 = x_51662 & x_51665;
assign x_51667 = x_20377 & x_20378;
assign x_51668 = x_20379 & x_20380;
assign x_51669 = x_51667 & x_51668;
assign x_51670 = x_20381 & x_20382;
assign x_51671 = x_20383 & x_20384;
assign x_51672 = x_51670 & x_51671;
assign x_51673 = x_51669 & x_51672;
assign x_51674 = x_51666 & x_51673;
assign x_51675 = x_51660 & x_51674;
assign x_51676 = x_20386 & x_20387;
assign x_51677 = x_20385 & x_51676;
assign x_51678 = x_20388 & x_20389;
assign x_51679 = x_20390 & x_20391;
assign x_51680 = x_51678 & x_51679;
assign x_51681 = x_51677 & x_51680;
assign x_51682 = x_20392 & x_20393;
assign x_51683 = x_20394 & x_20395;
assign x_51684 = x_51682 & x_51683;
assign x_51685 = x_20396 & x_20397;
assign x_51686 = x_20398 & x_20399;
assign x_51687 = x_51685 & x_51686;
assign x_51688 = x_51684 & x_51687;
assign x_51689 = x_51681 & x_51688;
assign x_51690 = x_20400 & x_20401;
assign x_51691 = x_20402 & x_20403;
assign x_51692 = x_51690 & x_51691;
assign x_51693 = x_20404 & x_20405;
assign x_51694 = x_20406 & x_20407;
assign x_51695 = x_51693 & x_51694;
assign x_51696 = x_51692 & x_51695;
assign x_51697 = x_20408 & x_20409;
assign x_51698 = x_20410 & x_20411;
assign x_51699 = x_51697 & x_51698;
assign x_51700 = x_20412 & x_20413;
assign x_51701 = x_20414 & x_20415;
assign x_51702 = x_51700 & x_51701;
assign x_51703 = x_51699 & x_51702;
assign x_51704 = x_51696 & x_51703;
assign x_51705 = x_51689 & x_51704;
assign x_51706 = x_51675 & x_51705;
assign x_51707 = x_51646 & x_51706;
assign x_51708 = x_20417 & x_20418;
assign x_51709 = x_20416 & x_51708;
assign x_51710 = x_20419 & x_20420;
assign x_51711 = x_20421 & x_20422;
assign x_51712 = x_51710 & x_51711;
assign x_51713 = x_51709 & x_51712;
assign x_51714 = x_20423 & x_20424;
assign x_51715 = x_20425 & x_20426;
assign x_51716 = x_51714 & x_51715;
assign x_51717 = x_20427 & x_20428;
assign x_51718 = x_20429 & x_20430;
assign x_51719 = x_51717 & x_51718;
assign x_51720 = x_51716 & x_51719;
assign x_51721 = x_51713 & x_51720;
assign x_51722 = x_20432 & x_20433;
assign x_51723 = x_20431 & x_51722;
assign x_51724 = x_20434 & x_20435;
assign x_51725 = x_20436 & x_20437;
assign x_51726 = x_51724 & x_51725;
assign x_51727 = x_51723 & x_51726;
assign x_51728 = x_20438 & x_20439;
assign x_51729 = x_20440 & x_20441;
assign x_51730 = x_51728 & x_51729;
assign x_51731 = x_20442 & x_20443;
assign x_51732 = x_20444 & x_20445;
assign x_51733 = x_51731 & x_51732;
assign x_51734 = x_51730 & x_51733;
assign x_51735 = x_51727 & x_51734;
assign x_51736 = x_51721 & x_51735;
assign x_51737 = x_20447 & x_20448;
assign x_51738 = x_20446 & x_51737;
assign x_51739 = x_20449 & x_20450;
assign x_51740 = x_20451 & x_20452;
assign x_51741 = x_51739 & x_51740;
assign x_51742 = x_51738 & x_51741;
assign x_51743 = x_20453 & x_20454;
assign x_51744 = x_20455 & x_20456;
assign x_51745 = x_51743 & x_51744;
assign x_51746 = x_20457 & x_20458;
assign x_51747 = x_20459 & x_20460;
assign x_51748 = x_51746 & x_51747;
assign x_51749 = x_51745 & x_51748;
assign x_51750 = x_51742 & x_51749;
assign x_51751 = x_20461 & x_20462;
assign x_51752 = x_20463 & x_20464;
assign x_51753 = x_51751 & x_51752;
assign x_51754 = x_20465 & x_20466;
assign x_51755 = x_20467 & x_20468;
assign x_51756 = x_51754 & x_51755;
assign x_51757 = x_51753 & x_51756;
assign x_51758 = x_20469 & x_20470;
assign x_51759 = x_20471 & x_20472;
assign x_51760 = x_51758 & x_51759;
assign x_51761 = x_20473 & x_20474;
assign x_51762 = x_20475 & x_20476;
assign x_51763 = x_51761 & x_51762;
assign x_51764 = x_51760 & x_51763;
assign x_51765 = x_51757 & x_51764;
assign x_51766 = x_51750 & x_51765;
assign x_51767 = x_51736 & x_51766;
assign x_51768 = x_20478 & x_20479;
assign x_51769 = x_20477 & x_51768;
assign x_51770 = x_20480 & x_20481;
assign x_51771 = x_20482 & x_20483;
assign x_51772 = x_51770 & x_51771;
assign x_51773 = x_51769 & x_51772;
assign x_51774 = x_20484 & x_20485;
assign x_51775 = x_20486 & x_20487;
assign x_51776 = x_51774 & x_51775;
assign x_51777 = x_20488 & x_20489;
assign x_51778 = x_20490 & x_20491;
assign x_51779 = x_51777 & x_51778;
assign x_51780 = x_51776 & x_51779;
assign x_51781 = x_51773 & x_51780;
assign x_51782 = x_20492 & x_20493;
assign x_51783 = x_20494 & x_20495;
assign x_51784 = x_51782 & x_51783;
assign x_51785 = x_20496 & x_20497;
assign x_51786 = x_20498 & x_20499;
assign x_51787 = x_51785 & x_51786;
assign x_51788 = x_51784 & x_51787;
assign x_51789 = x_20500 & x_20501;
assign x_51790 = x_20502 & x_20503;
assign x_51791 = x_51789 & x_51790;
assign x_51792 = x_20504 & x_20505;
assign x_51793 = x_20506 & x_20507;
assign x_51794 = x_51792 & x_51793;
assign x_51795 = x_51791 & x_51794;
assign x_51796 = x_51788 & x_51795;
assign x_51797 = x_51781 & x_51796;
assign x_51798 = x_20509 & x_20510;
assign x_51799 = x_20508 & x_51798;
assign x_51800 = x_20511 & x_20512;
assign x_51801 = x_20513 & x_20514;
assign x_51802 = x_51800 & x_51801;
assign x_51803 = x_51799 & x_51802;
assign x_51804 = x_20515 & x_20516;
assign x_51805 = x_20517 & x_20518;
assign x_51806 = x_51804 & x_51805;
assign x_51807 = x_20519 & x_20520;
assign x_51808 = x_20521 & x_20522;
assign x_51809 = x_51807 & x_51808;
assign x_51810 = x_51806 & x_51809;
assign x_51811 = x_51803 & x_51810;
assign x_51812 = x_20523 & x_20524;
assign x_51813 = x_20525 & x_20526;
assign x_51814 = x_51812 & x_51813;
assign x_51815 = x_20527 & x_20528;
assign x_51816 = x_20529 & x_20530;
assign x_51817 = x_51815 & x_51816;
assign x_51818 = x_51814 & x_51817;
assign x_51819 = x_20531 & x_20532;
assign x_51820 = x_20533 & x_20534;
assign x_51821 = x_51819 & x_51820;
assign x_51822 = x_20535 & x_20536;
assign x_51823 = x_20537 & x_20538;
assign x_51824 = x_51822 & x_51823;
assign x_51825 = x_51821 & x_51824;
assign x_51826 = x_51818 & x_51825;
assign x_51827 = x_51811 & x_51826;
assign x_51828 = x_51797 & x_51827;
assign x_51829 = x_51767 & x_51828;
assign x_51830 = x_51707 & x_51829;
assign x_51831 = x_51586 & x_51830;
assign x_51832 = x_51343 & x_51831;
assign x_51833 = x_20540 & x_20541;
assign x_51834 = x_20539 & x_51833;
assign x_51835 = x_20542 & x_20543;
assign x_51836 = x_20544 & x_20545;
assign x_51837 = x_51835 & x_51836;
assign x_51838 = x_51834 & x_51837;
assign x_51839 = x_20546 & x_20547;
assign x_51840 = x_20548 & x_20549;
assign x_51841 = x_51839 & x_51840;
assign x_51842 = x_20550 & x_20551;
assign x_51843 = x_20552 & x_20553;
assign x_51844 = x_51842 & x_51843;
assign x_51845 = x_51841 & x_51844;
assign x_51846 = x_51838 & x_51845;
assign x_51847 = x_20555 & x_20556;
assign x_51848 = x_20554 & x_51847;
assign x_51849 = x_20557 & x_20558;
assign x_51850 = x_20559 & x_20560;
assign x_51851 = x_51849 & x_51850;
assign x_51852 = x_51848 & x_51851;
assign x_51853 = x_20561 & x_20562;
assign x_51854 = x_20563 & x_20564;
assign x_51855 = x_51853 & x_51854;
assign x_51856 = x_20565 & x_20566;
assign x_51857 = x_20567 & x_20568;
assign x_51858 = x_51856 & x_51857;
assign x_51859 = x_51855 & x_51858;
assign x_51860 = x_51852 & x_51859;
assign x_51861 = x_51846 & x_51860;
assign x_51862 = x_20570 & x_20571;
assign x_51863 = x_20569 & x_51862;
assign x_51864 = x_20572 & x_20573;
assign x_51865 = x_20574 & x_20575;
assign x_51866 = x_51864 & x_51865;
assign x_51867 = x_51863 & x_51866;
assign x_51868 = x_20576 & x_20577;
assign x_51869 = x_20578 & x_20579;
assign x_51870 = x_51868 & x_51869;
assign x_51871 = x_20580 & x_20581;
assign x_51872 = x_20582 & x_20583;
assign x_51873 = x_51871 & x_51872;
assign x_51874 = x_51870 & x_51873;
assign x_51875 = x_51867 & x_51874;
assign x_51876 = x_20584 & x_20585;
assign x_51877 = x_20586 & x_20587;
assign x_51878 = x_51876 & x_51877;
assign x_51879 = x_20588 & x_20589;
assign x_51880 = x_20590 & x_20591;
assign x_51881 = x_51879 & x_51880;
assign x_51882 = x_51878 & x_51881;
assign x_51883 = x_20592 & x_20593;
assign x_51884 = x_20594 & x_20595;
assign x_51885 = x_51883 & x_51884;
assign x_51886 = x_20596 & x_20597;
assign x_51887 = x_20598 & x_20599;
assign x_51888 = x_51886 & x_51887;
assign x_51889 = x_51885 & x_51888;
assign x_51890 = x_51882 & x_51889;
assign x_51891 = x_51875 & x_51890;
assign x_51892 = x_51861 & x_51891;
assign x_51893 = x_20601 & x_20602;
assign x_51894 = x_20600 & x_51893;
assign x_51895 = x_20603 & x_20604;
assign x_51896 = x_20605 & x_20606;
assign x_51897 = x_51895 & x_51896;
assign x_51898 = x_51894 & x_51897;
assign x_51899 = x_20607 & x_20608;
assign x_51900 = x_20609 & x_20610;
assign x_51901 = x_51899 & x_51900;
assign x_51902 = x_20611 & x_20612;
assign x_51903 = x_20613 & x_20614;
assign x_51904 = x_51902 & x_51903;
assign x_51905 = x_51901 & x_51904;
assign x_51906 = x_51898 & x_51905;
assign x_51907 = x_20616 & x_20617;
assign x_51908 = x_20615 & x_51907;
assign x_51909 = x_20618 & x_20619;
assign x_51910 = x_20620 & x_20621;
assign x_51911 = x_51909 & x_51910;
assign x_51912 = x_51908 & x_51911;
assign x_51913 = x_20622 & x_20623;
assign x_51914 = x_20624 & x_20625;
assign x_51915 = x_51913 & x_51914;
assign x_51916 = x_20626 & x_20627;
assign x_51917 = x_20628 & x_20629;
assign x_51918 = x_51916 & x_51917;
assign x_51919 = x_51915 & x_51918;
assign x_51920 = x_51912 & x_51919;
assign x_51921 = x_51906 & x_51920;
assign x_51922 = x_20631 & x_20632;
assign x_51923 = x_20630 & x_51922;
assign x_51924 = x_20633 & x_20634;
assign x_51925 = x_20635 & x_20636;
assign x_51926 = x_51924 & x_51925;
assign x_51927 = x_51923 & x_51926;
assign x_51928 = x_20637 & x_20638;
assign x_51929 = x_20639 & x_20640;
assign x_51930 = x_51928 & x_51929;
assign x_51931 = x_20641 & x_20642;
assign x_51932 = x_20643 & x_20644;
assign x_51933 = x_51931 & x_51932;
assign x_51934 = x_51930 & x_51933;
assign x_51935 = x_51927 & x_51934;
assign x_51936 = x_20645 & x_20646;
assign x_51937 = x_20647 & x_20648;
assign x_51938 = x_51936 & x_51937;
assign x_51939 = x_20649 & x_20650;
assign x_51940 = x_20651 & x_20652;
assign x_51941 = x_51939 & x_51940;
assign x_51942 = x_51938 & x_51941;
assign x_51943 = x_20653 & x_20654;
assign x_51944 = x_20655 & x_20656;
assign x_51945 = x_51943 & x_51944;
assign x_51946 = x_20657 & x_20658;
assign x_51947 = x_20659 & x_20660;
assign x_51948 = x_51946 & x_51947;
assign x_51949 = x_51945 & x_51948;
assign x_51950 = x_51942 & x_51949;
assign x_51951 = x_51935 & x_51950;
assign x_51952 = x_51921 & x_51951;
assign x_51953 = x_51892 & x_51952;
assign x_51954 = x_20662 & x_20663;
assign x_51955 = x_20661 & x_51954;
assign x_51956 = x_20664 & x_20665;
assign x_51957 = x_20666 & x_20667;
assign x_51958 = x_51956 & x_51957;
assign x_51959 = x_51955 & x_51958;
assign x_51960 = x_20668 & x_20669;
assign x_51961 = x_20670 & x_20671;
assign x_51962 = x_51960 & x_51961;
assign x_51963 = x_20672 & x_20673;
assign x_51964 = x_20674 & x_20675;
assign x_51965 = x_51963 & x_51964;
assign x_51966 = x_51962 & x_51965;
assign x_51967 = x_51959 & x_51966;
assign x_51968 = x_20677 & x_20678;
assign x_51969 = x_20676 & x_51968;
assign x_51970 = x_20679 & x_20680;
assign x_51971 = x_20681 & x_20682;
assign x_51972 = x_51970 & x_51971;
assign x_51973 = x_51969 & x_51972;
assign x_51974 = x_20683 & x_20684;
assign x_51975 = x_20685 & x_20686;
assign x_51976 = x_51974 & x_51975;
assign x_51977 = x_20687 & x_20688;
assign x_51978 = x_20689 & x_20690;
assign x_51979 = x_51977 & x_51978;
assign x_51980 = x_51976 & x_51979;
assign x_51981 = x_51973 & x_51980;
assign x_51982 = x_51967 & x_51981;
assign x_51983 = x_20692 & x_20693;
assign x_51984 = x_20691 & x_51983;
assign x_51985 = x_20694 & x_20695;
assign x_51986 = x_20696 & x_20697;
assign x_51987 = x_51985 & x_51986;
assign x_51988 = x_51984 & x_51987;
assign x_51989 = x_20698 & x_20699;
assign x_51990 = x_20700 & x_20701;
assign x_51991 = x_51989 & x_51990;
assign x_51992 = x_20702 & x_20703;
assign x_51993 = x_20704 & x_20705;
assign x_51994 = x_51992 & x_51993;
assign x_51995 = x_51991 & x_51994;
assign x_51996 = x_51988 & x_51995;
assign x_51997 = x_20706 & x_20707;
assign x_51998 = x_20708 & x_20709;
assign x_51999 = x_51997 & x_51998;
assign x_52000 = x_20710 & x_20711;
assign x_52001 = x_20712 & x_20713;
assign x_52002 = x_52000 & x_52001;
assign x_52003 = x_51999 & x_52002;
assign x_52004 = x_20714 & x_20715;
assign x_52005 = x_20716 & x_20717;
assign x_52006 = x_52004 & x_52005;
assign x_52007 = x_20718 & x_20719;
assign x_52008 = x_20720 & x_20721;
assign x_52009 = x_52007 & x_52008;
assign x_52010 = x_52006 & x_52009;
assign x_52011 = x_52003 & x_52010;
assign x_52012 = x_51996 & x_52011;
assign x_52013 = x_51982 & x_52012;
assign x_52014 = x_20723 & x_20724;
assign x_52015 = x_20722 & x_52014;
assign x_52016 = x_20725 & x_20726;
assign x_52017 = x_20727 & x_20728;
assign x_52018 = x_52016 & x_52017;
assign x_52019 = x_52015 & x_52018;
assign x_52020 = x_20729 & x_20730;
assign x_52021 = x_20731 & x_20732;
assign x_52022 = x_52020 & x_52021;
assign x_52023 = x_20733 & x_20734;
assign x_52024 = x_20735 & x_20736;
assign x_52025 = x_52023 & x_52024;
assign x_52026 = x_52022 & x_52025;
assign x_52027 = x_52019 & x_52026;
assign x_52028 = x_20738 & x_20739;
assign x_52029 = x_20737 & x_52028;
assign x_52030 = x_20740 & x_20741;
assign x_52031 = x_20742 & x_20743;
assign x_52032 = x_52030 & x_52031;
assign x_52033 = x_52029 & x_52032;
assign x_52034 = x_20744 & x_20745;
assign x_52035 = x_20746 & x_20747;
assign x_52036 = x_52034 & x_52035;
assign x_52037 = x_20748 & x_20749;
assign x_52038 = x_20750 & x_20751;
assign x_52039 = x_52037 & x_52038;
assign x_52040 = x_52036 & x_52039;
assign x_52041 = x_52033 & x_52040;
assign x_52042 = x_52027 & x_52041;
assign x_52043 = x_20753 & x_20754;
assign x_52044 = x_20752 & x_52043;
assign x_52045 = x_20755 & x_20756;
assign x_52046 = x_20757 & x_20758;
assign x_52047 = x_52045 & x_52046;
assign x_52048 = x_52044 & x_52047;
assign x_52049 = x_20759 & x_20760;
assign x_52050 = x_20761 & x_20762;
assign x_52051 = x_52049 & x_52050;
assign x_52052 = x_20763 & x_20764;
assign x_52053 = x_20765 & x_20766;
assign x_52054 = x_52052 & x_52053;
assign x_52055 = x_52051 & x_52054;
assign x_52056 = x_52048 & x_52055;
assign x_52057 = x_20767 & x_20768;
assign x_52058 = x_20769 & x_20770;
assign x_52059 = x_52057 & x_52058;
assign x_52060 = x_20771 & x_20772;
assign x_52061 = x_20773 & x_20774;
assign x_52062 = x_52060 & x_52061;
assign x_52063 = x_52059 & x_52062;
assign x_52064 = x_20775 & x_20776;
assign x_52065 = x_20777 & x_20778;
assign x_52066 = x_52064 & x_52065;
assign x_52067 = x_20779 & x_20780;
assign x_52068 = x_20781 & x_20782;
assign x_52069 = x_52067 & x_52068;
assign x_52070 = x_52066 & x_52069;
assign x_52071 = x_52063 & x_52070;
assign x_52072 = x_52056 & x_52071;
assign x_52073 = x_52042 & x_52072;
assign x_52074 = x_52013 & x_52073;
assign x_52075 = x_51953 & x_52074;
assign x_52076 = x_20784 & x_20785;
assign x_52077 = x_20783 & x_52076;
assign x_52078 = x_20786 & x_20787;
assign x_52079 = x_20788 & x_20789;
assign x_52080 = x_52078 & x_52079;
assign x_52081 = x_52077 & x_52080;
assign x_52082 = x_20790 & x_20791;
assign x_52083 = x_20792 & x_20793;
assign x_52084 = x_52082 & x_52083;
assign x_52085 = x_20794 & x_20795;
assign x_52086 = x_20796 & x_20797;
assign x_52087 = x_52085 & x_52086;
assign x_52088 = x_52084 & x_52087;
assign x_52089 = x_52081 & x_52088;
assign x_52090 = x_20799 & x_20800;
assign x_52091 = x_20798 & x_52090;
assign x_52092 = x_20801 & x_20802;
assign x_52093 = x_20803 & x_20804;
assign x_52094 = x_52092 & x_52093;
assign x_52095 = x_52091 & x_52094;
assign x_52096 = x_20805 & x_20806;
assign x_52097 = x_20807 & x_20808;
assign x_52098 = x_52096 & x_52097;
assign x_52099 = x_20809 & x_20810;
assign x_52100 = x_20811 & x_20812;
assign x_52101 = x_52099 & x_52100;
assign x_52102 = x_52098 & x_52101;
assign x_52103 = x_52095 & x_52102;
assign x_52104 = x_52089 & x_52103;
assign x_52105 = x_20814 & x_20815;
assign x_52106 = x_20813 & x_52105;
assign x_52107 = x_20816 & x_20817;
assign x_52108 = x_20818 & x_20819;
assign x_52109 = x_52107 & x_52108;
assign x_52110 = x_52106 & x_52109;
assign x_52111 = x_20820 & x_20821;
assign x_52112 = x_20822 & x_20823;
assign x_52113 = x_52111 & x_52112;
assign x_52114 = x_20824 & x_20825;
assign x_52115 = x_20826 & x_20827;
assign x_52116 = x_52114 & x_52115;
assign x_52117 = x_52113 & x_52116;
assign x_52118 = x_52110 & x_52117;
assign x_52119 = x_20828 & x_20829;
assign x_52120 = x_20830 & x_20831;
assign x_52121 = x_52119 & x_52120;
assign x_52122 = x_20832 & x_20833;
assign x_52123 = x_20834 & x_20835;
assign x_52124 = x_52122 & x_52123;
assign x_52125 = x_52121 & x_52124;
assign x_52126 = x_20836 & x_20837;
assign x_52127 = x_20838 & x_20839;
assign x_52128 = x_52126 & x_52127;
assign x_52129 = x_20840 & x_20841;
assign x_52130 = x_20842 & x_20843;
assign x_52131 = x_52129 & x_52130;
assign x_52132 = x_52128 & x_52131;
assign x_52133 = x_52125 & x_52132;
assign x_52134 = x_52118 & x_52133;
assign x_52135 = x_52104 & x_52134;
assign x_52136 = x_20845 & x_20846;
assign x_52137 = x_20844 & x_52136;
assign x_52138 = x_20847 & x_20848;
assign x_52139 = x_20849 & x_20850;
assign x_52140 = x_52138 & x_52139;
assign x_52141 = x_52137 & x_52140;
assign x_52142 = x_20851 & x_20852;
assign x_52143 = x_20853 & x_20854;
assign x_52144 = x_52142 & x_52143;
assign x_52145 = x_20855 & x_20856;
assign x_52146 = x_20857 & x_20858;
assign x_52147 = x_52145 & x_52146;
assign x_52148 = x_52144 & x_52147;
assign x_52149 = x_52141 & x_52148;
assign x_52150 = x_20860 & x_20861;
assign x_52151 = x_20859 & x_52150;
assign x_52152 = x_20862 & x_20863;
assign x_52153 = x_20864 & x_20865;
assign x_52154 = x_52152 & x_52153;
assign x_52155 = x_52151 & x_52154;
assign x_52156 = x_20866 & x_20867;
assign x_52157 = x_20868 & x_20869;
assign x_52158 = x_52156 & x_52157;
assign x_52159 = x_20870 & x_20871;
assign x_52160 = x_20872 & x_20873;
assign x_52161 = x_52159 & x_52160;
assign x_52162 = x_52158 & x_52161;
assign x_52163 = x_52155 & x_52162;
assign x_52164 = x_52149 & x_52163;
assign x_52165 = x_20875 & x_20876;
assign x_52166 = x_20874 & x_52165;
assign x_52167 = x_20877 & x_20878;
assign x_52168 = x_20879 & x_20880;
assign x_52169 = x_52167 & x_52168;
assign x_52170 = x_52166 & x_52169;
assign x_52171 = x_20881 & x_20882;
assign x_52172 = x_20883 & x_20884;
assign x_52173 = x_52171 & x_52172;
assign x_52174 = x_20885 & x_20886;
assign x_52175 = x_20887 & x_20888;
assign x_52176 = x_52174 & x_52175;
assign x_52177 = x_52173 & x_52176;
assign x_52178 = x_52170 & x_52177;
assign x_52179 = x_20889 & x_20890;
assign x_52180 = x_20891 & x_20892;
assign x_52181 = x_52179 & x_52180;
assign x_52182 = x_20893 & x_20894;
assign x_52183 = x_20895 & x_20896;
assign x_52184 = x_52182 & x_52183;
assign x_52185 = x_52181 & x_52184;
assign x_52186 = x_20897 & x_20898;
assign x_52187 = x_20899 & x_20900;
assign x_52188 = x_52186 & x_52187;
assign x_52189 = x_20901 & x_20902;
assign x_52190 = x_20903 & x_20904;
assign x_52191 = x_52189 & x_52190;
assign x_52192 = x_52188 & x_52191;
assign x_52193 = x_52185 & x_52192;
assign x_52194 = x_52178 & x_52193;
assign x_52195 = x_52164 & x_52194;
assign x_52196 = x_52135 & x_52195;
assign x_52197 = x_20906 & x_20907;
assign x_52198 = x_20905 & x_52197;
assign x_52199 = x_20908 & x_20909;
assign x_52200 = x_20910 & x_20911;
assign x_52201 = x_52199 & x_52200;
assign x_52202 = x_52198 & x_52201;
assign x_52203 = x_20912 & x_20913;
assign x_52204 = x_20914 & x_20915;
assign x_52205 = x_52203 & x_52204;
assign x_52206 = x_20916 & x_20917;
assign x_52207 = x_20918 & x_20919;
assign x_52208 = x_52206 & x_52207;
assign x_52209 = x_52205 & x_52208;
assign x_52210 = x_52202 & x_52209;
assign x_52211 = x_20921 & x_20922;
assign x_52212 = x_20920 & x_52211;
assign x_52213 = x_20923 & x_20924;
assign x_52214 = x_20925 & x_20926;
assign x_52215 = x_52213 & x_52214;
assign x_52216 = x_52212 & x_52215;
assign x_52217 = x_20927 & x_20928;
assign x_52218 = x_20929 & x_20930;
assign x_52219 = x_52217 & x_52218;
assign x_52220 = x_20931 & x_20932;
assign x_52221 = x_20933 & x_20934;
assign x_52222 = x_52220 & x_52221;
assign x_52223 = x_52219 & x_52222;
assign x_52224 = x_52216 & x_52223;
assign x_52225 = x_52210 & x_52224;
assign x_52226 = x_20936 & x_20937;
assign x_52227 = x_20935 & x_52226;
assign x_52228 = x_20938 & x_20939;
assign x_52229 = x_20940 & x_20941;
assign x_52230 = x_52228 & x_52229;
assign x_52231 = x_52227 & x_52230;
assign x_52232 = x_20942 & x_20943;
assign x_52233 = x_20944 & x_20945;
assign x_52234 = x_52232 & x_52233;
assign x_52235 = x_20946 & x_20947;
assign x_52236 = x_20948 & x_20949;
assign x_52237 = x_52235 & x_52236;
assign x_52238 = x_52234 & x_52237;
assign x_52239 = x_52231 & x_52238;
assign x_52240 = x_20950 & x_20951;
assign x_52241 = x_20952 & x_20953;
assign x_52242 = x_52240 & x_52241;
assign x_52243 = x_20954 & x_20955;
assign x_52244 = x_20956 & x_20957;
assign x_52245 = x_52243 & x_52244;
assign x_52246 = x_52242 & x_52245;
assign x_52247 = x_20958 & x_20959;
assign x_52248 = x_20960 & x_20961;
assign x_52249 = x_52247 & x_52248;
assign x_52250 = x_20962 & x_20963;
assign x_52251 = x_20964 & x_20965;
assign x_52252 = x_52250 & x_52251;
assign x_52253 = x_52249 & x_52252;
assign x_52254 = x_52246 & x_52253;
assign x_52255 = x_52239 & x_52254;
assign x_52256 = x_52225 & x_52255;
assign x_52257 = x_20967 & x_20968;
assign x_52258 = x_20966 & x_52257;
assign x_52259 = x_20969 & x_20970;
assign x_52260 = x_20971 & x_20972;
assign x_52261 = x_52259 & x_52260;
assign x_52262 = x_52258 & x_52261;
assign x_52263 = x_20973 & x_20974;
assign x_52264 = x_20975 & x_20976;
assign x_52265 = x_52263 & x_52264;
assign x_52266 = x_20977 & x_20978;
assign x_52267 = x_20979 & x_20980;
assign x_52268 = x_52266 & x_52267;
assign x_52269 = x_52265 & x_52268;
assign x_52270 = x_52262 & x_52269;
assign x_52271 = x_20981 & x_20982;
assign x_52272 = x_20983 & x_20984;
assign x_52273 = x_52271 & x_52272;
assign x_52274 = x_20985 & x_20986;
assign x_52275 = x_20987 & x_20988;
assign x_52276 = x_52274 & x_52275;
assign x_52277 = x_52273 & x_52276;
assign x_52278 = x_20989 & x_20990;
assign x_52279 = x_20991 & x_20992;
assign x_52280 = x_52278 & x_52279;
assign x_52281 = x_20993 & x_20994;
assign x_52282 = x_20995 & x_20996;
assign x_52283 = x_52281 & x_52282;
assign x_52284 = x_52280 & x_52283;
assign x_52285 = x_52277 & x_52284;
assign x_52286 = x_52270 & x_52285;
assign x_52287 = x_20998 & x_20999;
assign x_52288 = x_20997 & x_52287;
assign x_52289 = x_21000 & x_21001;
assign x_52290 = x_21002 & x_21003;
assign x_52291 = x_52289 & x_52290;
assign x_52292 = x_52288 & x_52291;
assign x_52293 = x_21004 & x_21005;
assign x_52294 = x_21006 & x_21007;
assign x_52295 = x_52293 & x_52294;
assign x_52296 = x_21008 & x_21009;
assign x_52297 = x_21010 & x_21011;
assign x_52298 = x_52296 & x_52297;
assign x_52299 = x_52295 & x_52298;
assign x_52300 = x_52292 & x_52299;
assign x_52301 = x_21012 & x_21013;
assign x_52302 = x_21014 & x_21015;
assign x_52303 = x_52301 & x_52302;
assign x_52304 = x_21016 & x_21017;
assign x_52305 = x_21018 & x_21019;
assign x_52306 = x_52304 & x_52305;
assign x_52307 = x_52303 & x_52306;
assign x_52308 = x_21020 & x_21021;
assign x_52309 = x_21022 & x_21023;
assign x_52310 = x_52308 & x_52309;
assign x_52311 = x_21024 & x_21025;
assign x_52312 = x_21026 & x_21027;
assign x_52313 = x_52311 & x_52312;
assign x_52314 = x_52310 & x_52313;
assign x_52315 = x_52307 & x_52314;
assign x_52316 = x_52300 & x_52315;
assign x_52317 = x_52286 & x_52316;
assign x_52318 = x_52256 & x_52317;
assign x_52319 = x_52196 & x_52318;
assign x_52320 = x_52075 & x_52319;
assign x_52321 = x_21029 & x_21030;
assign x_52322 = x_21028 & x_52321;
assign x_52323 = x_21031 & x_21032;
assign x_52324 = x_21033 & x_21034;
assign x_52325 = x_52323 & x_52324;
assign x_52326 = x_52322 & x_52325;
assign x_52327 = x_21035 & x_21036;
assign x_52328 = x_21037 & x_21038;
assign x_52329 = x_52327 & x_52328;
assign x_52330 = x_21039 & x_21040;
assign x_52331 = x_21041 & x_21042;
assign x_52332 = x_52330 & x_52331;
assign x_52333 = x_52329 & x_52332;
assign x_52334 = x_52326 & x_52333;
assign x_52335 = x_21044 & x_21045;
assign x_52336 = x_21043 & x_52335;
assign x_52337 = x_21046 & x_21047;
assign x_52338 = x_21048 & x_21049;
assign x_52339 = x_52337 & x_52338;
assign x_52340 = x_52336 & x_52339;
assign x_52341 = x_21050 & x_21051;
assign x_52342 = x_21052 & x_21053;
assign x_52343 = x_52341 & x_52342;
assign x_52344 = x_21054 & x_21055;
assign x_52345 = x_21056 & x_21057;
assign x_52346 = x_52344 & x_52345;
assign x_52347 = x_52343 & x_52346;
assign x_52348 = x_52340 & x_52347;
assign x_52349 = x_52334 & x_52348;
assign x_52350 = x_21059 & x_21060;
assign x_52351 = x_21058 & x_52350;
assign x_52352 = x_21061 & x_21062;
assign x_52353 = x_21063 & x_21064;
assign x_52354 = x_52352 & x_52353;
assign x_52355 = x_52351 & x_52354;
assign x_52356 = x_21065 & x_21066;
assign x_52357 = x_21067 & x_21068;
assign x_52358 = x_52356 & x_52357;
assign x_52359 = x_21069 & x_21070;
assign x_52360 = x_21071 & x_21072;
assign x_52361 = x_52359 & x_52360;
assign x_52362 = x_52358 & x_52361;
assign x_52363 = x_52355 & x_52362;
assign x_52364 = x_21073 & x_21074;
assign x_52365 = x_21075 & x_21076;
assign x_52366 = x_52364 & x_52365;
assign x_52367 = x_21077 & x_21078;
assign x_52368 = x_21079 & x_21080;
assign x_52369 = x_52367 & x_52368;
assign x_52370 = x_52366 & x_52369;
assign x_52371 = x_21081 & x_21082;
assign x_52372 = x_21083 & x_21084;
assign x_52373 = x_52371 & x_52372;
assign x_52374 = x_21085 & x_21086;
assign x_52375 = x_21087 & x_21088;
assign x_52376 = x_52374 & x_52375;
assign x_52377 = x_52373 & x_52376;
assign x_52378 = x_52370 & x_52377;
assign x_52379 = x_52363 & x_52378;
assign x_52380 = x_52349 & x_52379;
assign x_52381 = x_21090 & x_21091;
assign x_52382 = x_21089 & x_52381;
assign x_52383 = x_21092 & x_21093;
assign x_52384 = x_21094 & x_21095;
assign x_52385 = x_52383 & x_52384;
assign x_52386 = x_52382 & x_52385;
assign x_52387 = x_21096 & x_21097;
assign x_52388 = x_21098 & x_21099;
assign x_52389 = x_52387 & x_52388;
assign x_52390 = x_21100 & x_21101;
assign x_52391 = x_21102 & x_21103;
assign x_52392 = x_52390 & x_52391;
assign x_52393 = x_52389 & x_52392;
assign x_52394 = x_52386 & x_52393;
assign x_52395 = x_21105 & x_21106;
assign x_52396 = x_21104 & x_52395;
assign x_52397 = x_21107 & x_21108;
assign x_52398 = x_21109 & x_21110;
assign x_52399 = x_52397 & x_52398;
assign x_52400 = x_52396 & x_52399;
assign x_52401 = x_21111 & x_21112;
assign x_52402 = x_21113 & x_21114;
assign x_52403 = x_52401 & x_52402;
assign x_52404 = x_21115 & x_21116;
assign x_52405 = x_21117 & x_21118;
assign x_52406 = x_52404 & x_52405;
assign x_52407 = x_52403 & x_52406;
assign x_52408 = x_52400 & x_52407;
assign x_52409 = x_52394 & x_52408;
assign x_52410 = x_21120 & x_21121;
assign x_52411 = x_21119 & x_52410;
assign x_52412 = x_21122 & x_21123;
assign x_52413 = x_21124 & x_21125;
assign x_52414 = x_52412 & x_52413;
assign x_52415 = x_52411 & x_52414;
assign x_52416 = x_21126 & x_21127;
assign x_52417 = x_21128 & x_21129;
assign x_52418 = x_52416 & x_52417;
assign x_52419 = x_21130 & x_21131;
assign x_52420 = x_21132 & x_21133;
assign x_52421 = x_52419 & x_52420;
assign x_52422 = x_52418 & x_52421;
assign x_52423 = x_52415 & x_52422;
assign x_52424 = x_21134 & x_21135;
assign x_52425 = x_21136 & x_21137;
assign x_52426 = x_52424 & x_52425;
assign x_52427 = x_21138 & x_21139;
assign x_52428 = x_21140 & x_21141;
assign x_52429 = x_52427 & x_52428;
assign x_52430 = x_52426 & x_52429;
assign x_52431 = x_21142 & x_21143;
assign x_52432 = x_21144 & x_21145;
assign x_52433 = x_52431 & x_52432;
assign x_52434 = x_21146 & x_21147;
assign x_52435 = x_21148 & x_21149;
assign x_52436 = x_52434 & x_52435;
assign x_52437 = x_52433 & x_52436;
assign x_52438 = x_52430 & x_52437;
assign x_52439 = x_52423 & x_52438;
assign x_52440 = x_52409 & x_52439;
assign x_52441 = x_52380 & x_52440;
assign x_52442 = x_21151 & x_21152;
assign x_52443 = x_21150 & x_52442;
assign x_52444 = x_21153 & x_21154;
assign x_52445 = x_21155 & x_21156;
assign x_52446 = x_52444 & x_52445;
assign x_52447 = x_52443 & x_52446;
assign x_52448 = x_21157 & x_21158;
assign x_52449 = x_21159 & x_21160;
assign x_52450 = x_52448 & x_52449;
assign x_52451 = x_21161 & x_21162;
assign x_52452 = x_21163 & x_21164;
assign x_52453 = x_52451 & x_52452;
assign x_52454 = x_52450 & x_52453;
assign x_52455 = x_52447 & x_52454;
assign x_52456 = x_21166 & x_21167;
assign x_52457 = x_21165 & x_52456;
assign x_52458 = x_21168 & x_21169;
assign x_52459 = x_21170 & x_21171;
assign x_52460 = x_52458 & x_52459;
assign x_52461 = x_52457 & x_52460;
assign x_52462 = x_21172 & x_21173;
assign x_52463 = x_21174 & x_21175;
assign x_52464 = x_52462 & x_52463;
assign x_52465 = x_21176 & x_21177;
assign x_52466 = x_21178 & x_21179;
assign x_52467 = x_52465 & x_52466;
assign x_52468 = x_52464 & x_52467;
assign x_52469 = x_52461 & x_52468;
assign x_52470 = x_52455 & x_52469;
assign x_52471 = x_21181 & x_21182;
assign x_52472 = x_21180 & x_52471;
assign x_52473 = x_21183 & x_21184;
assign x_52474 = x_21185 & x_21186;
assign x_52475 = x_52473 & x_52474;
assign x_52476 = x_52472 & x_52475;
assign x_52477 = x_21187 & x_21188;
assign x_52478 = x_21189 & x_21190;
assign x_52479 = x_52477 & x_52478;
assign x_52480 = x_21191 & x_21192;
assign x_52481 = x_21193 & x_21194;
assign x_52482 = x_52480 & x_52481;
assign x_52483 = x_52479 & x_52482;
assign x_52484 = x_52476 & x_52483;
assign x_52485 = x_21195 & x_21196;
assign x_52486 = x_21197 & x_21198;
assign x_52487 = x_52485 & x_52486;
assign x_52488 = x_21199 & x_21200;
assign x_52489 = x_21201 & x_21202;
assign x_52490 = x_52488 & x_52489;
assign x_52491 = x_52487 & x_52490;
assign x_52492 = x_21203 & x_21204;
assign x_52493 = x_21205 & x_21206;
assign x_52494 = x_52492 & x_52493;
assign x_52495 = x_21207 & x_21208;
assign x_52496 = x_21209 & x_21210;
assign x_52497 = x_52495 & x_52496;
assign x_52498 = x_52494 & x_52497;
assign x_52499 = x_52491 & x_52498;
assign x_52500 = x_52484 & x_52499;
assign x_52501 = x_52470 & x_52500;
assign x_52502 = x_21212 & x_21213;
assign x_52503 = x_21211 & x_52502;
assign x_52504 = x_21214 & x_21215;
assign x_52505 = x_21216 & x_21217;
assign x_52506 = x_52504 & x_52505;
assign x_52507 = x_52503 & x_52506;
assign x_52508 = x_21218 & x_21219;
assign x_52509 = x_21220 & x_21221;
assign x_52510 = x_52508 & x_52509;
assign x_52511 = x_21222 & x_21223;
assign x_52512 = x_21224 & x_21225;
assign x_52513 = x_52511 & x_52512;
assign x_52514 = x_52510 & x_52513;
assign x_52515 = x_52507 & x_52514;
assign x_52516 = x_21227 & x_21228;
assign x_52517 = x_21226 & x_52516;
assign x_52518 = x_21229 & x_21230;
assign x_52519 = x_21231 & x_21232;
assign x_52520 = x_52518 & x_52519;
assign x_52521 = x_52517 & x_52520;
assign x_52522 = x_21233 & x_21234;
assign x_52523 = x_21235 & x_21236;
assign x_52524 = x_52522 & x_52523;
assign x_52525 = x_21237 & x_21238;
assign x_52526 = x_21239 & x_21240;
assign x_52527 = x_52525 & x_52526;
assign x_52528 = x_52524 & x_52527;
assign x_52529 = x_52521 & x_52528;
assign x_52530 = x_52515 & x_52529;
assign x_52531 = x_21242 & x_21243;
assign x_52532 = x_21241 & x_52531;
assign x_52533 = x_21244 & x_21245;
assign x_52534 = x_21246 & x_21247;
assign x_52535 = x_52533 & x_52534;
assign x_52536 = x_52532 & x_52535;
assign x_52537 = x_21248 & x_21249;
assign x_52538 = x_21250 & x_21251;
assign x_52539 = x_52537 & x_52538;
assign x_52540 = x_21252 & x_21253;
assign x_52541 = x_21254 & x_21255;
assign x_52542 = x_52540 & x_52541;
assign x_52543 = x_52539 & x_52542;
assign x_52544 = x_52536 & x_52543;
assign x_52545 = x_21256 & x_21257;
assign x_52546 = x_21258 & x_21259;
assign x_52547 = x_52545 & x_52546;
assign x_52548 = x_21260 & x_21261;
assign x_52549 = x_21262 & x_21263;
assign x_52550 = x_52548 & x_52549;
assign x_52551 = x_52547 & x_52550;
assign x_52552 = x_21264 & x_21265;
assign x_52553 = x_21266 & x_21267;
assign x_52554 = x_52552 & x_52553;
assign x_52555 = x_21268 & x_21269;
assign x_52556 = x_21270 & x_21271;
assign x_52557 = x_52555 & x_52556;
assign x_52558 = x_52554 & x_52557;
assign x_52559 = x_52551 & x_52558;
assign x_52560 = x_52544 & x_52559;
assign x_52561 = x_52530 & x_52560;
assign x_52562 = x_52501 & x_52561;
assign x_52563 = x_52441 & x_52562;
assign x_52564 = x_21273 & x_21274;
assign x_52565 = x_21272 & x_52564;
assign x_52566 = x_21275 & x_21276;
assign x_52567 = x_21277 & x_21278;
assign x_52568 = x_52566 & x_52567;
assign x_52569 = x_52565 & x_52568;
assign x_52570 = x_21279 & x_21280;
assign x_52571 = x_21281 & x_21282;
assign x_52572 = x_52570 & x_52571;
assign x_52573 = x_21283 & x_21284;
assign x_52574 = x_21285 & x_21286;
assign x_52575 = x_52573 & x_52574;
assign x_52576 = x_52572 & x_52575;
assign x_52577 = x_52569 & x_52576;
assign x_52578 = x_21288 & x_21289;
assign x_52579 = x_21287 & x_52578;
assign x_52580 = x_21290 & x_21291;
assign x_52581 = x_21292 & x_21293;
assign x_52582 = x_52580 & x_52581;
assign x_52583 = x_52579 & x_52582;
assign x_52584 = x_21294 & x_21295;
assign x_52585 = x_21296 & x_21297;
assign x_52586 = x_52584 & x_52585;
assign x_52587 = x_21298 & x_21299;
assign x_52588 = x_21300 & x_21301;
assign x_52589 = x_52587 & x_52588;
assign x_52590 = x_52586 & x_52589;
assign x_52591 = x_52583 & x_52590;
assign x_52592 = x_52577 & x_52591;
assign x_52593 = x_21303 & x_21304;
assign x_52594 = x_21302 & x_52593;
assign x_52595 = x_21305 & x_21306;
assign x_52596 = x_21307 & x_21308;
assign x_52597 = x_52595 & x_52596;
assign x_52598 = x_52594 & x_52597;
assign x_52599 = x_21309 & x_21310;
assign x_52600 = x_21311 & x_21312;
assign x_52601 = x_52599 & x_52600;
assign x_52602 = x_21313 & x_21314;
assign x_52603 = x_21315 & x_21316;
assign x_52604 = x_52602 & x_52603;
assign x_52605 = x_52601 & x_52604;
assign x_52606 = x_52598 & x_52605;
assign x_52607 = x_21317 & x_21318;
assign x_52608 = x_21319 & x_21320;
assign x_52609 = x_52607 & x_52608;
assign x_52610 = x_21321 & x_21322;
assign x_52611 = x_21323 & x_21324;
assign x_52612 = x_52610 & x_52611;
assign x_52613 = x_52609 & x_52612;
assign x_52614 = x_21325 & x_21326;
assign x_52615 = x_21327 & x_21328;
assign x_52616 = x_52614 & x_52615;
assign x_52617 = x_21329 & x_21330;
assign x_52618 = x_21331 & x_21332;
assign x_52619 = x_52617 & x_52618;
assign x_52620 = x_52616 & x_52619;
assign x_52621 = x_52613 & x_52620;
assign x_52622 = x_52606 & x_52621;
assign x_52623 = x_52592 & x_52622;
assign x_52624 = x_21334 & x_21335;
assign x_52625 = x_21333 & x_52624;
assign x_52626 = x_21336 & x_21337;
assign x_52627 = x_21338 & x_21339;
assign x_52628 = x_52626 & x_52627;
assign x_52629 = x_52625 & x_52628;
assign x_52630 = x_21340 & x_21341;
assign x_52631 = x_21342 & x_21343;
assign x_52632 = x_52630 & x_52631;
assign x_52633 = x_21344 & x_21345;
assign x_52634 = x_21346 & x_21347;
assign x_52635 = x_52633 & x_52634;
assign x_52636 = x_52632 & x_52635;
assign x_52637 = x_52629 & x_52636;
assign x_52638 = x_21349 & x_21350;
assign x_52639 = x_21348 & x_52638;
assign x_52640 = x_21351 & x_21352;
assign x_52641 = x_21353 & x_21354;
assign x_52642 = x_52640 & x_52641;
assign x_52643 = x_52639 & x_52642;
assign x_52644 = x_21355 & x_21356;
assign x_52645 = x_21357 & x_21358;
assign x_52646 = x_52644 & x_52645;
assign x_52647 = x_21359 & x_21360;
assign x_52648 = x_21361 & x_21362;
assign x_52649 = x_52647 & x_52648;
assign x_52650 = x_52646 & x_52649;
assign x_52651 = x_52643 & x_52650;
assign x_52652 = x_52637 & x_52651;
assign x_52653 = x_21364 & x_21365;
assign x_52654 = x_21363 & x_52653;
assign x_52655 = x_21366 & x_21367;
assign x_52656 = x_21368 & x_21369;
assign x_52657 = x_52655 & x_52656;
assign x_52658 = x_52654 & x_52657;
assign x_52659 = x_21370 & x_21371;
assign x_52660 = x_21372 & x_21373;
assign x_52661 = x_52659 & x_52660;
assign x_52662 = x_21374 & x_21375;
assign x_52663 = x_21376 & x_21377;
assign x_52664 = x_52662 & x_52663;
assign x_52665 = x_52661 & x_52664;
assign x_52666 = x_52658 & x_52665;
assign x_52667 = x_21378 & x_21379;
assign x_52668 = x_21380 & x_21381;
assign x_52669 = x_52667 & x_52668;
assign x_52670 = x_21382 & x_21383;
assign x_52671 = x_21384 & x_21385;
assign x_52672 = x_52670 & x_52671;
assign x_52673 = x_52669 & x_52672;
assign x_52674 = x_21386 & x_21387;
assign x_52675 = x_21388 & x_21389;
assign x_52676 = x_52674 & x_52675;
assign x_52677 = x_21390 & x_21391;
assign x_52678 = x_21392 & x_21393;
assign x_52679 = x_52677 & x_52678;
assign x_52680 = x_52676 & x_52679;
assign x_52681 = x_52673 & x_52680;
assign x_52682 = x_52666 & x_52681;
assign x_52683 = x_52652 & x_52682;
assign x_52684 = x_52623 & x_52683;
assign x_52685 = x_21395 & x_21396;
assign x_52686 = x_21394 & x_52685;
assign x_52687 = x_21397 & x_21398;
assign x_52688 = x_21399 & x_21400;
assign x_52689 = x_52687 & x_52688;
assign x_52690 = x_52686 & x_52689;
assign x_52691 = x_21401 & x_21402;
assign x_52692 = x_21403 & x_21404;
assign x_52693 = x_52691 & x_52692;
assign x_52694 = x_21405 & x_21406;
assign x_52695 = x_21407 & x_21408;
assign x_52696 = x_52694 & x_52695;
assign x_52697 = x_52693 & x_52696;
assign x_52698 = x_52690 & x_52697;
assign x_52699 = x_21410 & x_21411;
assign x_52700 = x_21409 & x_52699;
assign x_52701 = x_21412 & x_21413;
assign x_52702 = x_21414 & x_21415;
assign x_52703 = x_52701 & x_52702;
assign x_52704 = x_52700 & x_52703;
assign x_52705 = x_21416 & x_21417;
assign x_52706 = x_21418 & x_21419;
assign x_52707 = x_52705 & x_52706;
assign x_52708 = x_21420 & x_21421;
assign x_52709 = x_21422 & x_21423;
assign x_52710 = x_52708 & x_52709;
assign x_52711 = x_52707 & x_52710;
assign x_52712 = x_52704 & x_52711;
assign x_52713 = x_52698 & x_52712;
assign x_52714 = x_21425 & x_21426;
assign x_52715 = x_21424 & x_52714;
assign x_52716 = x_21427 & x_21428;
assign x_52717 = x_21429 & x_21430;
assign x_52718 = x_52716 & x_52717;
assign x_52719 = x_52715 & x_52718;
assign x_52720 = x_21431 & x_21432;
assign x_52721 = x_21433 & x_21434;
assign x_52722 = x_52720 & x_52721;
assign x_52723 = x_21435 & x_21436;
assign x_52724 = x_21437 & x_21438;
assign x_52725 = x_52723 & x_52724;
assign x_52726 = x_52722 & x_52725;
assign x_52727 = x_52719 & x_52726;
assign x_52728 = x_21439 & x_21440;
assign x_52729 = x_21441 & x_21442;
assign x_52730 = x_52728 & x_52729;
assign x_52731 = x_21443 & x_21444;
assign x_52732 = x_21445 & x_21446;
assign x_52733 = x_52731 & x_52732;
assign x_52734 = x_52730 & x_52733;
assign x_52735 = x_21447 & x_21448;
assign x_52736 = x_21449 & x_21450;
assign x_52737 = x_52735 & x_52736;
assign x_52738 = x_21451 & x_21452;
assign x_52739 = x_21453 & x_21454;
assign x_52740 = x_52738 & x_52739;
assign x_52741 = x_52737 & x_52740;
assign x_52742 = x_52734 & x_52741;
assign x_52743 = x_52727 & x_52742;
assign x_52744 = x_52713 & x_52743;
assign x_52745 = x_21456 & x_21457;
assign x_52746 = x_21455 & x_52745;
assign x_52747 = x_21458 & x_21459;
assign x_52748 = x_21460 & x_21461;
assign x_52749 = x_52747 & x_52748;
assign x_52750 = x_52746 & x_52749;
assign x_52751 = x_21462 & x_21463;
assign x_52752 = x_21464 & x_21465;
assign x_52753 = x_52751 & x_52752;
assign x_52754 = x_21466 & x_21467;
assign x_52755 = x_21468 & x_21469;
assign x_52756 = x_52754 & x_52755;
assign x_52757 = x_52753 & x_52756;
assign x_52758 = x_52750 & x_52757;
assign x_52759 = x_21470 & x_21471;
assign x_52760 = x_21472 & x_21473;
assign x_52761 = x_52759 & x_52760;
assign x_52762 = x_21474 & x_21475;
assign x_52763 = x_21476 & x_21477;
assign x_52764 = x_52762 & x_52763;
assign x_52765 = x_52761 & x_52764;
assign x_52766 = x_21478 & x_21479;
assign x_52767 = x_21480 & x_21481;
assign x_52768 = x_52766 & x_52767;
assign x_52769 = x_21482 & x_21483;
assign x_52770 = x_21484 & x_21485;
assign x_52771 = x_52769 & x_52770;
assign x_52772 = x_52768 & x_52771;
assign x_52773 = x_52765 & x_52772;
assign x_52774 = x_52758 & x_52773;
assign x_52775 = x_21487 & x_21488;
assign x_52776 = x_21486 & x_52775;
assign x_52777 = x_21489 & x_21490;
assign x_52778 = x_21491 & x_21492;
assign x_52779 = x_52777 & x_52778;
assign x_52780 = x_52776 & x_52779;
assign x_52781 = x_21493 & x_21494;
assign x_52782 = x_21495 & x_21496;
assign x_52783 = x_52781 & x_52782;
assign x_52784 = x_21497 & x_21498;
assign x_52785 = x_21499 & x_21500;
assign x_52786 = x_52784 & x_52785;
assign x_52787 = x_52783 & x_52786;
assign x_52788 = x_52780 & x_52787;
assign x_52789 = x_21501 & x_21502;
assign x_52790 = x_21503 & x_21504;
assign x_52791 = x_52789 & x_52790;
assign x_52792 = x_21505 & x_21506;
assign x_52793 = x_21507 & x_21508;
assign x_52794 = x_52792 & x_52793;
assign x_52795 = x_52791 & x_52794;
assign x_52796 = x_21509 & x_21510;
assign x_52797 = x_21511 & x_21512;
assign x_52798 = x_52796 & x_52797;
assign x_52799 = x_21513 & x_21514;
assign x_52800 = x_21515 & x_21516;
assign x_52801 = x_52799 & x_52800;
assign x_52802 = x_52798 & x_52801;
assign x_52803 = x_52795 & x_52802;
assign x_52804 = x_52788 & x_52803;
assign x_52805 = x_52774 & x_52804;
assign x_52806 = x_52744 & x_52805;
assign x_52807 = x_52684 & x_52806;
assign x_52808 = x_52563 & x_52807;
assign x_52809 = x_52320 & x_52808;
assign x_52810 = x_51832 & x_52809;
assign x_52811 = x_21518 & x_21519;
assign x_52812 = x_21517 & x_52811;
assign x_52813 = x_21520 & x_21521;
assign x_52814 = x_21522 & x_21523;
assign x_52815 = x_52813 & x_52814;
assign x_52816 = x_52812 & x_52815;
assign x_52817 = x_21524 & x_21525;
assign x_52818 = x_21526 & x_21527;
assign x_52819 = x_52817 & x_52818;
assign x_52820 = x_21528 & x_21529;
assign x_52821 = x_21530 & x_21531;
assign x_52822 = x_52820 & x_52821;
assign x_52823 = x_52819 & x_52822;
assign x_52824 = x_52816 & x_52823;
assign x_52825 = x_21533 & x_21534;
assign x_52826 = x_21532 & x_52825;
assign x_52827 = x_21535 & x_21536;
assign x_52828 = x_21537 & x_21538;
assign x_52829 = x_52827 & x_52828;
assign x_52830 = x_52826 & x_52829;
assign x_52831 = x_21539 & x_21540;
assign x_52832 = x_21541 & x_21542;
assign x_52833 = x_52831 & x_52832;
assign x_52834 = x_21543 & x_21544;
assign x_52835 = x_21545 & x_21546;
assign x_52836 = x_52834 & x_52835;
assign x_52837 = x_52833 & x_52836;
assign x_52838 = x_52830 & x_52837;
assign x_52839 = x_52824 & x_52838;
assign x_52840 = x_21548 & x_21549;
assign x_52841 = x_21547 & x_52840;
assign x_52842 = x_21550 & x_21551;
assign x_52843 = x_21552 & x_21553;
assign x_52844 = x_52842 & x_52843;
assign x_52845 = x_52841 & x_52844;
assign x_52846 = x_21554 & x_21555;
assign x_52847 = x_21556 & x_21557;
assign x_52848 = x_52846 & x_52847;
assign x_52849 = x_21558 & x_21559;
assign x_52850 = x_21560 & x_21561;
assign x_52851 = x_52849 & x_52850;
assign x_52852 = x_52848 & x_52851;
assign x_52853 = x_52845 & x_52852;
assign x_52854 = x_21562 & x_21563;
assign x_52855 = x_21564 & x_21565;
assign x_52856 = x_52854 & x_52855;
assign x_52857 = x_21566 & x_21567;
assign x_52858 = x_21568 & x_21569;
assign x_52859 = x_52857 & x_52858;
assign x_52860 = x_52856 & x_52859;
assign x_52861 = x_21570 & x_21571;
assign x_52862 = x_21572 & x_21573;
assign x_52863 = x_52861 & x_52862;
assign x_52864 = x_21574 & x_21575;
assign x_52865 = x_21576 & x_21577;
assign x_52866 = x_52864 & x_52865;
assign x_52867 = x_52863 & x_52866;
assign x_52868 = x_52860 & x_52867;
assign x_52869 = x_52853 & x_52868;
assign x_52870 = x_52839 & x_52869;
assign x_52871 = x_21579 & x_21580;
assign x_52872 = x_21578 & x_52871;
assign x_52873 = x_21581 & x_21582;
assign x_52874 = x_21583 & x_21584;
assign x_52875 = x_52873 & x_52874;
assign x_52876 = x_52872 & x_52875;
assign x_52877 = x_21585 & x_21586;
assign x_52878 = x_21587 & x_21588;
assign x_52879 = x_52877 & x_52878;
assign x_52880 = x_21589 & x_21590;
assign x_52881 = x_21591 & x_21592;
assign x_52882 = x_52880 & x_52881;
assign x_52883 = x_52879 & x_52882;
assign x_52884 = x_52876 & x_52883;
assign x_52885 = x_21594 & x_21595;
assign x_52886 = x_21593 & x_52885;
assign x_52887 = x_21596 & x_21597;
assign x_52888 = x_21598 & x_21599;
assign x_52889 = x_52887 & x_52888;
assign x_52890 = x_52886 & x_52889;
assign x_52891 = x_21600 & x_21601;
assign x_52892 = x_21602 & x_21603;
assign x_52893 = x_52891 & x_52892;
assign x_52894 = x_21604 & x_21605;
assign x_52895 = x_21606 & x_21607;
assign x_52896 = x_52894 & x_52895;
assign x_52897 = x_52893 & x_52896;
assign x_52898 = x_52890 & x_52897;
assign x_52899 = x_52884 & x_52898;
assign x_52900 = x_21609 & x_21610;
assign x_52901 = x_21608 & x_52900;
assign x_52902 = x_21611 & x_21612;
assign x_52903 = x_21613 & x_21614;
assign x_52904 = x_52902 & x_52903;
assign x_52905 = x_52901 & x_52904;
assign x_52906 = x_21615 & x_21616;
assign x_52907 = x_21617 & x_21618;
assign x_52908 = x_52906 & x_52907;
assign x_52909 = x_21619 & x_21620;
assign x_52910 = x_21621 & x_21622;
assign x_52911 = x_52909 & x_52910;
assign x_52912 = x_52908 & x_52911;
assign x_52913 = x_52905 & x_52912;
assign x_52914 = x_21623 & x_21624;
assign x_52915 = x_21625 & x_21626;
assign x_52916 = x_52914 & x_52915;
assign x_52917 = x_21627 & x_21628;
assign x_52918 = x_21629 & x_21630;
assign x_52919 = x_52917 & x_52918;
assign x_52920 = x_52916 & x_52919;
assign x_52921 = x_21631 & x_21632;
assign x_52922 = x_21633 & x_21634;
assign x_52923 = x_52921 & x_52922;
assign x_52924 = x_21635 & x_21636;
assign x_52925 = x_21637 & x_21638;
assign x_52926 = x_52924 & x_52925;
assign x_52927 = x_52923 & x_52926;
assign x_52928 = x_52920 & x_52927;
assign x_52929 = x_52913 & x_52928;
assign x_52930 = x_52899 & x_52929;
assign x_52931 = x_52870 & x_52930;
assign x_52932 = x_21640 & x_21641;
assign x_52933 = x_21639 & x_52932;
assign x_52934 = x_21642 & x_21643;
assign x_52935 = x_21644 & x_21645;
assign x_52936 = x_52934 & x_52935;
assign x_52937 = x_52933 & x_52936;
assign x_52938 = x_21646 & x_21647;
assign x_52939 = x_21648 & x_21649;
assign x_52940 = x_52938 & x_52939;
assign x_52941 = x_21650 & x_21651;
assign x_52942 = x_21652 & x_21653;
assign x_52943 = x_52941 & x_52942;
assign x_52944 = x_52940 & x_52943;
assign x_52945 = x_52937 & x_52944;
assign x_52946 = x_21655 & x_21656;
assign x_52947 = x_21654 & x_52946;
assign x_52948 = x_21657 & x_21658;
assign x_52949 = x_21659 & x_21660;
assign x_52950 = x_52948 & x_52949;
assign x_52951 = x_52947 & x_52950;
assign x_52952 = x_21661 & x_21662;
assign x_52953 = x_21663 & x_21664;
assign x_52954 = x_52952 & x_52953;
assign x_52955 = x_21665 & x_21666;
assign x_52956 = x_21667 & x_21668;
assign x_52957 = x_52955 & x_52956;
assign x_52958 = x_52954 & x_52957;
assign x_52959 = x_52951 & x_52958;
assign x_52960 = x_52945 & x_52959;
assign x_52961 = x_21670 & x_21671;
assign x_52962 = x_21669 & x_52961;
assign x_52963 = x_21672 & x_21673;
assign x_52964 = x_21674 & x_21675;
assign x_52965 = x_52963 & x_52964;
assign x_52966 = x_52962 & x_52965;
assign x_52967 = x_21676 & x_21677;
assign x_52968 = x_21678 & x_21679;
assign x_52969 = x_52967 & x_52968;
assign x_52970 = x_21680 & x_21681;
assign x_52971 = x_21682 & x_21683;
assign x_52972 = x_52970 & x_52971;
assign x_52973 = x_52969 & x_52972;
assign x_52974 = x_52966 & x_52973;
assign x_52975 = x_21684 & x_21685;
assign x_52976 = x_21686 & x_21687;
assign x_52977 = x_52975 & x_52976;
assign x_52978 = x_21688 & x_21689;
assign x_52979 = x_21690 & x_21691;
assign x_52980 = x_52978 & x_52979;
assign x_52981 = x_52977 & x_52980;
assign x_52982 = x_21692 & x_21693;
assign x_52983 = x_21694 & x_21695;
assign x_52984 = x_52982 & x_52983;
assign x_52985 = x_21696 & x_21697;
assign x_52986 = x_21698 & x_21699;
assign x_52987 = x_52985 & x_52986;
assign x_52988 = x_52984 & x_52987;
assign x_52989 = x_52981 & x_52988;
assign x_52990 = x_52974 & x_52989;
assign x_52991 = x_52960 & x_52990;
assign x_52992 = x_21701 & x_21702;
assign x_52993 = x_21700 & x_52992;
assign x_52994 = x_21703 & x_21704;
assign x_52995 = x_21705 & x_21706;
assign x_52996 = x_52994 & x_52995;
assign x_52997 = x_52993 & x_52996;
assign x_52998 = x_21707 & x_21708;
assign x_52999 = x_21709 & x_21710;
assign x_53000 = x_52998 & x_52999;
assign x_53001 = x_21711 & x_21712;
assign x_53002 = x_21713 & x_21714;
assign x_53003 = x_53001 & x_53002;
assign x_53004 = x_53000 & x_53003;
assign x_53005 = x_52997 & x_53004;
assign x_53006 = x_21716 & x_21717;
assign x_53007 = x_21715 & x_53006;
assign x_53008 = x_21718 & x_21719;
assign x_53009 = x_21720 & x_21721;
assign x_53010 = x_53008 & x_53009;
assign x_53011 = x_53007 & x_53010;
assign x_53012 = x_21722 & x_21723;
assign x_53013 = x_21724 & x_21725;
assign x_53014 = x_53012 & x_53013;
assign x_53015 = x_21726 & x_21727;
assign x_53016 = x_21728 & x_21729;
assign x_53017 = x_53015 & x_53016;
assign x_53018 = x_53014 & x_53017;
assign x_53019 = x_53011 & x_53018;
assign x_53020 = x_53005 & x_53019;
assign x_53021 = x_21731 & x_21732;
assign x_53022 = x_21730 & x_53021;
assign x_53023 = x_21733 & x_21734;
assign x_53024 = x_21735 & x_21736;
assign x_53025 = x_53023 & x_53024;
assign x_53026 = x_53022 & x_53025;
assign x_53027 = x_21737 & x_21738;
assign x_53028 = x_21739 & x_21740;
assign x_53029 = x_53027 & x_53028;
assign x_53030 = x_21741 & x_21742;
assign x_53031 = x_21743 & x_21744;
assign x_53032 = x_53030 & x_53031;
assign x_53033 = x_53029 & x_53032;
assign x_53034 = x_53026 & x_53033;
assign x_53035 = x_21745 & x_21746;
assign x_53036 = x_21747 & x_21748;
assign x_53037 = x_53035 & x_53036;
assign x_53038 = x_21749 & x_21750;
assign x_53039 = x_21751 & x_21752;
assign x_53040 = x_53038 & x_53039;
assign x_53041 = x_53037 & x_53040;
assign x_53042 = x_21753 & x_21754;
assign x_53043 = x_21755 & x_21756;
assign x_53044 = x_53042 & x_53043;
assign x_53045 = x_21757 & x_21758;
assign x_53046 = x_21759 & x_21760;
assign x_53047 = x_53045 & x_53046;
assign x_53048 = x_53044 & x_53047;
assign x_53049 = x_53041 & x_53048;
assign x_53050 = x_53034 & x_53049;
assign x_53051 = x_53020 & x_53050;
assign x_53052 = x_52991 & x_53051;
assign x_53053 = x_52931 & x_53052;
assign x_53054 = x_21762 & x_21763;
assign x_53055 = x_21761 & x_53054;
assign x_53056 = x_21764 & x_21765;
assign x_53057 = x_21766 & x_21767;
assign x_53058 = x_53056 & x_53057;
assign x_53059 = x_53055 & x_53058;
assign x_53060 = x_21768 & x_21769;
assign x_53061 = x_21770 & x_21771;
assign x_53062 = x_53060 & x_53061;
assign x_53063 = x_21772 & x_21773;
assign x_53064 = x_21774 & x_21775;
assign x_53065 = x_53063 & x_53064;
assign x_53066 = x_53062 & x_53065;
assign x_53067 = x_53059 & x_53066;
assign x_53068 = x_21777 & x_21778;
assign x_53069 = x_21776 & x_53068;
assign x_53070 = x_21779 & x_21780;
assign x_53071 = x_21781 & x_21782;
assign x_53072 = x_53070 & x_53071;
assign x_53073 = x_53069 & x_53072;
assign x_53074 = x_21783 & x_21784;
assign x_53075 = x_21785 & x_21786;
assign x_53076 = x_53074 & x_53075;
assign x_53077 = x_21787 & x_21788;
assign x_53078 = x_21789 & x_21790;
assign x_53079 = x_53077 & x_53078;
assign x_53080 = x_53076 & x_53079;
assign x_53081 = x_53073 & x_53080;
assign x_53082 = x_53067 & x_53081;
assign x_53083 = x_21792 & x_21793;
assign x_53084 = x_21791 & x_53083;
assign x_53085 = x_21794 & x_21795;
assign x_53086 = x_21796 & x_21797;
assign x_53087 = x_53085 & x_53086;
assign x_53088 = x_53084 & x_53087;
assign x_53089 = x_21798 & x_21799;
assign x_53090 = x_21800 & x_21801;
assign x_53091 = x_53089 & x_53090;
assign x_53092 = x_21802 & x_21803;
assign x_53093 = x_21804 & x_21805;
assign x_53094 = x_53092 & x_53093;
assign x_53095 = x_53091 & x_53094;
assign x_53096 = x_53088 & x_53095;
assign x_53097 = x_21806 & x_21807;
assign x_53098 = x_21808 & x_21809;
assign x_53099 = x_53097 & x_53098;
assign x_53100 = x_21810 & x_21811;
assign x_53101 = x_21812 & x_21813;
assign x_53102 = x_53100 & x_53101;
assign x_53103 = x_53099 & x_53102;
assign x_53104 = x_21814 & x_21815;
assign x_53105 = x_21816 & x_21817;
assign x_53106 = x_53104 & x_53105;
assign x_53107 = x_21818 & x_21819;
assign x_53108 = x_21820 & x_21821;
assign x_53109 = x_53107 & x_53108;
assign x_53110 = x_53106 & x_53109;
assign x_53111 = x_53103 & x_53110;
assign x_53112 = x_53096 & x_53111;
assign x_53113 = x_53082 & x_53112;
assign x_53114 = x_21823 & x_21824;
assign x_53115 = x_21822 & x_53114;
assign x_53116 = x_21825 & x_21826;
assign x_53117 = x_21827 & x_21828;
assign x_53118 = x_53116 & x_53117;
assign x_53119 = x_53115 & x_53118;
assign x_53120 = x_21829 & x_21830;
assign x_53121 = x_21831 & x_21832;
assign x_53122 = x_53120 & x_53121;
assign x_53123 = x_21833 & x_21834;
assign x_53124 = x_21835 & x_21836;
assign x_53125 = x_53123 & x_53124;
assign x_53126 = x_53122 & x_53125;
assign x_53127 = x_53119 & x_53126;
assign x_53128 = x_21838 & x_21839;
assign x_53129 = x_21837 & x_53128;
assign x_53130 = x_21840 & x_21841;
assign x_53131 = x_21842 & x_21843;
assign x_53132 = x_53130 & x_53131;
assign x_53133 = x_53129 & x_53132;
assign x_53134 = x_21844 & x_21845;
assign x_53135 = x_21846 & x_21847;
assign x_53136 = x_53134 & x_53135;
assign x_53137 = x_21848 & x_21849;
assign x_53138 = x_21850 & x_21851;
assign x_53139 = x_53137 & x_53138;
assign x_53140 = x_53136 & x_53139;
assign x_53141 = x_53133 & x_53140;
assign x_53142 = x_53127 & x_53141;
assign x_53143 = x_21853 & x_21854;
assign x_53144 = x_21852 & x_53143;
assign x_53145 = x_21855 & x_21856;
assign x_53146 = x_21857 & x_21858;
assign x_53147 = x_53145 & x_53146;
assign x_53148 = x_53144 & x_53147;
assign x_53149 = x_21859 & x_21860;
assign x_53150 = x_21861 & x_21862;
assign x_53151 = x_53149 & x_53150;
assign x_53152 = x_21863 & x_21864;
assign x_53153 = x_21865 & x_21866;
assign x_53154 = x_53152 & x_53153;
assign x_53155 = x_53151 & x_53154;
assign x_53156 = x_53148 & x_53155;
assign x_53157 = x_21867 & x_21868;
assign x_53158 = x_21869 & x_21870;
assign x_53159 = x_53157 & x_53158;
assign x_53160 = x_21871 & x_21872;
assign x_53161 = x_21873 & x_21874;
assign x_53162 = x_53160 & x_53161;
assign x_53163 = x_53159 & x_53162;
assign x_53164 = x_21875 & x_21876;
assign x_53165 = x_21877 & x_21878;
assign x_53166 = x_53164 & x_53165;
assign x_53167 = x_21879 & x_21880;
assign x_53168 = x_21881 & x_21882;
assign x_53169 = x_53167 & x_53168;
assign x_53170 = x_53166 & x_53169;
assign x_53171 = x_53163 & x_53170;
assign x_53172 = x_53156 & x_53171;
assign x_53173 = x_53142 & x_53172;
assign x_53174 = x_53113 & x_53173;
assign x_53175 = x_21884 & x_21885;
assign x_53176 = x_21883 & x_53175;
assign x_53177 = x_21886 & x_21887;
assign x_53178 = x_21888 & x_21889;
assign x_53179 = x_53177 & x_53178;
assign x_53180 = x_53176 & x_53179;
assign x_53181 = x_21890 & x_21891;
assign x_53182 = x_21892 & x_21893;
assign x_53183 = x_53181 & x_53182;
assign x_53184 = x_21894 & x_21895;
assign x_53185 = x_21896 & x_21897;
assign x_53186 = x_53184 & x_53185;
assign x_53187 = x_53183 & x_53186;
assign x_53188 = x_53180 & x_53187;
assign x_53189 = x_21899 & x_21900;
assign x_53190 = x_21898 & x_53189;
assign x_53191 = x_21901 & x_21902;
assign x_53192 = x_21903 & x_21904;
assign x_53193 = x_53191 & x_53192;
assign x_53194 = x_53190 & x_53193;
assign x_53195 = x_21905 & x_21906;
assign x_53196 = x_21907 & x_21908;
assign x_53197 = x_53195 & x_53196;
assign x_53198 = x_21909 & x_21910;
assign x_53199 = x_21911 & x_21912;
assign x_53200 = x_53198 & x_53199;
assign x_53201 = x_53197 & x_53200;
assign x_53202 = x_53194 & x_53201;
assign x_53203 = x_53188 & x_53202;
assign x_53204 = x_21914 & x_21915;
assign x_53205 = x_21913 & x_53204;
assign x_53206 = x_21916 & x_21917;
assign x_53207 = x_21918 & x_21919;
assign x_53208 = x_53206 & x_53207;
assign x_53209 = x_53205 & x_53208;
assign x_53210 = x_21920 & x_21921;
assign x_53211 = x_21922 & x_21923;
assign x_53212 = x_53210 & x_53211;
assign x_53213 = x_21924 & x_21925;
assign x_53214 = x_21926 & x_21927;
assign x_53215 = x_53213 & x_53214;
assign x_53216 = x_53212 & x_53215;
assign x_53217 = x_53209 & x_53216;
assign x_53218 = x_21928 & x_21929;
assign x_53219 = x_21930 & x_21931;
assign x_53220 = x_53218 & x_53219;
assign x_53221 = x_21932 & x_21933;
assign x_53222 = x_21934 & x_21935;
assign x_53223 = x_53221 & x_53222;
assign x_53224 = x_53220 & x_53223;
assign x_53225 = x_21936 & x_21937;
assign x_53226 = x_21938 & x_21939;
assign x_53227 = x_53225 & x_53226;
assign x_53228 = x_21940 & x_21941;
assign x_53229 = x_21942 & x_21943;
assign x_53230 = x_53228 & x_53229;
assign x_53231 = x_53227 & x_53230;
assign x_53232 = x_53224 & x_53231;
assign x_53233 = x_53217 & x_53232;
assign x_53234 = x_53203 & x_53233;
assign x_53235 = x_21945 & x_21946;
assign x_53236 = x_21944 & x_53235;
assign x_53237 = x_21947 & x_21948;
assign x_53238 = x_21949 & x_21950;
assign x_53239 = x_53237 & x_53238;
assign x_53240 = x_53236 & x_53239;
assign x_53241 = x_21951 & x_21952;
assign x_53242 = x_21953 & x_21954;
assign x_53243 = x_53241 & x_53242;
assign x_53244 = x_21955 & x_21956;
assign x_53245 = x_21957 & x_21958;
assign x_53246 = x_53244 & x_53245;
assign x_53247 = x_53243 & x_53246;
assign x_53248 = x_53240 & x_53247;
assign x_53249 = x_21959 & x_21960;
assign x_53250 = x_21961 & x_21962;
assign x_53251 = x_53249 & x_53250;
assign x_53252 = x_21963 & x_21964;
assign x_53253 = x_21965 & x_21966;
assign x_53254 = x_53252 & x_53253;
assign x_53255 = x_53251 & x_53254;
assign x_53256 = x_21967 & x_21968;
assign x_53257 = x_21969 & x_21970;
assign x_53258 = x_53256 & x_53257;
assign x_53259 = x_21971 & x_21972;
assign x_53260 = x_21973 & x_21974;
assign x_53261 = x_53259 & x_53260;
assign x_53262 = x_53258 & x_53261;
assign x_53263 = x_53255 & x_53262;
assign x_53264 = x_53248 & x_53263;
assign x_53265 = x_21976 & x_21977;
assign x_53266 = x_21975 & x_53265;
assign x_53267 = x_21978 & x_21979;
assign x_53268 = x_21980 & x_21981;
assign x_53269 = x_53267 & x_53268;
assign x_53270 = x_53266 & x_53269;
assign x_53271 = x_21982 & x_21983;
assign x_53272 = x_21984 & x_21985;
assign x_53273 = x_53271 & x_53272;
assign x_53274 = x_21986 & x_21987;
assign x_53275 = x_21988 & x_21989;
assign x_53276 = x_53274 & x_53275;
assign x_53277 = x_53273 & x_53276;
assign x_53278 = x_53270 & x_53277;
assign x_53279 = x_21990 & x_21991;
assign x_53280 = x_21992 & x_21993;
assign x_53281 = x_53279 & x_53280;
assign x_53282 = x_21994 & x_21995;
assign x_53283 = x_21996 & x_21997;
assign x_53284 = x_53282 & x_53283;
assign x_53285 = x_53281 & x_53284;
assign x_53286 = x_21998 & x_21999;
assign x_53287 = x_22000 & x_22001;
assign x_53288 = x_53286 & x_53287;
assign x_53289 = x_22002 & x_22003;
assign x_53290 = x_22004 & x_22005;
assign x_53291 = x_53289 & x_53290;
assign x_53292 = x_53288 & x_53291;
assign x_53293 = x_53285 & x_53292;
assign x_53294 = x_53278 & x_53293;
assign x_53295 = x_53264 & x_53294;
assign x_53296 = x_53234 & x_53295;
assign x_53297 = x_53174 & x_53296;
assign x_53298 = x_53053 & x_53297;
assign x_53299 = x_22007 & x_22008;
assign x_53300 = x_22006 & x_53299;
assign x_53301 = x_22009 & x_22010;
assign x_53302 = x_22011 & x_22012;
assign x_53303 = x_53301 & x_53302;
assign x_53304 = x_53300 & x_53303;
assign x_53305 = x_22013 & x_22014;
assign x_53306 = x_22015 & x_22016;
assign x_53307 = x_53305 & x_53306;
assign x_53308 = x_22017 & x_22018;
assign x_53309 = x_22019 & x_22020;
assign x_53310 = x_53308 & x_53309;
assign x_53311 = x_53307 & x_53310;
assign x_53312 = x_53304 & x_53311;
assign x_53313 = x_22022 & x_22023;
assign x_53314 = x_22021 & x_53313;
assign x_53315 = x_22024 & x_22025;
assign x_53316 = x_22026 & x_22027;
assign x_53317 = x_53315 & x_53316;
assign x_53318 = x_53314 & x_53317;
assign x_53319 = x_22028 & x_22029;
assign x_53320 = x_22030 & x_22031;
assign x_53321 = x_53319 & x_53320;
assign x_53322 = x_22032 & x_22033;
assign x_53323 = x_22034 & x_22035;
assign x_53324 = x_53322 & x_53323;
assign x_53325 = x_53321 & x_53324;
assign x_53326 = x_53318 & x_53325;
assign x_53327 = x_53312 & x_53326;
assign x_53328 = x_22037 & x_22038;
assign x_53329 = x_22036 & x_53328;
assign x_53330 = x_22039 & x_22040;
assign x_53331 = x_22041 & x_22042;
assign x_53332 = x_53330 & x_53331;
assign x_53333 = x_53329 & x_53332;
assign x_53334 = x_22043 & x_22044;
assign x_53335 = x_22045 & x_22046;
assign x_53336 = x_53334 & x_53335;
assign x_53337 = x_22047 & x_22048;
assign x_53338 = x_22049 & x_22050;
assign x_53339 = x_53337 & x_53338;
assign x_53340 = x_53336 & x_53339;
assign x_53341 = x_53333 & x_53340;
assign x_53342 = x_22051 & x_22052;
assign x_53343 = x_22053 & x_22054;
assign x_53344 = x_53342 & x_53343;
assign x_53345 = x_22055 & x_22056;
assign x_53346 = x_22057 & x_22058;
assign x_53347 = x_53345 & x_53346;
assign x_53348 = x_53344 & x_53347;
assign x_53349 = x_22059 & x_22060;
assign x_53350 = x_22061 & x_22062;
assign x_53351 = x_53349 & x_53350;
assign x_53352 = x_22063 & x_22064;
assign x_53353 = x_22065 & x_22066;
assign x_53354 = x_53352 & x_53353;
assign x_53355 = x_53351 & x_53354;
assign x_53356 = x_53348 & x_53355;
assign x_53357 = x_53341 & x_53356;
assign x_53358 = x_53327 & x_53357;
assign x_53359 = x_22068 & x_22069;
assign x_53360 = x_22067 & x_53359;
assign x_53361 = x_22070 & x_22071;
assign x_53362 = x_22072 & x_22073;
assign x_53363 = x_53361 & x_53362;
assign x_53364 = x_53360 & x_53363;
assign x_53365 = x_22074 & x_22075;
assign x_53366 = x_22076 & x_22077;
assign x_53367 = x_53365 & x_53366;
assign x_53368 = x_22078 & x_22079;
assign x_53369 = x_22080 & x_22081;
assign x_53370 = x_53368 & x_53369;
assign x_53371 = x_53367 & x_53370;
assign x_53372 = x_53364 & x_53371;
assign x_53373 = x_22083 & x_22084;
assign x_53374 = x_22082 & x_53373;
assign x_53375 = x_22085 & x_22086;
assign x_53376 = x_22087 & x_22088;
assign x_53377 = x_53375 & x_53376;
assign x_53378 = x_53374 & x_53377;
assign x_53379 = x_22089 & x_22090;
assign x_53380 = x_22091 & x_22092;
assign x_53381 = x_53379 & x_53380;
assign x_53382 = x_22093 & x_22094;
assign x_53383 = x_22095 & x_22096;
assign x_53384 = x_53382 & x_53383;
assign x_53385 = x_53381 & x_53384;
assign x_53386 = x_53378 & x_53385;
assign x_53387 = x_53372 & x_53386;
assign x_53388 = x_22098 & x_22099;
assign x_53389 = x_22097 & x_53388;
assign x_53390 = x_22100 & x_22101;
assign x_53391 = x_22102 & x_22103;
assign x_53392 = x_53390 & x_53391;
assign x_53393 = x_53389 & x_53392;
assign x_53394 = x_22104 & x_22105;
assign x_53395 = x_22106 & x_22107;
assign x_53396 = x_53394 & x_53395;
assign x_53397 = x_22108 & x_22109;
assign x_53398 = x_22110 & x_22111;
assign x_53399 = x_53397 & x_53398;
assign x_53400 = x_53396 & x_53399;
assign x_53401 = x_53393 & x_53400;
assign x_53402 = x_22112 & x_22113;
assign x_53403 = x_22114 & x_22115;
assign x_53404 = x_53402 & x_53403;
assign x_53405 = x_22116 & x_22117;
assign x_53406 = x_22118 & x_22119;
assign x_53407 = x_53405 & x_53406;
assign x_53408 = x_53404 & x_53407;
assign x_53409 = x_22120 & x_22121;
assign x_53410 = x_22122 & x_22123;
assign x_53411 = x_53409 & x_53410;
assign x_53412 = x_22124 & x_22125;
assign x_53413 = x_22126 & x_22127;
assign x_53414 = x_53412 & x_53413;
assign x_53415 = x_53411 & x_53414;
assign x_53416 = x_53408 & x_53415;
assign x_53417 = x_53401 & x_53416;
assign x_53418 = x_53387 & x_53417;
assign x_53419 = x_53358 & x_53418;
assign x_53420 = x_22129 & x_22130;
assign x_53421 = x_22128 & x_53420;
assign x_53422 = x_22131 & x_22132;
assign x_53423 = x_22133 & x_22134;
assign x_53424 = x_53422 & x_53423;
assign x_53425 = x_53421 & x_53424;
assign x_53426 = x_22135 & x_22136;
assign x_53427 = x_22137 & x_22138;
assign x_53428 = x_53426 & x_53427;
assign x_53429 = x_22139 & x_22140;
assign x_53430 = x_22141 & x_22142;
assign x_53431 = x_53429 & x_53430;
assign x_53432 = x_53428 & x_53431;
assign x_53433 = x_53425 & x_53432;
assign x_53434 = x_22144 & x_22145;
assign x_53435 = x_22143 & x_53434;
assign x_53436 = x_22146 & x_22147;
assign x_53437 = x_22148 & x_22149;
assign x_53438 = x_53436 & x_53437;
assign x_53439 = x_53435 & x_53438;
assign x_53440 = x_22150 & x_22151;
assign x_53441 = x_22152 & x_22153;
assign x_53442 = x_53440 & x_53441;
assign x_53443 = x_22154 & x_22155;
assign x_53444 = x_22156 & x_22157;
assign x_53445 = x_53443 & x_53444;
assign x_53446 = x_53442 & x_53445;
assign x_53447 = x_53439 & x_53446;
assign x_53448 = x_53433 & x_53447;
assign x_53449 = x_22159 & x_22160;
assign x_53450 = x_22158 & x_53449;
assign x_53451 = x_22161 & x_22162;
assign x_53452 = x_22163 & x_22164;
assign x_53453 = x_53451 & x_53452;
assign x_53454 = x_53450 & x_53453;
assign x_53455 = x_22165 & x_22166;
assign x_53456 = x_22167 & x_22168;
assign x_53457 = x_53455 & x_53456;
assign x_53458 = x_22169 & x_22170;
assign x_53459 = x_22171 & x_22172;
assign x_53460 = x_53458 & x_53459;
assign x_53461 = x_53457 & x_53460;
assign x_53462 = x_53454 & x_53461;
assign x_53463 = x_22173 & x_22174;
assign x_53464 = x_22175 & x_22176;
assign x_53465 = x_53463 & x_53464;
assign x_53466 = x_22177 & x_22178;
assign x_53467 = x_22179 & x_22180;
assign x_53468 = x_53466 & x_53467;
assign x_53469 = x_53465 & x_53468;
assign x_53470 = x_22181 & x_22182;
assign x_53471 = x_22183 & x_22184;
assign x_53472 = x_53470 & x_53471;
assign x_53473 = x_22185 & x_22186;
assign x_53474 = x_22187 & x_22188;
assign x_53475 = x_53473 & x_53474;
assign x_53476 = x_53472 & x_53475;
assign x_53477 = x_53469 & x_53476;
assign x_53478 = x_53462 & x_53477;
assign x_53479 = x_53448 & x_53478;
assign x_53480 = x_22190 & x_22191;
assign x_53481 = x_22189 & x_53480;
assign x_53482 = x_22192 & x_22193;
assign x_53483 = x_22194 & x_22195;
assign x_53484 = x_53482 & x_53483;
assign x_53485 = x_53481 & x_53484;
assign x_53486 = x_22196 & x_22197;
assign x_53487 = x_22198 & x_22199;
assign x_53488 = x_53486 & x_53487;
assign x_53489 = x_22200 & x_22201;
assign x_53490 = x_22202 & x_22203;
assign x_53491 = x_53489 & x_53490;
assign x_53492 = x_53488 & x_53491;
assign x_53493 = x_53485 & x_53492;
assign x_53494 = x_22205 & x_22206;
assign x_53495 = x_22204 & x_53494;
assign x_53496 = x_22207 & x_22208;
assign x_53497 = x_22209 & x_22210;
assign x_53498 = x_53496 & x_53497;
assign x_53499 = x_53495 & x_53498;
assign x_53500 = x_22211 & x_22212;
assign x_53501 = x_22213 & x_22214;
assign x_53502 = x_53500 & x_53501;
assign x_53503 = x_22215 & x_22216;
assign x_53504 = x_22217 & x_22218;
assign x_53505 = x_53503 & x_53504;
assign x_53506 = x_53502 & x_53505;
assign x_53507 = x_53499 & x_53506;
assign x_53508 = x_53493 & x_53507;
assign x_53509 = x_22220 & x_22221;
assign x_53510 = x_22219 & x_53509;
assign x_53511 = x_22222 & x_22223;
assign x_53512 = x_22224 & x_22225;
assign x_53513 = x_53511 & x_53512;
assign x_53514 = x_53510 & x_53513;
assign x_53515 = x_22226 & x_22227;
assign x_53516 = x_22228 & x_22229;
assign x_53517 = x_53515 & x_53516;
assign x_53518 = x_22230 & x_22231;
assign x_53519 = x_22232 & x_22233;
assign x_53520 = x_53518 & x_53519;
assign x_53521 = x_53517 & x_53520;
assign x_53522 = x_53514 & x_53521;
assign x_53523 = x_22234 & x_22235;
assign x_53524 = x_22236 & x_22237;
assign x_53525 = x_53523 & x_53524;
assign x_53526 = x_22238 & x_22239;
assign x_53527 = x_22240 & x_22241;
assign x_53528 = x_53526 & x_53527;
assign x_53529 = x_53525 & x_53528;
assign x_53530 = x_22242 & x_22243;
assign x_53531 = x_22244 & x_22245;
assign x_53532 = x_53530 & x_53531;
assign x_53533 = x_22246 & x_22247;
assign x_53534 = x_22248 & x_22249;
assign x_53535 = x_53533 & x_53534;
assign x_53536 = x_53532 & x_53535;
assign x_53537 = x_53529 & x_53536;
assign x_53538 = x_53522 & x_53537;
assign x_53539 = x_53508 & x_53538;
assign x_53540 = x_53479 & x_53539;
assign x_53541 = x_53419 & x_53540;
assign x_53542 = x_22251 & x_22252;
assign x_53543 = x_22250 & x_53542;
assign x_53544 = x_22253 & x_22254;
assign x_53545 = x_22255 & x_22256;
assign x_53546 = x_53544 & x_53545;
assign x_53547 = x_53543 & x_53546;
assign x_53548 = x_22257 & x_22258;
assign x_53549 = x_22259 & x_22260;
assign x_53550 = x_53548 & x_53549;
assign x_53551 = x_22261 & x_22262;
assign x_53552 = x_22263 & x_22264;
assign x_53553 = x_53551 & x_53552;
assign x_53554 = x_53550 & x_53553;
assign x_53555 = x_53547 & x_53554;
assign x_53556 = x_22266 & x_22267;
assign x_53557 = x_22265 & x_53556;
assign x_53558 = x_22268 & x_22269;
assign x_53559 = x_22270 & x_22271;
assign x_53560 = x_53558 & x_53559;
assign x_53561 = x_53557 & x_53560;
assign x_53562 = x_22272 & x_22273;
assign x_53563 = x_22274 & x_22275;
assign x_53564 = x_53562 & x_53563;
assign x_53565 = x_22276 & x_22277;
assign x_53566 = x_22278 & x_22279;
assign x_53567 = x_53565 & x_53566;
assign x_53568 = x_53564 & x_53567;
assign x_53569 = x_53561 & x_53568;
assign x_53570 = x_53555 & x_53569;
assign x_53571 = x_22281 & x_22282;
assign x_53572 = x_22280 & x_53571;
assign x_53573 = x_22283 & x_22284;
assign x_53574 = x_22285 & x_22286;
assign x_53575 = x_53573 & x_53574;
assign x_53576 = x_53572 & x_53575;
assign x_53577 = x_22287 & x_22288;
assign x_53578 = x_22289 & x_22290;
assign x_53579 = x_53577 & x_53578;
assign x_53580 = x_22291 & x_22292;
assign x_53581 = x_22293 & x_22294;
assign x_53582 = x_53580 & x_53581;
assign x_53583 = x_53579 & x_53582;
assign x_53584 = x_53576 & x_53583;
assign x_53585 = x_22295 & x_22296;
assign x_53586 = x_22297 & x_22298;
assign x_53587 = x_53585 & x_53586;
assign x_53588 = x_22299 & x_22300;
assign x_53589 = x_22301 & x_22302;
assign x_53590 = x_53588 & x_53589;
assign x_53591 = x_53587 & x_53590;
assign x_53592 = x_22303 & x_22304;
assign x_53593 = x_22305 & x_22306;
assign x_53594 = x_53592 & x_53593;
assign x_53595 = x_22307 & x_22308;
assign x_53596 = x_22309 & x_22310;
assign x_53597 = x_53595 & x_53596;
assign x_53598 = x_53594 & x_53597;
assign x_53599 = x_53591 & x_53598;
assign x_53600 = x_53584 & x_53599;
assign x_53601 = x_53570 & x_53600;
assign x_53602 = x_22312 & x_22313;
assign x_53603 = x_22311 & x_53602;
assign x_53604 = x_22314 & x_22315;
assign x_53605 = x_22316 & x_22317;
assign x_53606 = x_53604 & x_53605;
assign x_53607 = x_53603 & x_53606;
assign x_53608 = x_22318 & x_22319;
assign x_53609 = x_22320 & x_22321;
assign x_53610 = x_53608 & x_53609;
assign x_53611 = x_22322 & x_22323;
assign x_53612 = x_22324 & x_22325;
assign x_53613 = x_53611 & x_53612;
assign x_53614 = x_53610 & x_53613;
assign x_53615 = x_53607 & x_53614;
assign x_53616 = x_22327 & x_22328;
assign x_53617 = x_22326 & x_53616;
assign x_53618 = x_22329 & x_22330;
assign x_53619 = x_22331 & x_22332;
assign x_53620 = x_53618 & x_53619;
assign x_53621 = x_53617 & x_53620;
assign x_53622 = x_22333 & x_22334;
assign x_53623 = x_22335 & x_22336;
assign x_53624 = x_53622 & x_53623;
assign x_53625 = x_22337 & x_22338;
assign x_53626 = x_22339 & x_22340;
assign x_53627 = x_53625 & x_53626;
assign x_53628 = x_53624 & x_53627;
assign x_53629 = x_53621 & x_53628;
assign x_53630 = x_53615 & x_53629;
assign x_53631 = x_22342 & x_22343;
assign x_53632 = x_22341 & x_53631;
assign x_53633 = x_22344 & x_22345;
assign x_53634 = x_22346 & x_22347;
assign x_53635 = x_53633 & x_53634;
assign x_53636 = x_53632 & x_53635;
assign x_53637 = x_22348 & x_22349;
assign x_53638 = x_22350 & x_22351;
assign x_53639 = x_53637 & x_53638;
assign x_53640 = x_22352 & x_22353;
assign x_53641 = x_22354 & x_22355;
assign x_53642 = x_53640 & x_53641;
assign x_53643 = x_53639 & x_53642;
assign x_53644 = x_53636 & x_53643;
assign x_53645 = x_22356 & x_22357;
assign x_53646 = x_22358 & x_22359;
assign x_53647 = x_53645 & x_53646;
assign x_53648 = x_22360 & x_22361;
assign x_53649 = x_22362 & x_22363;
assign x_53650 = x_53648 & x_53649;
assign x_53651 = x_53647 & x_53650;
assign x_53652 = x_22364 & x_22365;
assign x_53653 = x_22366 & x_22367;
assign x_53654 = x_53652 & x_53653;
assign x_53655 = x_22368 & x_22369;
assign x_53656 = x_22370 & x_22371;
assign x_53657 = x_53655 & x_53656;
assign x_53658 = x_53654 & x_53657;
assign x_53659 = x_53651 & x_53658;
assign x_53660 = x_53644 & x_53659;
assign x_53661 = x_53630 & x_53660;
assign x_53662 = x_53601 & x_53661;
assign x_53663 = x_22373 & x_22374;
assign x_53664 = x_22372 & x_53663;
assign x_53665 = x_22375 & x_22376;
assign x_53666 = x_22377 & x_22378;
assign x_53667 = x_53665 & x_53666;
assign x_53668 = x_53664 & x_53667;
assign x_53669 = x_22379 & x_22380;
assign x_53670 = x_22381 & x_22382;
assign x_53671 = x_53669 & x_53670;
assign x_53672 = x_22383 & x_22384;
assign x_53673 = x_22385 & x_22386;
assign x_53674 = x_53672 & x_53673;
assign x_53675 = x_53671 & x_53674;
assign x_53676 = x_53668 & x_53675;
assign x_53677 = x_22388 & x_22389;
assign x_53678 = x_22387 & x_53677;
assign x_53679 = x_22390 & x_22391;
assign x_53680 = x_22392 & x_22393;
assign x_53681 = x_53679 & x_53680;
assign x_53682 = x_53678 & x_53681;
assign x_53683 = x_22394 & x_22395;
assign x_53684 = x_22396 & x_22397;
assign x_53685 = x_53683 & x_53684;
assign x_53686 = x_22398 & x_22399;
assign x_53687 = x_22400 & x_22401;
assign x_53688 = x_53686 & x_53687;
assign x_53689 = x_53685 & x_53688;
assign x_53690 = x_53682 & x_53689;
assign x_53691 = x_53676 & x_53690;
assign x_53692 = x_22403 & x_22404;
assign x_53693 = x_22402 & x_53692;
assign x_53694 = x_22405 & x_22406;
assign x_53695 = x_22407 & x_22408;
assign x_53696 = x_53694 & x_53695;
assign x_53697 = x_53693 & x_53696;
assign x_53698 = x_22409 & x_22410;
assign x_53699 = x_22411 & x_22412;
assign x_53700 = x_53698 & x_53699;
assign x_53701 = x_22413 & x_22414;
assign x_53702 = x_22415 & x_22416;
assign x_53703 = x_53701 & x_53702;
assign x_53704 = x_53700 & x_53703;
assign x_53705 = x_53697 & x_53704;
assign x_53706 = x_22417 & x_22418;
assign x_53707 = x_22419 & x_22420;
assign x_53708 = x_53706 & x_53707;
assign x_53709 = x_22421 & x_22422;
assign x_53710 = x_22423 & x_22424;
assign x_53711 = x_53709 & x_53710;
assign x_53712 = x_53708 & x_53711;
assign x_53713 = x_22425 & x_22426;
assign x_53714 = x_22427 & x_22428;
assign x_53715 = x_53713 & x_53714;
assign x_53716 = x_22429 & x_22430;
assign x_53717 = x_22431 & x_22432;
assign x_53718 = x_53716 & x_53717;
assign x_53719 = x_53715 & x_53718;
assign x_53720 = x_53712 & x_53719;
assign x_53721 = x_53705 & x_53720;
assign x_53722 = x_53691 & x_53721;
assign x_53723 = x_22434 & x_22435;
assign x_53724 = x_22433 & x_53723;
assign x_53725 = x_22436 & x_22437;
assign x_53726 = x_22438 & x_22439;
assign x_53727 = x_53725 & x_53726;
assign x_53728 = x_53724 & x_53727;
assign x_53729 = x_22440 & x_22441;
assign x_53730 = x_22442 & x_22443;
assign x_53731 = x_53729 & x_53730;
assign x_53732 = x_22444 & x_22445;
assign x_53733 = x_22446 & x_22447;
assign x_53734 = x_53732 & x_53733;
assign x_53735 = x_53731 & x_53734;
assign x_53736 = x_53728 & x_53735;
assign x_53737 = x_22448 & x_22449;
assign x_53738 = x_22450 & x_22451;
assign x_53739 = x_53737 & x_53738;
assign x_53740 = x_22452 & x_22453;
assign x_53741 = x_22454 & x_22455;
assign x_53742 = x_53740 & x_53741;
assign x_53743 = x_53739 & x_53742;
assign x_53744 = x_22456 & x_22457;
assign x_53745 = x_22458 & x_22459;
assign x_53746 = x_53744 & x_53745;
assign x_53747 = x_22460 & x_22461;
assign x_53748 = x_22462 & x_22463;
assign x_53749 = x_53747 & x_53748;
assign x_53750 = x_53746 & x_53749;
assign x_53751 = x_53743 & x_53750;
assign x_53752 = x_53736 & x_53751;
assign x_53753 = x_22465 & x_22466;
assign x_53754 = x_22464 & x_53753;
assign x_53755 = x_22467 & x_22468;
assign x_53756 = x_22469 & x_22470;
assign x_53757 = x_53755 & x_53756;
assign x_53758 = x_53754 & x_53757;
assign x_53759 = x_22471 & x_22472;
assign x_53760 = x_22473 & x_22474;
assign x_53761 = x_53759 & x_53760;
assign x_53762 = x_22475 & x_22476;
assign x_53763 = x_22477 & x_22478;
assign x_53764 = x_53762 & x_53763;
assign x_53765 = x_53761 & x_53764;
assign x_53766 = x_53758 & x_53765;
assign x_53767 = x_22479 & x_22480;
assign x_53768 = x_22481 & x_22482;
assign x_53769 = x_53767 & x_53768;
assign x_53770 = x_22483 & x_22484;
assign x_53771 = x_22485 & x_22486;
assign x_53772 = x_53770 & x_53771;
assign x_53773 = x_53769 & x_53772;
assign x_53774 = x_22487 & x_22488;
assign x_53775 = x_22489 & x_22490;
assign x_53776 = x_53774 & x_53775;
assign x_53777 = x_22491 & x_22492;
assign x_53778 = x_22493 & x_22494;
assign x_53779 = x_53777 & x_53778;
assign x_53780 = x_53776 & x_53779;
assign x_53781 = x_53773 & x_53780;
assign x_53782 = x_53766 & x_53781;
assign x_53783 = x_53752 & x_53782;
assign x_53784 = x_53722 & x_53783;
assign x_53785 = x_53662 & x_53784;
assign x_53786 = x_53541 & x_53785;
assign x_53787 = x_53298 & x_53786;
assign x_53788 = x_22496 & x_22497;
assign x_53789 = x_22495 & x_53788;
assign x_53790 = x_22498 & x_22499;
assign x_53791 = x_22500 & x_22501;
assign x_53792 = x_53790 & x_53791;
assign x_53793 = x_53789 & x_53792;
assign x_53794 = x_22502 & x_22503;
assign x_53795 = x_22504 & x_22505;
assign x_53796 = x_53794 & x_53795;
assign x_53797 = x_22506 & x_22507;
assign x_53798 = x_22508 & x_22509;
assign x_53799 = x_53797 & x_53798;
assign x_53800 = x_53796 & x_53799;
assign x_53801 = x_53793 & x_53800;
assign x_53802 = x_22511 & x_22512;
assign x_53803 = x_22510 & x_53802;
assign x_53804 = x_22513 & x_22514;
assign x_53805 = x_22515 & x_22516;
assign x_53806 = x_53804 & x_53805;
assign x_53807 = x_53803 & x_53806;
assign x_53808 = x_22517 & x_22518;
assign x_53809 = x_22519 & x_22520;
assign x_53810 = x_53808 & x_53809;
assign x_53811 = x_22521 & x_22522;
assign x_53812 = x_22523 & x_22524;
assign x_53813 = x_53811 & x_53812;
assign x_53814 = x_53810 & x_53813;
assign x_53815 = x_53807 & x_53814;
assign x_53816 = x_53801 & x_53815;
assign x_53817 = x_22526 & x_22527;
assign x_53818 = x_22525 & x_53817;
assign x_53819 = x_22528 & x_22529;
assign x_53820 = x_22530 & x_22531;
assign x_53821 = x_53819 & x_53820;
assign x_53822 = x_53818 & x_53821;
assign x_53823 = x_22532 & x_22533;
assign x_53824 = x_22534 & x_22535;
assign x_53825 = x_53823 & x_53824;
assign x_53826 = x_22536 & x_22537;
assign x_53827 = x_22538 & x_22539;
assign x_53828 = x_53826 & x_53827;
assign x_53829 = x_53825 & x_53828;
assign x_53830 = x_53822 & x_53829;
assign x_53831 = x_22540 & x_22541;
assign x_53832 = x_22542 & x_22543;
assign x_53833 = x_53831 & x_53832;
assign x_53834 = x_22544 & x_22545;
assign x_53835 = x_22546 & x_22547;
assign x_53836 = x_53834 & x_53835;
assign x_53837 = x_53833 & x_53836;
assign x_53838 = x_22548 & x_22549;
assign x_53839 = x_22550 & x_22551;
assign x_53840 = x_53838 & x_53839;
assign x_53841 = x_22552 & x_22553;
assign x_53842 = x_22554 & x_22555;
assign x_53843 = x_53841 & x_53842;
assign x_53844 = x_53840 & x_53843;
assign x_53845 = x_53837 & x_53844;
assign x_53846 = x_53830 & x_53845;
assign x_53847 = x_53816 & x_53846;
assign x_53848 = x_22557 & x_22558;
assign x_53849 = x_22556 & x_53848;
assign x_53850 = x_22559 & x_22560;
assign x_53851 = x_22561 & x_22562;
assign x_53852 = x_53850 & x_53851;
assign x_53853 = x_53849 & x_53852;
assign x_53854 = x_22563 & x_22564;
assign x_53855 = x_22565 & x_22566;
assign x_53856 = x_53854 & x_53855;
assign x_53857 = x_22567 & x_22568;
assign x_53858 = x_22569 & x_22570;
assign x_53859 = x_53857 & x_53858;
assign x_53860 = x_53856 & x_53859;
assign x_53861 = x_53853 & x_53860;
assign x_53862 = x_22572 & x_22573;
assign x_53863 = x_22571 & x_53862;
assign x_53864 = x_22574 & x_22575;
assign x_53865 = x_22576 & x_22577;
assign x_53866 = x_53864 & x_53865;
assign x_53867 = x_53863 & x_53866;
assign x_53868 = x_22578 & x_22579;
assign x_53869 = x_22580 & x_22581;
assign x_53870 = x_53868 & x_53869;
assign x_53871 = x_22582 & x_22583;
assign x_53872 = x_22584 & x_22585;
assign x_53873 = x_53871 & x_53872;
assign x_53874 = x_53870 & x_53873;
assign x_53875 = x_53867 & x_53874;
assign x_53876 = x_53861 & x_53875;
assign x_53877 = x_22587 & x_22588;
assign x_53878 = x_22586 & x_53877;
assign x_53879 = x_22589 & x_22590;
assign x_53880 = x_22591 & x_22592;
assign x_53881 = x_53879 & x_53880;
assign x_53882 = x_53878 & x_53881;
assign x_53883 = x_22593 & x_22594;
assign x_53884 = x_22595 & x_22596;
assign x_53885 = x_53883 & x_53884;
assign x_53886 = x_22597 & x_22598;
assign x_53887 = x_22599 & x_22600;
assign x_53888 = x_53886 & x_53887;
assign x_53889 = x_53885 & x_53888;
assign x_53890 = x_53882 & x_53889;
assign x_53891 = x_22601 & x_22602;
assign x_53892 = x_22603 & x_22604;
assign x_53893 = x_53891 & x_53892;
assign x_53894 = x_22605 & x_22606;
assign x_53895 = x_22607 & x_22608;
assign x_53896 = x_53894 & x_53895;
assign x_53897 = x_53893 & x_53896;
assign x_53898 = x_22609 & x_22610;
assign x_53899 = x_22611 & x_22612;
assign x_53900 = x_53898 & x_53899;
assign x_53901 = x_22613 & x_22614;
assign x_53902 = x_22615 & x_22616;
assign x_53903 = x_53901 & x_53902;
assign x_53904 = x_53900 & x_53903;
assign x_53905 = x_53897 & x_53904;
assign x_53906 = x_53890 & x_53905;
assign x_53907 = x_53876 & x_53906;
assign x_53908 = x_53847 & x_53907;
assign x_53909 = x_22618 & x_22619;
assign x_53910 = x_22617 & x_53909;
assign x_53911 = x_22620 & x_22621;
assign x_53912 = x_22622 & x_22623;
assign x_53913 = x_53911 & x_53912;
assign x_53914 = x_53910 & x_53913;
assign x_53915 = x_22624 & x_22625;
assign x_53916 = x_22626 & x_22627;
assign x_53917 = x_53915 & x_53916;
assign x_53918 = x_22628 & x_22629;
assign x_53919 = x_22630 & x_22631;
assign x_53920 = x_53918 & x_53919;
assign x_53921 = x_53917 & x_53920;
assign x_53922 = x_53914 & x_53921;
assign x_53923 = x_22633 & x_22634;
assign x_53924 = x_22632 & x_53923;
assign x_53925 = x_22635 & x_22636;
assign x_53926 = x_22637 & x_22638;
assign x_53927 = x_53925 & x_53926;
assign x_53928 = x_53924 & x_53927;
assign x_53929 = x_22639 & x_22640;
assign x_53930 = x_22641 & x_22642;
assign x_53931 = x_53929 & x_53930;
assign x_53932 = x_22643 & x_22644;
assign x_53933 = x_22645 & x_22646;
assign x_53934 = x_53932 & x_53933;
assign x_53935 = x_53931 & x_53934;
assign x_53936 = x_53928 & x_53935;
assign x_53937 = x_53922 & x_53936;
assign x_53938 = x_22648 & x_22649;
assign x_53939 = x_22647 & x_53938;
assign x_53940 = x_22650 & x_22651;
assign x_53941 = x_22652 & x_22653;
assign x_53942 = x_53940 & x_53941;
assign x_53943 = x_53939 & x_53942;
assign x_53944 = x_22654 & x_22655;
assign x_53945 = x_22656 & x_22657;
assign x_53946 = x_53944 & x_53945;
assign x_53947 = x_22658 & x_22659;
assign x_53948 = x_22660 & x_22661;
assign x_53949 = x_53947 & x_53948;
assign x_53950 = x_53946 & x_53949;
assign x_53951 = x_53943 & x_53950;
assign x_53952 = x_22662 & x_22663;
assign x_53953 = x_22664 & x_22665;
assign x_53954 = x_53952 & x_53953;
assign x_53955 = x_22666 & x_22667;
assign x_53956 = x_22668 & x_22669;
assign x_53957 = x_53955 & x_53956;
assign x_53958 = x_53954 & x_53957;
assign x_53959 = x_22670 & x_22671;
assign x_53960 = x_22672 & x_22673;
assign x_53961 = x_53959 & x_53960;
assign x_53962 = x_22674 & x_22675;
assign x_53963 = x_22676 & x_22677;
assign x_53964 = x_53962 & x_53963;
assign x_53965 = x_53961 & x_53964;
assign x_53966 = x_53958 & x_53965;
assign x_53967 = x_53951 & x_53966;
assign x_53968 = x_53937 & x_53967;
assign x_53969 = x_22679 & x_22680;
assign x_53970 = x_22678 & x_53969;
assign x_53971 = x_22681 & x_22682;
assign x_53972 = x_22683 & x_22684;
assign x_53973 = x_53971 & x_53972;
assign x_53974 = x_53970 & x_53973;
assign x_53975 = x_22685 & x_22686;
assign x_53976 = x_22687 & x_22688;
assign x_53977 = x_53975 & x_53976;
assign x_53978 = x_22689 & x_22690;
assign x_53979 = x_22691 & x_22692;
assign x_53980 = x_53978 & x_53979;
assign x_53981 = x_53977 & x_53980;
assign x_53982 = x_53974 & x_53981;
assign x_53983 = x_22694 & x_22695;
assign x_53984 = x_22693 & x_53983;
assign x_53985 = x_22696 & x_22697;
assign x_53986 = x_22698 & x_22699;
assign x_53987 = x_53985 & x_53986;
assign x_53988 = x_53984 & x_53987;
assign x_53989 = x_22700 & x_22701;
assign x_53990 = x_22702 & x_22703;
assign x_53991 = x_53989 & x_53990;
assign x_53992 = x_22704 & x_22705;
assign x_53993 = x_22706 & x_22707;
assign x_53994 = x_53992 & x_53993;
assign x_53995 = x_53991 & x_53994;
assign x_53996 = x_53988 & x_53995;
assign x_53997 = x_53982 & x_53996;
assign x_53998 = x_22709 & x_22710;
assign x_53999 = x_22708 & x_53998;
assign x_54000 = x_22711 & x_22712;
assign x_54001 = x_22713 & x_22714;
assign x_54002 = x_54000 & x_54001;
assign x_54003 = x_53999 & x_54002;
assign x_54004 = x_22715 & x_22716;
assign x_54005 = x_22717 & x_22718;
assign x_54006 = x_54004 & x_54005;
assign x_54007 = x_22719 & x_22720;
assign x_54008 = x_22721 & x_22722;
assign x_54009 = x_54007 & x_54008;
assign x_54010 = x_54006 & x_54009;
assign x_54011 = x_54003 & x_54010;
assign x_54012 = x_22723 & x_22724;
assign x_54013 = x_22725 & x_22726;
assign x_54014 = x_54012 & x_54013;
assign x_54015 = x_22727 & x_22728;
assign x_54016 = x_22729 & x_22730;
assign x_54017 = x_54015 & x_54016;
assign x_54018 = x_54014 & x_54017;
assign x_54019 = x_22731 & x_22732;
assign x_54020 = x_22733 & x_22734;
assign x_54021 = x_54019 & x_54020;
assign x_54022 = x_22735 & x_22736;
assign x_54023 = x_22737 & x_22738;
assign x_54024 = x_54022 & x_54023;
assign x_54025 = x_54021 & x_54024;
assign x_54026 = x_54018 & x_54025;
assign x_54027 = x_54011 & x_54026;
assign x_54028 = x_53997 & x_54027;
assign x_54029 = x_53968 & x_54028;
assign x_54030 = x_53908 & x_54029;
assign x_54031 = x_22740 & x_22741;
assign x_54032 = x_22739 & x_54031;
assign x_54033 = x_22742 & x_22743;
assign x_54034 = x_22744 & x_22745;
assign x_54035 = x_54033 & x_54034;
assign x_54036 = x_54032 & x_54035;
assign x_54037 = x_22746 & x_22747;
assign x_54038 = x_22748 & x_22749;
assign x_54039 = x_54037 & x_54038;
assign x_54040 = x_22750 & x_22751;
assign x_54041 = x_22752 & x_22753;
assign x_54042 = x_54040 & x_54041;
assign x_54043 = x_54039 & x_54042;
assign x_54044 = x_54036 & x_54043;
assign x_54045 = x_22755 & x_22756;
assign x_54046 = x_22754 & x_54045;
assign x_54047 = x_22757 & x_22758;
assign x_54048 = x_22759 & x_22760;
assign x_54049 = x_54047 & x_54048;
assign x_54050 = x_54046 & x_54049;
assign x_54051 = x_22761 & x_22762;
assign x_54052 = x_22763 & x_22764;
assign x_54053 = x_54051 & x_54052;
assign x_54054 = x_22765 & x_22766;
assign x_54055 = x_22767 & x_22768;
assign x_54056 = x_54054 & x_54055;
assign x_54057 = x_54053 & x_54056;
assign x_54058 = x_54050 & x_54057;
assign x_54059 = x_54044 & x_54058;
assign x_54060 = x_22770 & x_22771;
assign x_54061 = x_22769 & x_54060;
assign x_54062 = x_22772 & x_22773;
assign x_54063 = x_22774 & x_22775;
assign x_54064 = x_54062 & x_54063;
assign x_54065 = x_54061 & x_54064;
assign x_54066 = x_22776 & x_22777;
assign x_54067 = x_22778 & x_22779;
assign x_54068 = x_54066 & x_54067;
assign x_54069 = x_22780 & x_22781;
assign x_54070 = x_22782 & x_22783;
assign x_54071 = x_54069 & x_54070;
assign x_54072 = x_54068 & x_54071;
assign x_54073 = x_54065 & x_54072;
assign x_54074 = x_22784 & x_22785;
assign x_54075 = x_22786 & x_22787;
assign x_54076 = x_54074 & x_54075;
assign x_54077 = x_22788 & x_22789;
assign x_54078 = x_22790 & x_22791;
assign x_54079 = x_54077 & x_54078;
assign x_54080 = x_54076 & x_54079;
assign x_54081 = x_22792 & x_22793;
assign x_54082 = x_22794 & x_22795;
assign x_54083 = x_54081 & x_54082;
assign x_54084 = x_22796 & x_22797;
assign x_54085 = x_22798 & x_22799;
assign x_54086 = x_54084 & x_54085;
assign x_54087 = x_54083 & x_54086;
assign x_54088 = x_54080 & x_54087;
assign x_54089 = x_54073 & x_54088;
assign x_54090 = x_54059 & x_54089;
assign x_54091 = x_22801 & x_22802;
assign x_54092 = x_22800 & x_54091;
assign x_54093 = x_22803 & x_22804;
assign x_54094 = x_22805 & x_22806;
assign x_54095 = x_54093 & x_54094;
assign x_54096 = x_54092 & x_54095;
assign x_54097 = x_22807 & x_22808;
assign x_54098 = x_22809 & x_22810;
assign x_54099 = x_54097 & x_54098;
assign x_54100 = x_22811 & x_22812;
assign x_54101 = x_22813 & x_22814;
assign x_54102 = x_54100 & x_54101;
assign x_54103 = x_54099 & x_54102;
assign x_54104 = x_54096 & x_54103;
assign x_54105 = x_22816 & x_22817;
assign x_54106 = x_22815 & x_54105;
assign x_54107 = x_22818 & x_22819;
assign x_54108 = x_22820 & x_22821;
assign x_54109 = x_54107 & x_54108;
assign x_54110 = x_54106 & x_54109;
assign x_54111 = x_22822 & x_22823;
assign x_54112 = x_22824 & x_22825;
assign x_54113 = x_54111 & x_54112;
assign x_54114 = x_22826 & x_22827;
assign x_54115 = x_22828 & x_22829;
assign x_54116 = x_54114 & x_54115;
assign x_54117 = x_54113 & x_54116;
assign x_54118 = x_54110 & x_54117;
assign x_54119 = x_54104 & x_54118;
assign x_54120 = x_22831 & x_22832;
assign x_54121 = x_22830 & x_54120;
assign x_54122 = x_22833 & x_22834;
assign x_54123 = x_22835 & x_22836;
assign x_54124 = x_54122 & x_54123;
assign x_54125 = x_54121 & x_54124;
assign x_54126 = x_22837 & x_22838;
assign x_54127 = x_22839 & x_22840;
assign x_54128 = x_54126 & x_54127;
assign x_54129 = x_22841 & x_22842;
assign x_54130 = x_22843 & x_22844;
assign x_54131 = x_54129 & x_54130;
assign x_54132 = x_54128 & x_54131;
assign x_54133 = x_54125 & x_54132;
assign x_54134 = x_22845 & x_22846;
assign x_54135 = x_22847 & x_22848;
assign x_54136 = x_54134 & x_54135;
assign x_54137 = x_22849 & x_22850;
assign x_54138 = x_22851 & x_22852;
assign x_54139 = x_54137 & x_54138;
assign x_54140 = x_54136 & x_54139;
assign x_54141 = x_22853 & x_22854;
assign x_54142 = x_22855 & x_22856;
assign x_54143 = x_54141 & x_54142;
assign x_54144 = x_22857 & x_22858;
assign x_54145 = x_22859 & x_22860;
assign x_54146 = x_54144 & x_54145;
assign x_54147 = x_54143 & x_54146;
assign x_54148 = x_54140 & x_54147;
assign x_54149 = x_54133 & x_54148;
assign x_54150 = x_54119 & x_54149;
assign x_54151 = x_54090 & x_54150;
assign x_54152 = x_22862 & x_22863;
assign x_54153 = x_22861 & x_54152;
assign x_54154 = x_22864 & x_22865;
assign x_54155 = x_22866 & x_22867;
assign x_54156 = x_54154 & x_54155;
assign x_54157 = x_54153 & x_54156;
assign x_54158 = x_22868 & x_22869;
assign x_54159 = x_22870 & x_22871;
assign x_54160 = x_54158 & x_54159;
assign x_54161 = x_22872 & x_22873;
assign x_54162 = x_22874 & x_22875;
assign x_54163 = x_54161 & x_54162;
assign x_54164 = x_54160 & x_54163;
assign x_54165 = x_54157 & x_54164;
assign x_54166 = x_22877 & x_22878;
assign x_54167 = x_22876 & x_54166;
assign x_54168 = x_22879 & x_22880;
assign x_54169 = x_22881 & x_22882;
assign x_54170 = x_54168 & x_54169;
assign x_54171 = x_54167 & x_54170;
assign x_54172 = x_22883 & x_22884;
assign x_54173 = x_22885 & x_22886;
assign x_54174 = x_54172 & x_54173;
assign x_54175 = x_22887 & x_22888;
assign x_54176 = x_22889 & x_22890;
assign x_54177 = x_54175 & x_54176;
assign x_54178 = x_54174 & x_54177;
assign x_54179 = x_54171 & x_54178;
assign x_54180 = x_54165 & x_54179;
assign x_54181 = x_22892 & x_22893;
assign x_54182 = x_22891 & x_54181;
assign x_54183 = x_22894 & x_22895;
assign x_54184 = x_22896 & x_22897;
assign x_54185 = x_54183 & x_54184;
assign x_54186 = x_54182 & x_54185;
assign x_54187 = x_22898 & x_22899;
assign x_54188 = x_22900 & x_22901;
assign x_54189 = x_54187 & x_54188;
assign x_54190 = x_22902 & x_22903;
assign x_54191 = x_22904 & x_22905;
assign x_54192 = x_54190 & x_54191;
assign x_54193 = x_54189 & x_54192;
assign x_54194 = x_54186 & x_54193;
assign x_54195 = x_22906 & x_22907;
assign x_54196 = x_22908 & x_22909;
assign x_54197 = x_54195 & x_54196;
assign x_54198 = x_22910 & x_22911;
assign x_54199 = x_22912 & x_22913;
assign x_54200 = x_54198 & x_54199;
assign x_54201 = x_54197 & x_54200;
assign x_54202 = x_22914 & x_22915;
assign x_54203 = x_22916 & x_22917;
assign x_54204 = x_54202 & x_54203;
assign x_54205 = x_22918 & x_22919;
assign x_54206 = x_22920 & x_22921;
assign x_54207 = x_54205 & x_54206;
assign x_54208 = x_54204 & x_54207;
assign x_54209 = x_54201 & x_54208;
assign x_54210 = x_54194 & x_54209;
assign x_54211 = x_54180 & x_54210;
assign x_54212 = x_22923 & x_22924;
assign x_54213 = x_22922 & x_54212;
assign x_54214 = x_22925 & x_22926;
assign x_54215 = x_22927 & x_22928;
assign x_54216 = x_54214 & x_54215;
assign x_54217 = x_54213 & x_54216;
assign x_54218 = x_22929 & x_22930;
assign x_54219 = x_22931 & x_22932;
assign x_54220 = x_54218 & x_54219;
assign x_54221 = x_22933 & x_22934;
assign x_54222 = x_22935 & x_22936;
assign x_54223 = x_54221 & x_54222;
assign x_54224 = x_54220 & x_54223;
assign x_54225 = x_54217 & x_54224;
assign x_54226 = x_22937 & x_22938;
assign x_54227 = x_22939 & x_22940;
assign x_54228 = x_54226 & x_54227;
assign x_54229 = x_22941 & x_22942;
assign x_54230 = x_22943 & x_22944;
assign x_54231 = x_54229 & x_54230;
assign x_54232 = x_54228 & x_54231;
assign x_54233 = x_22945 & x_22946;
assign x_54234 = x_22947 & x_22948;
assign x_54235 = x_54233 & x_54234;
assign x_54236 = x_22949 & x_22950;
assign x_54237 = x_22951 & x_22952;
assign x_54238 = x_54236 & x_54237;
assign x_54239 = x_54235 & x_54238;
assign x_54240 = x_54232 & x_54239;
assign x_54241 = x_54225 & x_54240;
assign x_54242 = x_22954 & x_22955;
assign x_54243 = x_22953 & x_54242;
assign x_54244 = x_22956 & x_22957;
assign x_54245 = x_22958 & x_22959;
assign x_54246 = x_54244 & x_54245;
assign x_54247 = x_54243 & x_54246;
assign x_54248 = x_22960 & x_22961;
assign x_54249 = x_22962 & x_22963;
assign x_54250 = x_54248 & x_54249;
assign x_54251 = x_22964 & x_22965;
assign x_54252 = x_22966 & x_22967;
assign x_54253 = x_54251 & x_54252;
assign x_54254 = x_54250 & x_54253;
assign x_54255 = x_54247 & x_54254;
assign x_54256 = x_22968 & x_22969;
assign x_54257 = x_22970 & x_22971;
assign x_54258 = x_54256 & x_54257;
assign x_54259 = x_22972 & x_22973;
assign x_54260 = x_22974 & x_22975;
assign x_54261 = x_54259 & x_54260;
assign x_54262 = x_54258 & x_54261;
assign x_54263 = x_22976 & x_22977;
assign x_54264 = x_22978 & x_22979;
assign x_54265 = x_54263 & x_54264;
assign x_54266 = x_22980 & x_22981;
assign x_54267 = x_22982 & x_22983;
assign x_54268 = x_54266 & x_54267;
assign x_54269 = x_54265 & x_54268;
assign x_54270 = x_54262 & x_54269;
assign x_54271 = x_54255 & x_54270;
assign x_54272 = x_54241 & x_54271;
assign x_54273 = x_54211 & x_54272;
assign x_54274 = x_54151 & x_54273;
assign x_54275 = x_54030 & x_54274;
assign x_54276 = x_22985 & x_22986;
assign x_54277 = x_22984 & x_54276;
assign x_54278 = x_22987 & x_22988;
assign x_54279 = x_22989 & x_22990;
assign x_54280 = x_54278 & x_54279;
assign x_54281 = x_54277 & x_54280;
assign x_54282 = x_22991 & x_22992;
assign x_54283 = x_22993 & x_22994;
assign x_54284 = x_54282 & x_54283;
assign x_54285 = x_22995 & x_22996;
assign x_54286 = x_22997 & x_22998;
assign x_54287 = x_54285 & x_54286;
assign x_54288 = x_54284 & x_54287;
assign x_54289 = x_54281 & x_54288;
assign x_54290 = x_23000 & x_23001;
assign x_54291 = x_22999 & x_54290;
assign x_54292 = x_23002 & x_23003;
assign x_54293 = x_23004 & x_23005;
assign x_54294 = x_54292 & x_54293;
assign x_54295 = x_54291 & x_54294;
assign x_54296 = x_23006 & x_23007;
assign x_54297 = x_23008 & x_23009;
assign x_54298 = x_54296 & x_54297;
assign x_54299 = x_23010 & x_23011;
assign x_54300 = x_23012 & x_23013;
assign x_54301 = x_54299 & x_54300;
assign x_54302 = x_54298 & x_54301;
assign x_54303 = x_54295 & x_54302;
assign x_54304 = x_54289 & x_54303;
assign x_54305 = x_23015 & x_23016;
assign x_54306 = x_23014 & x_54305;
assign x_54307 = x_23017 & x_23018;
assign x_54308 = x_23019 & x_23020;
assign x_54309 = x_54307 & x_54308;
assign x_54310 = x_54306 & x_54309;
assign x_54311 = x_23021 & x_23022;
assign x_54312 = x_23023 & x_23024;
assign x_54313 = x_54311 & x_54312;
assign x_54314 = x_23025 & x_23026;
assign x_54315 = x_23027 & x_23028;
assign x_54316 = x_54314 & x_54315;
assign x_54317 = x_54313 & x_54316;
assign x_54318 = x_54310 & x_54317;
assign x_54319 = x_23029 & x_23030;
assign x_54320 = x_23031 & x_23032;
assign x_54321 = x_54319 & x_54320;
assign x_54322 = x_23033 & x_23034;
assign x_54323 = x_23035 & x_23036;
assign x_54324 = x_54322 & x_54323;
assign x_54325 = x_54321 & x_54324;
assign x_54326 = x_23037 & x_23038;
assign x_54327 = x_23039 & x_23040;
assign x_54328 = x_54326 & x_54327;
assign x_54329 = x_23041 & x_23042;
assign x_54330 = x_23043 & x_23044;
assign x_54331 = x_54329 & x_54330;
assign x_54332 = x_54328 & x_54331;
assign x_54333 = x_54325 & x_54332;
assign x_54334 = x_54318 & x_54333;
assign x_54335 = x_54304 & x_54334;
assign x_54336 = x_23046 & x_23047;
assign x_54337 = x_23045 & x_54336;
assign x_54338 = x_23048 & x_23049;
assign x_54339 = x_23050 & x_23051;
assign x_54340 = x_54338 & x_54339;
assign x_54341 = x_54337 & x_54340;
assign x_54342 = x_23052 & x_23053;
assign x_54343 = x_23054 & x_23055;
assign x_54344 = x_54342 & x_54343;
assign x_54345 = x_23056 & x_23057;
assign x_54346 = x_23058 & x_23059;
assign x_54347 = x_54345 & x_54346;
assign x_54348 = x_54344 & x_54347;
assign x_54349 = x_54341 & x_54348;
assign x_54350 = x_23061 & x_23062;
assign x_54351 = x_23060 & x_54350;
assign x_54352 = x_23063 & x_23064;
assign x_54353 = x_23065 & x_23066;
assign x_54354 = x_54352 & x_54353;
assign x_54355 = x_54351 & x_54354;
assign x_54356 = x_23067 & x_23068;
assign x_54357 = x_23069 & x_23070;
assign x_54358 = x_54356 & x_54357;
assign x_54359 = x_23071 & x_23072;
assign x_54360 = x_23073 & x_23074;
assign x_54361 = x_54359 & x_54360;
assign x_54362 = x_54358 & x_54361;
assign x_54363 = x_54355 & x_54362;
assign x_54364 = x_54349 & x_54363;
assign x_54365 = x_23076 & x_23077;
assign x_54366 = x_23075 & x_54365;
assign x_54367 = x_23078 & x_23079;
assign x_54368 = x_23080 & x_23081;
assign x_54369 = x_54367 & x_54368;
assign x_54370 = x_54366 & x_54369;
assign x_54371 = x_23082 & x_23083;
assign x_54372 = x_23084 & x_23085;
assign x_54373 = x_54371 & x_54372;
assign x_54374 = x_23086 & x_23087;
assign x_54375 = x_23088 & x_23089;
assign x_54376 = x_54374 & x_54375;
assign x_54377 = x_54373 & x_54376;
assign x_54378 = x_54370 & x_54377;
assign x_54379 = x_23090 & x_23091;
assign x_54380 = x_23092 & x_23093;
assign x_54381 = x_54379 & x_54380;
assign x_54382 = x_23094 & x_23095;
assign x_54383 = x_23096 & x_23097;
assign x_54384 = x_54382 & x_54383;
assign x_54385 = x_54381 & x_54384;
assign x_54386 = x_23098 & x_23099;
assign x_54387 = x_23100 & x_23101;
assign x_54388 = x_54386 & x_54387;
assign x_54389 = x_23102 & x_23103;
assign x_54390 = x_23104 & x_23105;
assign x_54391 = x_54389 & x_54390;
assign x_54392 = x_54388 & x_54391;
assign x_54393 = x_54385 & x_54392;
assign x_54394 = x_54378 & x_54393;
assign x_54395 = x_54364 & x_54394;
assign x_54396 = x_54335 & x_54395;
assign x_54397 = x_23107 & x_23108;
assign x_54398 = x_23106 & x_54397;
assign x_54399 = x_23109 & x_23110;
assign x_54400 = x_23111 & x_23112;
assign x_54401 = x_54399 & x_54400;
assign x_54402 = x_54398 & x_54401;
assign x_54403 = x_23113 & x_23114;
assign x_54404 = x_23115 & x_23116;
assign x_54405 = x_54403 & x_54404;
assign x_54406 = x_23117 & x_23118;
assign x_54407 = x_23119 & x_23120;
assign x_54408 = x_54406 & x_54407;
assign x_54409 = x_54405 & x_54408;
assign x_54410 = x_54402 & x_54409;
assign x_54411 = x_23122 & x_23123;
assign x_54412 = x_23121 & x_54411;
assign x_54413 = x_23124 & x_23125;
assign x_54414 = x_23126 & x_23127;
assign x_54415 = x_54413 & x_54414;
assign x_54416 = x_54412 & x_54415;
assign x_54417 = x_23128 & x_23129;
assign x_54418 = x_23130 & x_23131;
assign x_54419 = x_54417 & x_54418;
assign x_54420 = x_23132 & x_23133;
assign x_54421 = x_23134 & x_23135;
assign x_54422 = x_54420 & x_54421;
assign x_54423 = x_54419 & x_54422;
assign x_54424 = x_54416 & x_54423;
assign x_54425 = x_54410 & x_54424;
assign x_54426 = x_23137 & x_23138;
assign x_54427 = x_23136 & x_54426;
assign x_54428 = x_23139 & x_23140;
assign x_54429 = x_23141 & x_23142;
assign x_54430 = x_54428 & x_54429;
assign x_54431 = x_54427 & x_54430;
assign x_54432 = x_23143 & x_23144;
assign x_54433 = x_23145 & x_23146;
assign x_54434 = x_54432 & x_54433;
assign x_54435 = x_23147 & x_23148;
assign x_54436 = x_23149 & x_23150;
assign x_54437 = x_54435 & x_54436;
assign x_54438 = x_54434 & x_54437;
assign x_54439 = x_54431 & x_54438;
assign x_54440 = x_23151 & x_23152;
assign x_54441 = x_23153 & x_23154;
assign x_54442 = x_54440 & x_54441;
assign x_54443 = x_23155 & x_23156;
assign x_54444 = x_23157 & x_23158;
assign x_54445 = x_54443 & x_54444;
assign x_54446 = x_54442 & x_54445;
assign x_54447 = x_23159 & x_23160;
assign x_54448 = x_23161 & x_23162;
assign x_54449 = x_54447 & x_54448;
assign x_54450 = x_23163 & x_23164;
assign x_54451 = x_23165 & x_23166;
assign x_54452 = x_54450 & x_54451;
assign x_54453 = x_54449 & x_54452;
assign x_54454 = x_54446 & x_54453;
assign x_54455 = x_54439 & x_54454;
assign x_54456 = x_54425 & x_54455;
assign x_54457 = x_23168 & x_23169;
assign x_54458 = x_23167 & x_54457;
assign x_54459 = x_23170 & x_23171;
assign x_54460 = x_23172 & x_23173;
assign x_54461 = x_54459 & x_54460;
assign x_54462 = x_54458 & x_54461;
assign x_54463 = x_23174 & x_23175;
assign x_54464 = x_23176 & x_23177;
assign x_54465 = x_54463 & x_54464;
assign x_54466 = x_23178 & x_23179;
assign x_54467 = x_23180 & x_23181;
assign x_54468 = x_54466 & x_54467;
assign x_54469 = x_54465 & x_54468;
assign x_54470 = x_54462 & x_54469;
assign x_54471 = x_23183 & x_23184;
assign x_54472 = x_23182 & x_54471;
assign x_54473 = x_23185 & x_23186;
assign x_54474 = x_23187 & x_23188;
assign x_54475 = x_54473 & x_54474;
assign x_54476 = x_54472 & x_54475;
assign x_54477 = x_23189 & x_23190;
assign x_54478 = x_23191 & x_23192;
assign x_54479 = x_54477 & x_54478;
assign x_54480 = x_23193 & x_23194;
assign x_54481 = x_23195 & x_23196;
assign x_54482 = x_54480 & x_54481;
assign x_54483 = x_54479 & x_54482;
assign x_54484 = x_54476 & x_54483;
assign x_54485 = x_54470 & x_54484;
assign x_54486 = x_23198 & x_23199;
assign x_54487 = x_23197 & x_54486;
assign x_54488 = x_23200 & x_23201;
assign x_54489 = x_23202 & x_23203;
assign x_54490 = x_54488 & x_54489;
assign x_54491 = x_54487 & x_54490;
assign x_54492 = x_23204 & x_23205;
assign x_54493 = x_23206 & x_23207;
assign x_54494 = x_54492 & x_54493;
assign x_54495 = x_23208 & x_23209;
assign x_54496 = x_23210 & x_23211;
assign x_54497 = x_54495 & x_54496;
assign x_54498 = x_54494 & x_54497;
assign x_54499 = x_54491 & x_54498;
assign x_54500 = x_23212 & x_23213;
assign x_54501 = x_23214 & x_23215;
assign x_54502 = x_54500 & x_54501;
assign x_54503 = x_23216 & x_23217;
assign x_54504 = x_23218 & x_23219;
assign x_54505 = x_54503 & x_54504;
assign x_54506 = x_54502 & x_54505;
assign x_54507 = x_23220 & x_23221;
assign x_54508 = x_23222 & x_23223;
assign x_54509 = x_54507 & x_54508;
assign x_54510 = x_23224 & x_23225;
assign x_54511 = x_23226 & x_23227;
assign x_54512 = x_54510 & x_54511;
assign x_54513 = x_54509 & x_54512;
assign x_54514 = x_54506 & x_54513;
assign x_54515 = x_54499 & x_54514;
assign x_54516 = x_54485 & x_54515;
assign x_54517 = x_54456 & x_54516;
assign x_54518 = x_54396 & x_54517;
assign x_54519 = x_23229 & x_23230;
assign x_54520 = x_23228 & x_54519;
assign x_54521 = x_23231 & x_23232;
assign x_54522 = x_23233 & x_23234;
assign x_54523 = x_54521 & x_54522;
assign x_54524 = x_54520 & x_54523;
assign x_54525 = x_23235 & x_23236;
assign x_54526 = x_23237 & x_23238;
assign x_54527 = x_54525 & x_54526;
assign x_54528 = x_23239 & x_23240;
assign x_54529 = x_23241 & x_23242;
assign x_54530 = x_54528 & x_54529;
assign x_54531 = x_54527 & x_54530;
assign x_54532 = x_54524 & x_54531;
assign x_54533 = x_23244 & x_23245;
assign x_54534 = x_23243 & x_54533;
assign x_54535 = x_23246 & x_23247;
assign x_54536 = x_23248 & x_23249;
assign x_54537 = x_54535 & x_54536;
assign x_54538 = x_54534 & x_54537;
assign x_54539 = x_23250 & x_23251;
assign x_54540 = x_23252 & x_23253;
assign x_54541 = x_54539 & x_54540;
assign x_54542 = x_23254 & x_23255;
assign x_54543 = x_23256 & x_23257;
assign x_54544 = x_54542 & x_54543;
assign x_54545 = x_54541 & x_54544;
assign x_54546 = x_54538 & x_54545;
assign x_54547 = x_54532 & x_54546;
assign x_54548 = x_23259 & x_23260;
assign x_54549 = x_23258 & x_54548;
assign x_54550 = x_23261 & x_23262;
assign x_54551 = x_23263 & x_23264;
assign x_54552 = x_54550 & x_54551;
assign x_54553 = x_54549 & x_54552;
assign x_54554 = x_23265 & x_23266;
assign x_54555 = x_23267 & x_23268;
assign x_54556 = x_54554 & x_54555;
assign x_54557 = x_23269 & x_23270;
assign x_54558 = x_23271 & x_23272;
assign x_54559 = x_54557 & x_54558;
assign x_54560 = x_54556 & x_54559;
assign x_54561 = x_54553 & x_54560;
assign x_54562 = x_23273 & x_23274;
assign x_54563 = x_23275 & x_23276;
assign x_54564 = x_54562 & x_54563;
assign x_54565 = x_23277 & x_23278;
assign x_54566 = x_23279 & x_23280;
assign x_54567 = x_54565 & x_54566;
assign x_54568 = x_54564 & x_54567;
assign x_54569 = x_23281 & x_23282;
assign x_54570 = x_23283 & x_23284;
assign x_54571 = x_54569 & x_54570;
assign x_54572 = x_23285 & x_23286;
assign x_54573 = x_23287 & x_23288;
assign x_54574 = x_54572 & x_54573;
assign x_54575 = x_54571 & x_54574;
assign x_54576 = x_54568 & x_54575;
assign x_54577 = x_54561 & x_54576;
assign x_54578 = x_54547 & x_54577;
assign x_54579 = x_23290 & x_23291;
assign x_54580 = x_23289 & x_54579;
assign x_54581 = x_23292 & x_23293;
assign x_54582 = x_23294 & x_23295;
assign x_54583 = x_54581 & x_54582;
assign x_54584 = x_54580 & x_54583;
assign x_54585 = x_23296 & x_23297;
assign x_54586 = x_23298 & x_23299;
assign x_54587 = x_54585 & x_54586;
assign x_54588 = x_23300 & x_23301;
assign x_54589 = x_23302 & x_23303;
assign x_54590 = x_54588 & x_54589;
assign x_54591 = x_54587 & x_54590;
assign x_54592 = x_54584 & x_54591;
assign x_54593 = x_23305 & x_23306;
assign x_54594 = x_23304 & x_54593;
assign x_54595 = x_23307 & x_23308;
assign x_54596 = x_23309 & x_23310;
assign x_54597 = x_54595 & x_54596;
assign x_54598 = x_54594 & x_54597;
assign x_54599 = x_23311 & x_23312;
assign x_54600 = x_23313 & x_23314;
assign x_54601 = x_54599 & x_54600;
assign x_54602 = x_23315 & x_23316;
assign x_54603 = x_23317 & x_23318;
assign x_54604 = x_54602 & x_54603;
assign x_54605 = x_54601 & x_54604;
assign x_54606 = x_54598 & x_54605;
assign x_54607 = x_54592 & x_54606;
assign x_54608 = x_23320 & x_23321;
assign x_54609 = x_23319 & x_54608;
assign x_54610 = x_23322 & x_23323;
assign x_54611 = x_23324 & x_23325;
assign x_54612 = x_54610 & x_54611;
assign x_54613 = x_54609 & x_54612;
assign x_54614 = x_23326 & x_23327;
assign x_54615 = x_23328 & x_23329;
assign x_54616 = x_54614 & x_54615;
assign x_54617 = x_23330 & x_23331;
assign x_54618 = x_23332 & x_23333;
assign x_54619 = x_54617 & x_54618;
assign x_54620 = x_54616 & x_54619;
assign x_54621 = x_54613 & x_54620;
assign x_54622 = x_23334 & x_23335;
assign x_54623 = x_23336 & x_23337;
assign x_54624 = x_54622 & x_54623;
assign x_54625 = x_23338 & x_23339;
assign x_54626 = x_23340 & x_23341;
assign x_54627 = x_54625 & x_54626;
assign x_54628 = x_54624 & x_54627;
assign x_54629 = x_23342 & x_23343;
assign x_54630 = x_23344 & x_23345;
assign x_54631 = x_54629 & x_54630;
assign x_54632 = x_23346 & x_23347;
assign x_54633 = x_23348 & x_23349;
assign x_54634 = x_54632 & x_54633;
assign x_54635 = x_54631 & x_54634;
assign x_54636 = x_54628 & x_54635;
assign x_54637 = x_54621 & x_54636;
assign x_54638 = x_54607 & x_54637;
assign x_54639 = x_54578 & x_54638;
assign x_54640 = x_23351 & x_23352;
assign x_54641 = x_23350 & x_54640;
assign x_54642 = x_23353 & x_23354;
assign x_54643 = x_23355 & x_23356;
assign x_54644 = x_54642 & x_54643;
assign x_54645 = x_54641 & x_54644;
assign x_54646 = x_23357 & x_23358;
assign x_54647 = x_23359 & x_23360;
assign x_54648 = x_54646 & x_54647;
assign x_54649 = x_23361 & x_23362;
assign x_54650 = x_23363 & x_23364;
assign x_54651 = x_54649 & x_54650;
assign x_54652 = x_54648 & x_54651;
assign x_54653 = x_54645 & x_54652;
assign x_54654 = x_23366 & x_23367;
assign x_54655 = x_23365 & x_54654;
assign x_54656 = x_23368 & x_23369;
assign x_54657 = x_23370 & x_23371;
assign x_54658 = x_54656 & x_54657;
assign x_54659 = x_54655 & x_54658;
assign x_54660 = x_23372 & x_23373;
assign x_54661 = x_23374 & x_23375;
assign x_54662 = x_54660 & x_54661;
assign x_54663 = x_23376 & x_23377;
assign x_54664 = x_23378 & x_23379;
assign x_54665 = x_54663 & x_54664;
assign x_54666 = x_54662 & x_54665;
assign x_54667 = x_54659 & x_54666;
assign x_54668 = x_54653 & x_54667;
assign x_54669 = x_23381 & x_23382;
assign x_54670 = x_23380 & x_54669;
assign x_54671 = x_23383 & x_23384;
assign x_54672 = x_23385 & x_23386;
assign x_54673 = x_54671 & x_54672;
assign x_54674 = x_54670 & x_54673;
assign x_54675 = x_23387 & x_23388;
assign x_54676 = x_23389 & x_23390;
assign x_54677 = x_54675 & x_54676;
assign x_54678 = x_23391 & x_23392;
assign x_54679 = x_23393 & x_23394;
assign x_54680 = x_54678 & x_54679;
assign x_54681 = x_54677 & x_54680;
assign x_54682 = x_54674 & x_54681;
assign x_54683 = x_23395 & x_23396;
assign x_54684 = x_23397 & x_23398;
assign x_54685 = x_54683 & x_54684;
assign x_54686 = x_23399 & x_23400;
assign x_54687 = x_23401 & x_23402;
assign x_54688 = x_54686 & x_54687;
assign x_54689 = x_54685 & x_54688;
assign x_54690 = x_23403 & x_23404;
assign x_54691 = x_23405 & x_23406;
assign x_54692 = x_54690 & x_54691;
assign x_54693 = x_23407 & x_23408;
assign x_54694 = x_23409 & x_23410;
assign x_54695 = x_54693 & x_54694;
assign x_54696 = x_54692 & x_54695;
assign x_54697 = x_54689 & x_54696;
assign x_54698 = x_54682 & x_54697;
assign x_54699 = x_54668 & x_54698;
assign x_54700 = x_23412 & x_23413;
assign x_54701 = x_23411 & x_54700;
assign x_54702 = x_23414 & x_23415;
assign x_54703 = x_23416 & x_23417;
assign x_54704 = x_54702 & x_54703;
assign x_54705 = x_54701 & x_54704;
assign x_54706 = x_23418 & x_23419;
assign x_54707 = x_23420 & x_23421;
assign x_54708 = x_54706 & x_54707;
assign x_54709 = x_23422 & x_23423;
assign x_54710 = x_23424 & x_23425;
assign x_54711 = x_54709 & x_54710;
assign x_54712 = x_54708 & x_54711;
assign x_54713 = x_54705 & x_54712;
assign x_54714 = x_23426 & x_23427;
assign x_54715 = x_23428 & x_23429;
assign x_54716 = x_54714 & x_54715;
assign x_54717 = x_23430 & x_23431;
assign x_54718 = x_23432 & x_23433;
assign x_54719 = x_54717 & x_54718;
assign x_54720 = x_54716 & x_54719;
assign x_54721 = x_23434 & x_23435;
assign x_54722 = x_23436 & x_23437;
assign x_54723 = x_54721 & x_54722;
assign x_54724 = x_23438 & x_23439;
assign x_54725 = x_23440 & x_23441;
assign x_54726 = x_54724 & x_54725;
assign x_54727 = x_54723 & x_54726;
assign x_54728 = x_54720 & x_54727;
assign x_54729 = x_54713 & x_54728;
assign x_54730 = x_23443 & x_23444;
assign x_54731 = x_23442 & x_54730;
assign x_54732 = x_23445 & x_23446;
assign x_54733 = x_23447 & x_23448;
assign x_54734 = x_54732 & x_54733;
assign x_54735 = x_54731 & x_54734;
assign x_54736 = x_23449 & x_23450;
assign x_54737 = x_23451 & x_23452;
assign x_54738 = x_54736 & x_54737;
assign x_54739 = x_23453 & x_23454;
assign x_54740 = x_23455 & x_23456;
assign x_54741 = x_54739 & x_54740;
assign x_54742 = x_54738 & x_54741;
assign x_54743 = x_54735 & x_54742;
assign x_54744 = x_23457 & x_23458;
assign x_54745 = x_23459 & x_23460;
assign x_54746 = x_54744 & x_54745;
assign x_54747 = x_23461 & x_23462;
assign x_54748 = x_23463 & x_23464;
assign x_54749 = x_54747 & x_54748;
assign x_54750 = x_54746 & x_54749;
assign x_54751 = x_23465 & x_23466;
assign x_54752 = x_23467 & x_23468;
assign x_54753 = x_54751 & x_54752;
assign x_54754 = x_23469 & x_23470;
assign x_54755 = x_23471 & x_23472;
assign x_54756 = x_54754 & x_54755;
assign x_54757 = x_54753 & x_54756;
assign x_54758 = x_54750 & x_54757;
assign x_54759 = x_54743 & x_54758;
assign x_54760 = x_54729 & x_54759;
assign x_54761 = x_54699 & x_54760;
assign x_54762 = x_54639 & x_54761;
assign x_54763 = x_54518 & x_54762;
assign x_54764 = x_54275 & x_54763;
assign x_54765 = x_53787 & x_54764;
assign x_54766 = x_52810 & x_54765;
assign x_54767 = x_50855 & x_54766;
assign x_54768 = x_23474 & x_23475;
assign x_54769 = x_23473 & x_54768;
assign x_54770 = x_23476 & x_23477;
assign x_54771 = x_23478 & x_23479;
assign x_54772 = x_54770 & x_54771;
assign x_54773 = x_54769 & x_54772;
assign x_54774 = x_23480 & x_23481;
assign x_54775 = x_23482 & x_23483;
assign x_54776 = x_54774 & x_54775;
assign x_54777 = x_23484 & x_23485;
assign x_54778 = x_23486 & x_23487;
assign x_54779 = x_54777 & x_54778;
assign x_54780 = x_54776 & x_54779;
assign x_54781 = x_54773 & x_54780;
assign x_54782 = x_23489 & x_23490;
assign x_54783 = x_23488 & x_54782;
assign x_54784 = x_23491 & x_23492;
assign x_54785 = x_23493 & x_23494;
assign x_54786 = x_54784 & x_54785;
assign x_54787 = x_54783 & x_54786;
assign x_54788 = x_23495 & x_23496;
assign x_54789 = x_23497 & x_23498;
assign x_54790 = x_54788 & x_54789;
assign x_54791 = x_23499 & x_23500;
assign x_54792 = x_23501 & x_23502;
assign x_54793 = x_54791 & x_54792;
assign x_54794 = x_54790 & x_54793;
assign x_54795 = x_54787 & x_54794;
assign x_54796 = x_54781 & x_54795;
assign x_54797 = x_23504 & x_23505;
assign x_54798 = x_23503 & x_54797;
assign x_54799 = x_23506 & x_23507;
assign x_54800 = x_23508 & x_23509;
assign x_54801 = x_54799 & x_54800;
assign x_54802 = x_54798 & x_54801;
assign x_54803 = x_23510 & x_23511;
assign x_54804 = x_23512 & x_23513;
assign x_54805 = x_54803 & x_54804;
assign x_54806 = x_23514 & x_23515;
assign x_54807 = x_23516 & x_23517;
assign x_54808 = x_54806 & x_54807;
assign x_54809 = x_54805 & x_54808;
assign x_54810 = x_54802 & x_54809;
assign x_54811 = x_23518 & x_23519;
assign x_54812 = x_23520 & x_23521;
assign x_54813 = x_54811 & x_54812;
assign x_54814 = x_23522 & x_23523;
assign x_54815 = x_23524 & x_23525;
assign x_54816 = x_54814 & x_54815;
assign x_54817 = x_54813 & x_54816;
assign x_54818 = x_23526 & x_23527;
assign x_54819 = x_23528 & x_23529;
assign x_54820 = x_54818 & x_54819;
assign x_54821 = x_23530 & x_23531;
assign x_54822 = x_23532 & x_23533;
assign x_54823 = x_54821 & x_54822;
assign x_54824 = x_54820 & x_54823;
assign x_54825 = x_54817 & x_54824;
assign x_54826 = x_54810 & x_54825;
assign x_54827 = x_54796 & x_54826;
assign x_54828 = x_23535 & x_23536;
assign x_54829 = x_23534 & x_54828;
assign x_54830 = x_23537 & x_23538;
assign x_54831 = x_23539 & x_23540;
assign x_54832 = x_54830 & x_54831;
assign x_54833 = x_54829 & x_54832;
assign x_54834 = x_23541 & x_23542;
assign x_54835 = x_23543 & x_23544;
assign x_54836 = x_54834 & x_54835;
assign x_54837 = x_23545 & x_23546;
assign x_54838 = x_23547 & x_23548;
assign x_54839 = x_54837 & x_54838;
assign x_54840 = x_54836 & x_54839;
assign x_54841 = x_54833 & x_54840;
assign x_54842 = x_23550 & x_23551;
assign x_54843 = x_23549 & x_54842;
assign x_54844 = x_23552 & x_23553;
assign x_54845 = x_23554 & x_23555;
assign x_54846 = x_54844 & x_54845;
assign x_54847 = x_54843 & x_54846;
assign x_54848 = x_23556 & x_23557;
assign x_54849 = x_23558 & x_23559;
assign x_54850 = x_54848 & x_54849;
assign x_54851 = x_23560 & x_23561;
assign x_54852 = x_23562 & x_23563;
assign x_54853 = x_54851 & x_54852;
assign x_54854 = x_54850 & x_54853;
assign x_54855 = x_54847 & x_54854;
assign x_54856 = x_54841 & x_54855;
assign x_54857 = x_23565 & x_23566;
assign x_54858 = x_23564 & x_54857;
assign x_54859 = x_23567 & x_23568;
assign x_54860 = x_23569 & x_23570;
assign x_54861 = x_54859 & x_54860;
assign x_54862 = x_54858 & x_54861;
assign x_54863 = x_23571 & x_23572;
assign x_54864 = x_23573 & x_23574;
assign x_54865 = x_54863 & x_54864;
assign x_54866 = x_23575 & x_23576;
assign x_54867 = x_23577 & x_23578;
assign x_54868 = x_54866 & x_54867;
assign x_54869 = x_54865 & x_54868;
assign x_54870 = x_54862 & x_54869;
assign x_54871 = x_23579 & x_23580;
assign x_54872 = x_23581 & x_23582;
assign x_54873 = x_54871 & x_54872;
assign x_54874 = x_23583 & x_23584;
assign x_54875 = x_23585 & x_23586;
assign x_54876 = x_54874 & x_54875;
assign x_54877 = x_54873 & x_54876;
assign x_54878 = x_23587 & x_23588;
assign x_54879 = x_23589 & x_23590;
assign x_54880 = x_54878 & x_54879;
assign x_54881 = x_23591 & x_23592;
assign x_54882 = x_23593 & x_23594;
assign x_54883 = x_54881 & x_54882;
assign x_54884 = x_54880 & x_54883;
assign x_54885 = x_54877 & x_54884;
assign x_54886 = x_54870 & x_54885;
assign x_54887 = x_54856 & x_54886;
assign x_54888 = x_54827 & x_54887;
assign x_54889 = x_23596 & x_23597;
assign x_54890 = x_23595 & x_54889;
assign x_54891 = x_23598 & x_23599;
assign x_54892 = x_23600 & x_23601;
assign x_54893 = x_54891 & x_54892;
assign x_54894 = x_54890 & x_54893;
assign x_54895 = x_23602 & x_23603;
assign x_54896 = x_23604 & x_23605;
assign x_54897 = x_54895 & x_54896;
assign x_54898 = x_23606 & x_23607;
assign x_54899 = x_23608 & x_23609;
assign x_54900 = x_54898 & x_54899;
assign x_54901 = x_54897 & x_54900;
assign x_54902 = x_54894 & x_54901;
assign x_54903 = x_23611 & x_23612;
assign x_54904 = x_23610 & x_54903;
assign x_54905 = x_23613 & x_23614;
assign x_54906 = x_23615 & x_23616;
assign x_54907 = x_54905 & x_54906;
assign x_54908 = x_54904 & x_54907;
assign x_54909 = x_23617 & x_23618;
assign x_54910 = x_23619 & x_23620;
assign x_54911 = x_54909 & x_54910;
assign x_54912 = x_23621 & x_23622;
assign x_54913 = x_23623 & x_23624;
assign x_54914 = x_54912 & x_54913;
assign x_54915 = x_54911 & x_54914;
assign x_54916 = x_54908 & x_54915;
assign x_54917 = x_54902 & x_54916;
assign x_54918 = x_23626 & x_23627;
assign x_54919 = x_23625 & x_54918;
assign x_54920 = x_23628 & x_23629;
assign x_54921 = x_23630 & x_23631;
assign x_54922 = x_54920 & x_54921;
assign x_54923 = x_54919 & x_54922;
assign x_54924 = x_23632 & x_23633;
assign x_54925 = x_23634 & x_23635;
assign x_54926 = x_54924 & x_54925;
assign x_54927 = x_23636 & x_23637;
assign x_54928 = x_23638 & x_23639;
assign x_54929 = x_54927 & x_54928;
assign x_54930 = x_54926 & x_54929;
assign x_54931 = x_54923 & x_54930;
assign x_54932 = x_23640 & x_23641;
assign x_54933 = x_23642 & x_23643;
assign x_54934 = x_54932 & x_54933;
assign x_54935 = x_23644 & x_23645;
assign x_54936 = x_23646 & x_23647;
assign x_54937 = x_54935 & x_54936;
assign x_54938 = x_54934 & x_54937;
assign x_54939 = x_23648 & x_23649;
assign x_54940 = x_23650 & x_23651;
assign x_54941 = x_54939 & x_54940;
assign x_54942 = x_23652 & x_23653;
assign x_54943 = x_23654 & x_23655;
assign x_54944 = x_54942 & x_54943;
assign x_54945 = x_54941 & x_54944;
assign x_54946 = x_54938 & x_54945;
assign x_54947 = x_54931 & x_54946;
assign x_54948 = x_54917 & x_54947;
assign x_54949 = x_23657 & x_23658;
assign x_54950 = x_23656 & x_54949;
assign x_54951 = x_23659 & x_23660;
assign x_54952 = x_23661 & x_23662;
assign x_54953 = x_54951 & x_54952;
assign x_54954 = x_54950 & x_54953;
assign x_54955 = x_23663 & x_23664;
assign x_54956 = x_23665 & x_23666;
assign x_54957 = x_54955 & x_54956;
assign x_54958 = x_23667 & x_23668;
assign x_54959 = x_23669 & x_23670;
assign x_54960 = x_54958 & x_54959;
assign x_54961 = x_54957 & x_54960;
assign x_54962 = x_54954 & x_54961;
assign x_54963 = x_23672 & x_23673;
assign x_54964 = x_23671 & x_54963;
assign x_54965 = x_23674 & x_23675;
assign x_54966 = x_23676 & x_23677;
assign x_54967 = x_54965 & x_54966;
assign x_54968 = x_54964 & x_54967;
assign x_54969 = x_23678 & x_23679;
assign x_54970 = x_23680 & x_23681;
assign x_54971 = x_54969 & x_54970;
assign x_54972 = x_23682 & x_23683;
assign x_54973 = x_23684 & x_23685;
assign x_54974 = x_54972 & x_54973;
assign x_54975 = x_54971 & x_54974;
assign x_54976 = x_54968 & x_54975;
assign x_54977 = x_54962 & x_54976;
assign x_54978 = x_23687 & x_23688;
assign x_54979 = x_23686 & x_54978;
assign x_54980 = x_23689 & x_23690;
assign x_54981 = x_23691 & x_23692;
assign x_54982 = x_54980 & x_54981;
assign x_54983 = x_54979 & x_54982;
assign x_54984 = x_23693 & x_23694;
assign x_54985 = x_23695 & x_23696;
assign x_54986 = x_54984 & x_54985;
assign x_54987 = x_23697 & x_23698;
assign x_54988 = x_23699 & x_23700;
assign x_54989 = x_54987 & x_54988;
assign x_54990 = x_54986 & x_54989;
assign x_54991 = x_54983 & x_54990;
assign x_54992 = x_23701 & x_23702;
assign x_54993 = x_23703 & x_23704;
assign x_54994 = x_54992 & x_54993;
assign x_54995 = x_23705 & x_23706;
assign x_54996 = x_23707 & x_23708;
assign x_54997 = x_54995 & x_54996;
assign x_54998 = x_54994 & x_54997;
assign x_54999 = x_23709 & x_23710;
assign x_55000 = x_23711 & x_23712;
assign x_55001 = x_54999 & x_55000;
assign x_55002 = x_23713 & x_23714;
assign x_55003 = x_23715 & x_23716;
assign x_55004 = x_55002 & x_55003;
assign x_55005 = x_55001 & x_55004;
assign x_55006 = x_54998 & x_55005;
assign x_55007 = x_54991 & x_55006;
assign x_55008 = x_54977 & x_55007;
assign x_55009 = x_54948 & x_55008;
assign x_55010 = x_54888 & x_55009;
assign x_55011 = x_23718 & x_23719;
assign x_55012 = x_23717 & x_55011;
assign x_55013 = x_23720 & x_23721;
assign x_55014 = x_23722 & x_23723;
assign x_55015 = x_55013 & x_55014;
assign x_55016 = x_55012 & x_55015;
assign x_55017 = x_23724 & x_23725;
assign x_55018 = x_23726 & x_23727;
assign x_55019 = x_55017 & x_55018;
assign x_55020 = x_23728 & x_23729;
assign x_55021 = x_23730 & x_23731;
assign x_55022 = x_55020 & x_55021;
assign x_55023 = x_55019 & x_55022;
assign x_55024 = x_55016 & x_55023;
assign x_55025 = x_23733 & x_23734;
assign x_55026 = x_23732 & x_55025;
assign x_55027 = x_23735 & x_23736;
assign x_55028 = x_23737 & x_23738;
assign x_55029 = x_55027 & x_55028;
assign x_55030 = x_55026 & x_55029;
assign x_55031 = x_23739 & x_23740;
assign x_55032 = x_23741 & x_23742;
assign x_55033 = x_55031 & x_55032;
assign x_55034 = x_23743 & x_23744;
assign x_55035 = x_23745 & x_23746;
assign x_55036 = x_55034 & x_55035;
assign x_55037 = x_55033 & x_55036;
assign x_55038 = x_55030 & x_55037;
assign x_55039 = x_55024 & x_55038;
assign x_55040 = x_23748 & x_23749;
assign x_55041 = x_23747 & x_55040;
assign x_55042 = x_23750 & x_23751;
assign x_55043 = x_23752 & x_23753;
assign x_55044 = x_55042 & x_55043;
assign x_55045 = x_55041 & x_55044;
assign x_55046 = x_23754 & x_23755;
assign x_55047 = x_23756 & x_23757;
assign x_55048 = x_55046 & x_55047;
assign x_55049 = x_23758 & x_23759;
assign x_55050 = x_23760 & x_23761;
assign x_55051 = x_55049 & x_55050;
assign x_55052 = x_55048 & x_55051;
assign x_55053 = x_55045 & x_55052;
assign x_55054 = x_23762 & x_23763;
assign x_55055 = x_23764 & x_23765;
assign x_55056 = x_55054 & x_55055;
assign x_55057 = x_23766 & x_23767;
assign x_55058 = x_23768 & x_23769;
assign x_55059 = x_55057 & x_55058;
assign x_55060 = x_55056 & x_55059;
assign x_55061 = x_23770 & x_23771;
assign x_55062 = x_23772 & x_23773;
assign x_55063 = x_55061 & x_55062;
assign x_55064 = x_23774 & x_23775;
assign x_55065 = x_23776 & x_23777;
assign x_55066 = x_55064 & x_55065;
assign x_55067 = x_55063 & x_55066;
assign x_55068 = x_55060 & x_55067;
assign x_55069 = x_55053 & x_55068;
assign x_55070 = x_55039 & x_55069;
assign x_55071 = x_23779 & x_23780;
assign x_55072 = x_23778 & x_55071;
assign x_55073 = x_23781 & x_23782;
assign x_55074 = x_23783 & x_23784;
assign x_55075 = x_55073 & x_55074;
assign x_55076 = x_55072 & x_55075;
assign x_55077 = x_23785 & x_23786;
assign x_55078 = x_23787 & x_23788;
assign x_55079 = x_55077 & x_55078;
assign x_55080 = x_23789 & x_23790;
assign x_55081 = x_23791 & x_23792;
assign x_55082 = x_55080 & x_55081;
assign x_55083 = x_55079 & x_55082;
assign x_55084 = x_55076 & x_55083;
assign x_55085 = x_23794 & x_23795;
assign x_55086 = x_23793 & x_55085;
assign x_55087 = x_23796 & x_23797;
assign x_55088 = x_23798 & x_23799;
assign x_55089 = x_55087 & x_55088;
assign x_55090 = x_55086 & x_55089;
assign x_55091 = x_23800 & x_23801;
assign x_55092 = x_23802 & x_23803;
assign x_55093 = x_55091 & x_55092;
assign x_55094 = x_23804 & x_23805;
assign x_55095 = x_23806 & x_23807;
assign x_55096 = x_55094 & x_55095;
assign x_55097 = x_55093 & x_55096;
assign x_55098 = x_55090 & x_55097;
assign x_55099 = x_55084 & x_55098;
assign x_55100 = x_23809 & x_23810;
assign x_55101 = x_23808 & x_55100;
assign x_55102 = x_23811 & x_23812;
assign x_55103 = x_23813 & x_23814;
assign x_55104 = x_55102 & x_55103;
assign x_55105 = x_55101 & x_55104;
assign x_55106 = x_23815 & x_23816;
assign x_55107 = x_23817 & x_23818;
assign x_55108 = x_55106 & x_55107;
assign x_55109 = x_23819 & x_23820;
assign x_55110 = x_23821 & x_23822;
assign x_55111 = x_55109 & x_55110;
assign x_55112 = x_55108 & x_55111;
assign x_55113 = x_55105 & x_55112;
assign x_55114 = x_23823 & x_23824;
assign x_55115 = x_23825 & x_23826;
assign x_55116 = x_55114 & x_55115;
assign x_55117 = x_23827 & x_23828;
assign x_55118 = x_23829 & x_23830;
assign x_55119 = x_55117 & x_55118;
assign x_55120 = x_55116 & x_55119;
assign x_55121 = x_23831 & x_23832;
assign x_55122 = x_23833 & x_23834;
assign x_55123 = x_55121 & x_55122;
assign x_55124 = x_23835 & x_23836;
assign x_55125 = x_23837 & x_23838;
assign x_55126 = x_55124 & x_55125;
assign x_55127 = x_55123 & x_55126;
assign x_55128 = x_55120 & x_55127;
assign x_55129 = x_55113 & x_55128;
assign x_55130 = x_55099 & x_55129;
assign x_55131 = x_55070 & x_55130;
assign x_55132 = x_23840 & x_23841;
assign x_55133 = x_23839 & x_55132;
assign x_55134 = x_23842 & x_23843;
assign x_55135 = x_23844 & x_23845;
assign x_55136 = x_55134 & x_55135;
assign x_55137 = x_55133 & x_55136;
assign x_55138 = x_23846 & x_23847;
assign x_55139 = x_23848 & x_23849;
assign x_55140 = x_55138 & x_55139;
assign x_55141 = x_23850 & x_23851;
assign x_55142 = x_23852 & x_23853;
assign x_55143 = x_55141 & x_55142;
assign x_55144 = x_55140 & x_55143;
assign x_55145 = x_55137 & x_55144;
assign x_55146 = x_23855 & x_23856;
assign x_55147 = x_23854 & x_55146;
assign x_55148 = x_23857 & x_23858;
assign x_55149 = x_23859 & x_23860;
assign x_55150 = x_55148 & x_55149;
assign x_55151 = x_55147 & x_55150;
assign x_55152 = x_23861 & x_23862;
assign x_55153 = x_23863 & x_23864;
assign x_55154 = x_55152 & x_55153;
assign x_55155 = x_23865 & x_23866;
assign x_55156 = x_23867 & x_23868;
assign x_55157 = x_55155 & x_55156;
assign x_55158 = x_55154 & x_55157;
assign x_55159 = x_55151 & x_55158;
assign x_55160 = x_55145 & x_55159;
assign x_55161 = x_23870 & x_23871;
assign x_55162 = x_23869 & x_55161;
assign x_55163 = x_23872 & x_23873;
assign x_55164 = x_23874 & x_23875;
assign x_55165 = x_55163 & x_55164;
assign x_55166 = x_55162 & x_55165;
assign x_55167 = x_23876 & x_23877;
assign x_55168 = x_23878 & x_23879;
assign x_55169 = x_55167 & x_55168;
assign x_55170 = x_23880 & x_23881;
assign x_55171 = x_23882 & x_23883;
assign x_55172 = x_55170 & x_55171;
assign x_55173 = x_55169 & x_55172;
assign x_55174 = x_55166 & x_55173;
assign x_55175 = x_23884 & x_23885;
assign x_55176 = x_23886 & x_23887;
assign x_55177 = x_55175 & x_55176;
assign x_55178 = x_23888 & x_23889;
assign x_55179 = x_23890 & x_23891;
assign x_55180 = x_55178 & x_55179;
assign x_55181 = x_55177 & x_55180;
assign x_55182 = x_23892 & x_23893;
assign x_55183 = x_23894 & x_23895;
assign x_55184 = x_55182 & x_55183;
assign x_55185 = x_23896 & x_23897;
assign x_55186 = x_23898 & x_23899;
assign x_55187 = x_55185 & x_55186;
assign x_55188 = x_55184 & x_55187;
assign x_55189 = x_55181 & x_55188;
assign x_55190 = x_55174 & x_55189;
assign x_55191 = x_55160 & x_55190;
assign x_55192 = x_23901 & x_23902;
assign x_55193 = x_23900 & x_55192;
assign x_55194 = x_23903 & x_23904;
assign x_55195 = x_23905 & x_23906;
assign x_55196 = x_55194 & x_55195;
assign x_55197 = x_55193 & x_55196;
assign x_55198 = x_23907 & x_23908;
assign x_55199 = x_23909 & x_23910;
assign x_55200 = x_55198 & x_55199;
assign x_55201 = x_23911 & x_23912;
assign x_55202 = x_23913 & x_23914;
assign x_55203 = x_55201 & x_55202;
assign x_55204 = x_55200 & x_55203;
assign x_55205 = x_55197 & x_55204;
assign x_55206 = x_23915 & x_23916;
assign x_55207 = x_23917 & x_23918;
assign x_55208 = x_55206 & x_55207;
assign x_55209 = x_23919 & x_23920;
assign x_55210 = x_23921 & x_23922;
assign x_55211 = x_55209 & x_55210;
assign x_55212 = x_55208 & x_55211;
assign x_55213 = x_23923 & x_23924;
assign x_55214 = x_23925 & x_23926;
assign x_55215 = x_55213 & x_55214;
assign x_55216 = x_23927 & x_23928;
assign x_55217 = x_23929 & x_23930;
assign x_55218 = x_55216 & x_55217;
assign x_55219 = x_55215 & x_55218;
assign x_55220 = x_55212 & x_55219;
assign x_55221 = x_55205 & x_55220;
assign x_55222 = x_23932 & x_23933;
assign x_55223 = x_23931 & x_55222;
assign x_55224 = x_23934 & x_23935;
assign x_55225 = x_23936 & x_23937;
assign x_55226 = x_55224 & x_55225;
assign x_55227 = x_55223 & x_55226;
assign x_55228 = x_23938 & x_23939;
assign x_55229 = x_23940 & x_23941;
assign x_55230 = x_55228 & x_55229;
assign x_55231 = x_23942 & x_23943;
assign x_55232 = x_23944 & x_23945;
assign x_55233 = x_55231 & x_55232;
assign x_55234 = x_55230 & x_55233;
assign x_55235 = x_55227 & x_55234;
assign x_55236 = x_23946 & x_23947;
assign x_55237 = x_23948 & x_23949;
assign x_55238 = x_55236 & x_55237;
assign x_55239 = x_23950 & x_23951;
assign x_55240 = x_23952 & x_23953;
assign x_55241 = x_55239 & x_55240;
assign x_55242 = x_55238 & x_55241;
assign x_55243 = x_23954 & x_23955;
assign x_55244 = x_23956 & x_23957;
assign x_55245 = x_55243 & x_55244;
assign x_55246 = x_23958 & x_23959;
assign x_55247 = x_23960 & x_23961;
assign x_55248 = x_55246 & x_55247;
assign x_55249 = x_55245 & x_55248;
assign x_55250 = x_55242 & x_55249;
assign x_55251 = x_55235 & x_55250;
assign x_55252 = x_55221 & x_55251;
assign x_55253 = x_55191 & x_55252;
assign x_55254 = x_55131 & x_55253;
assign x_55255 = x_55010 & x_55254;
assign x_55256 = x_23963 & x_23964;
assign x_55257 = x_23962 & x_55256;
assign x_55258 = x_23965 & x_23966;
assign x_55259 = x_23967 & x_23968;
assign x_55260 = x_55258 & x_55259;
assign x_55261 = x_55257 & x_55260;
assign x_55262 = x_23969 & x_23970;
assign x_55263 = x_23971 & x_23972;
assign x_55264 = x_55262 & x_55263;
assign x_55265 = x_23973 & x_23974;
assign x_55266 = x_23975 & x_23976;
assign x_55267 = x_55265 & x_55266;
assign x_55268 = x_55264 & x_55267;
assign x_55269 = x_55261 & x_55268;
assign x_55270 = x_23978 & x_23979;
assign x_55271 = x_23977 & x_55270;
assign x_55272 = x_23980 & x_23981;
assign x_55273 = x_23982 & x_23983;
assign x_55274 = x_55272 & x_55273;
assign x_55275 = x_55271 & x_55274;
assign x_55276 = x_23984 & x_23985;
assign x_55277 = x_23986 & x_23987;
assign x_55278 = x_55276 & x_55277;
assign x_55279 = x_23988 & x_23989;
assign x_55280 = x_23990 & x_23991;
assign x_55281 = x_55279 & x_55280;
assign x_55282 = x_55278 & x_55281;
assign x_55283 = x_55275 & x_55282;
assign x_55284 = x_55269 & x_55283;
assign x_55285 = x_23993 & x_23994;
assign x_55286 = x_23992 & x_55285;
assign x_55287 = x_23995 & x_23996;
assign x_55288 = x_23997 & x_23998;
assign x_55289 = x_55287 & x_55288;
assign x_55290 = x_55286 & x_55289;
assign x_55291 = x_23999 & x_24000;
assign x_55292 = x_24001 & x_24002;
assign x_55293 = x_55291 & x_55292;
assign x_55294 = x_24003 & x_24004;
assign x_55295 = x_24005 & x_24006;
assign x_55296 = x_55294 & x_55295;
assign x_55297 = x_55293 & x_55296;
assign x_55298 = x_55290 & x_55297;
assign x_55299 = x_24007 & x_24008;
assign x_55300 = x_24009 & x_24010;
assign x_55301 = x_55299 & x_55300;
assign x_55302 = x_24011 & x_24012;
assign x_55303 = x_24013 & x_24014;
assign x_55304 = x_55302 & x_55303;
assign x_55305 = x_55301 & x_55304;
assign x_55306 = x_24015 & x_24016;
assign x_55307 = x_24017 & x_24018;
assign x_55308 = x_55306 & x_55307;
assign x_55309 = x_24019 & x_24020;
assign x_55310 = x_24021 & x_24022;
assign x_55311 = x_55309 & x_55310;
assign x_55312 = x_55308 & x_55311;
assign x_55313 = x_55305 & x_55312;
assign x_55314 = x_55298 & x_55313;
assign x_55315 = x_55284 & x_55314;
assign x_55316 = x_24024 & x_24025;
assign x_55317 = x_24023 & x_55316;
assign x_55318 = x_24026 & x_24027;
assign x_55319 = x_24028 & x_24029;
assign x_55320 = x_55318 & x_55319;
assign x_55321 = x_55317 & x_55320;
assign x_55322 = x_24030 & x_24031;
assign x_55323 = x_24032 & x_24033;
assign x_55324 = x_55322 & x_55323;
assign x_55325 = x_24034 & x_24035;
assign x_55326 = x_24036 & x_24037;
assign x_55327 = x_55325 & x_55326;
assign x_55328 = x_55324 & x_55327;
assign x_55329 = x_55321 & x_55328;
assign x_55330 = x_24039 & x_24040;
assign x_55331 = x_24038 & x_55330;
assign x_55332 = x_24041 & x_24042;
assign x_55333 = x_24043 & x_24044;
assign x_55334 = x_55332 & x_55333;
assign x_55335 = x_55331 & x_55334;
assign x_55336 = x_24045 & x_24046;
assign x_55337 = x_24047 & x_24048;
assign x_55338 = x_55336 & x_55337;
assign x_55339 = x_24049 & x_24050;
assign x_55340 = x_24051 & x_24052;
assign x_55341 = x_55339 & x_55340;
assign x_55342 = x_55338 & x_55341;
assign x_55343 = x_55335 & x_55342;
assign x_55344 = x_55329 & x_55343;
assign x_55345 = x_24054 & x_24055;
assign x_55346 = x_24053 & x_55345;
assign x_55347 = x_24056 & x_24057;
assign x_55348 = x_24058 & x_24059;
assign x_55349 = x_55347 & x_55348;
assign x_55350 = x_55346 & x_55349;
assign x_55351 = x_24060 & x_24061;
assign x_55352 = x_24062 & x_24063;
assign x_55353 = x_55351 & x_55352;
assign x_55354 = x_24064 & x_24065;
assign x_55355 = x_24066 & x_24067;
assign x_55356 = x_55354 & x_55355;
assign x_55357 = x_55353 & x_55356;
assign x_55358 = x_55350 & x_55357;
assign x_55359 = x_24068 & x_24069;
assign x_55360 = x_24070 & x_24071;
assign x_55361 = x_55359 & x_55360;
assign x_55362 = x_24072 & x_24073;
assign x_55363 = x_24074 & x_24075;
assign x_55364 = x_55362 & x_55363;
assign x_55365 = x_55361 & x_55364;
assign x_55366 = x_24076 & x_24077;
assign x_55367 = x_24078 & x_24079;
assign x_55368 = x_55366 & x_55367;
assign x_55369 = x_24080 & x_24081;
assign x_55370 = x_24082 & x_24083;
assign x_55371 = x_55369 & x_55370;
assign x_55372 = x_55368 & x_55371;
assign x_55373 = x_55365 & x_55372;
assign x_55374 = x_55358 & x_55373;
assign x_55375 = x_55344 & x_55374;
assign x_55376 = x_55315 & x_55375;
assign x_55377 = x_24085 & x_24086;
assign x_55378 = x_24084 & x_55377;
assign x_55379 = x_24087 & x_24088;
assign x_55380 = x_24089 & x_24090;
assign x_55381 = x_55379 & x_55380;
assign x_55382 = x_55378 & x_55381;
assign x_55383 = x_24091 & x_24092;
assign x_55384 = x_24093 & x_24094;
assign x_55385 = x_55383 & x_55384;
assign x_55386 = x_24095 & x_24096;
assign x_55387 = x_24097 & x_24098;
assign x_55388 = x_55386 & x_55387;
assign x_55389 = x_55385 & x_55388;
assign x_55390 = x_55382 & x_55389;
assign x_55391 = x_24100 & x_24101;
assign x_55392 = x_24099 & x_55391;
assign x_55393 = x_24102 & x_24103;
assign x_55394 = x_24104 & x_24105;
assign x_55395 = x_55393 & x_55394;
assign x_55396 = x_55392 & x_55395;
assign x_55397 = x_24106 & x_24107;
assign x_55398 = x_24108 & x_24109;
assign x_55399 = x_55397 & x_55398;
assign x_55400 = x_24110 & x_24111;
assign x_55401 = x_24112 & x_24113;
assign x_55402 = x_55400 & x_55401;
assign x_55403 = x_55399 & x_55402;
assign x_55404 = x_55396 & x_55403;
assign x_55405 = x_55390 & x_55404;
assign x_55406 = x_24115 & x_24116;
assign x_55407 = x_24114 & x_55406;
assign x_55408 = x_24117 & x_24118;
assign x_55409 = x_24119 & x_24120;
assign x_55410 = x_55408 & x_55409;
assign x_55411 = x_55407 & x_55410;
assign x_55412 = x_24121 & x_24122;
assign x_55413 = x_24123 & x_24124;
assign x_55414 = x_55412 & x_55413;
assign x_55415 = x_24125 & x_24126;
assign x_55416 = x_24127 & x_24128;
assign x_55417 = x_55415 & x_55416;
assign x_55418 = x_55414 & x_55417;
assign x_55419 = x_55411 & x_55418;
assign x_55420 = x_24129 & x_24130;
assign x_55421 = x_24131 & x_24132;
assign x_55422 = x_55420 & x_55421;
assign x_55423 = x_24133 & x_24134;
assign x_55424 = x_24135 & x_24136;
assign x_55425 = x_55423 & x_55424;
assign x_55426 = x_55422 & x_55425;
assign x_55427 = x_24137 & x_24138;
assign x_55428 = x_24139 & x_24140;
assign x_55429 = x_55427 & x_55428;
assign x_55430 = x_24141 & x_24142;
assign x_55431 = x_24143 & x_24144;
assign x_55432 = x_55430 & x_55431;
assign x_55433 = x_55429 & x_55432;
assign x_55434 = x_55426 & x_55433;
assign x_55435 = x_55419 & x_55434;
assign x_55436 = x_55405 & x_55435;
assign x_55437 = x_24146 & x_24147;
assign x_55438 = x_24145 & x_55437;
assign x_55439 = x_24148 & x_24149;
assign x_55440 = x_24150 & x_24151;
assign x_55441 = x_55439 & x_55440;
assign x_55442 = x_55438 & x_55441;
assign x_55443 = x_24152 & x_24153;
assign x_55444 = x_24154 & x_24155;
assign x_55445 = x_55443 & x_55444;
assign x_55446 = x_24156 & x_24157;
assign x_55447 = x_24158 & x_24159;
assign x_55448 = x_55446 & x_55447;
assign x_55449 = x_55445 & x_55448;
assign x_55450 = x_55442 & x_55449;
assign x_55451 = x_24161 & x_24162;
assign x_55452 = x_24160 & x_55451;
assign x_55453 = x_24163 & x_24164;
assign x_55454 = x_24165 & x_24166;
assign x_55455 = x_55453 & x_55454;
assign x_55456 = x_55452 & x_55455;
assign x_55457 = x_24167 & x_24168;
assign x_55458 = x_24169 & x_24170;
assign x_55459 = x_55457 & x_55458;
assign x_55460 = x_24171 & x_24172;
assign x_55461 = x_24173 & x_24174;
assign x_55462 = x_55460 & x_55461;
assign x_55463 = x_55459 & x_55462;
assign x_55464 = x_55456 & x_55463;
assign x_55465 = x_55450 & x_55464;
assign x_55466 = x_24176 & x_24177;
assign x_55467 = x_24175 & x_55466;
assign x_55468 = x_24178 & x_24179;
assign x_55469 = x_24180 & x_24181;
assign x_55470 = x_55468 & x_55469;
assign x_55471 = x_55467 & x_55470;
assign x_55472 = x_24182 & x_24183;
assign x_55473 = x_24184 & x_24185;
assign x_55474 = x_55472 & x_55473;
assign x_55475 = x_24186 & x_24187;
assign x_55476 = x_24188 & x_24189;
assign x_55477 = x_55475 & x_55476;
assign x_55478 = x_55474 & x_55477;
assign x_55479 = x_55471 & x_55478;
assign x_55480 = x_24190 & x_24191;
assign x_55481 = x_24192 & x_24193;
assign x_55482 = x_55480 & x_55481;
assign x_55483 = x_24194 & x_24195;
assign x_55484 = x_24196 & x_24197;
assign x_55485 = x_55483 & x_55484;
assign x_55486 = x_55482 & x_55485;
assign x_55487 = x_24198 & x_24199;
assign x_55488 = x_24200 & x_24201;
assign x_55489 = x_55487 & x_55488;
assign x_55490 = x_24202 & x_24203;
assign x_55491 = x_24204 & x_24205;
assign x_55492 = x_55490 & x_55491;
assign x_55493 = x_55489 & x_55492;
assign x_55494 = x_55486 & x_55493;
assign x_55495 = x_55479 & x_55494;
assign x_55496 = x_55465 & x_55495;
assign x_55497 = x_55436 & x_55496;
assign x_55498 = x_55376 & x_55497;
assign x_55499 = x_24207 & x_24208;
assign x_55500 = x_24206 & x_55499;
assign x_55501 = x_24209 & x_24210;
assign x_55502 = x_24211 & x_24212;
assign x_55503 = x_55501 & x_55502;
assign x_55504 = x_55500 & x_55503;
assign x_55505 = x_24213 & x_24214;
assign x_55506 = x_24215 & x_24216;
assign x_55507 = x_55505 & x_55506;
assign x_55508 = x_24217 & x_24218;
assign x_55509 = x_24219 & x_24220;
assign x_55510 = x_55508 & x_55509;
assign x_55511 = x_55507 & x_55510;
assign x_55512 = x_55504 & x_55511;
assign x_55513 = x_24222 & x_24223;
assign x_55514 = x_24221 & x_55513;
assign x_55515 = x_24224 & x_24225;
assign x_55516 = x_24226 & x_24227;
assign x_55517 = x_55515 & x_55516;
assign x_55518 = x_55514 & x_55517;
assign x_55519 = x_24228 & x_24229;
assign x_55520 = x_24230 & x_24231;
assign x_55521 = x_55519 & x_55520;
assign x_55522 = x_24232 & x_24233;
assign x_55523 = x_24234 & x_24235;
assign x_55524 = x_55522 & x_55523;
assign x_55525 = x_55521 & x_55524;
assign x_55526 = x_55518 & x_55525;
assign x_55527 = x_55512 & x_55526;
assign x_55528 = x_24237 & x_24238;
assign x_55529 = x_24236 & x_55528;
assign x_55530 = x_24239 & x_24240;
assign x_55531 = x_24241 & x_24242;
assign x_55532 = x_55530 & x_55531;
assign x_55533 = x_55529 & x_55532;
assign x_55534 = x_24243 & x_24244;
assign x_55535 = x_24245 & x_24246;
assign x_55536 = x_55534 & x_55535;
assign x_55537 = x_24247 & x_24248;
assign x_55538 = x_24249 & x_24250;
assign x_55539 = x_55537 & x_55538;
assign x_55540 = x_55536 & x_55539;
assign x_55541 = x_55533 & x_55540;
assign x_55542 = x_24251 & x_24252;
assign x_55543 = x_24253 & x_24254;
assign x_55544 = x_55542 & x_55543;
assign x_55545 = x_24255 & x_24256;
assign x_55546 = x_24257 & x_24258;
assign x_55547 = x_55545 & x_55546;
assign x_55548 = x_55544 & x_55547;
assign x_55549 = x_24259 & x_24260;
assign x_55550 = x_24261 & x_24262;
assign x_55551 = x_55549 & x_55550;
assign x_55552 = x_24263 & x_24264;
assign x_55553 = x_24265 & x_24266;
assign x_55554 = x_55552 & x_55553;
assign x_55555 = x_55551 & x_55554;
assign x_55556 = x_55548 & x_55555;
assign x_55557 = x_55541 & x_55556;
assign x_55558 = x_55527 & x_55557;
assign x_55559 = x_24268 & x_24269;
assign x_55560 = x_24267 & x_55559;
assign x_55561 = x_24270 & x_24271;
assign x_55562 = x_24272 & x_24273;
assign x_55563 = x_55561 & x_55562;
assign x_55564 = x_55560 & x_55563;
assign x_55565 = x_24274 & x_24275;
assign x_55566 = x_24276 & x_24277;
assign x_55567 = x_55565 & x_55566;
assign x_55568 = x_24278 & x_24279;
assign x_55569 = x_24280 & x_24281;
assign x_55570 = x_55568 & x_55569;
assign x_55571 = x_55567 & x_55570;
assign x_55572 = x_55564 & x_55571;
assign x_55573 = x_24283 & x_24284;
assign x_55574 = x_24282 & x_55573;
assign x_55575 = x_24285 & x_24286;
assign x_55576 = x_24287 & x_24288;
assign x_55577 = x_55575 & x_55576;
assign x_55578 = x_55574 & x_55577;
assign x_55579 = x_24289 & x_24290;
assign x_55580 = x_24291 & x_24292;
assign x_55581 = x_55579 & x_55580;
assign x_55582 = x_24293 & x_24294;
assign x_55583 = x_24295 & x_24296;
assign x_55584 = x_55582 & x_55583;
assign x_55585 = x_55581 & x_55584;
assign x_55586 = x_55578 & x_55585;
assign x_55587 = x_55572 & x_55586;
assign x_55588 = x_24298 & x_24299;
assign x_55589 = x_24297 & x_55588;
assign x_55590 = x_24300 & x_24301;
assign x_55591 = x_24302 & x_24303;
assign x_55592 = x_55590 & x_55591;
assign x_55593 = x_55589 & x_55592;
assign x_55594 = x_24304 & x_24305;
assign x_55595 = x_24306 & x_24307;
assign x_55596 = x_55594 & x_55595;
assign x_55597 = x_24308 & x_24309;
assign x_55598 = x_24310 & x_24311;
assign x_55599 = x_55597 & x_55598;
assign x_55600 = x_55596 & x_55599;
assign x_55601 = x_55593 & x_55600;
assign x_55602 = x_24312 & x_24313;
assign x_55603 = x_24314 & x_24315;
assign x_55604 = x_55602 & x_55603;
assign x_55605 = x_24316 & x_24317;
assign x_55606 = x_24318 & x_24319;
assign x_55607 = x_55605 & x_55606;
assign x_55608 = x_55604 & x_55607;
assign x_55609 = x_24320 & x_24321;
assign x_55610 = x_24322 & x_24323;
assign x_55611 = x_55609 & x_55610;
assign x_55612 = x_24324 & x_24325;
assign x_55613 = x_24326 & x_24327;
assign x_55614 = x_55612 & x_55613;
assign x_55615 = x_55611 & x_55614;
assign x_55616 = x_55608 & x_55615;
assign x_55617 = x_55601 & x_55616;
assign x_55618 = x_55587 & x_55617;
assign x_55619 = x_55558 & x_55618;
assign x_55620 = x_24329 & x_24330;
assign x_55621 = x_24328 & x_55620;
assign x_55622 = x_24331 & x_24332;
assign x_55623 = x_24333 & x_24334;
assign x_55624 = x_55622 & x_55623;
assign x_55625 = x_55621 & x_55624;
assign x_55626 = x_24335 & x_24336;
assign x_55627 = x_24337 & x_24338;
assign x_55628 = x_55626 & x_55627;
assign x_55629 = x_24339 & x_24340;
assign x_55630 = x_24341 & x_24342;
assign x_55631 = x_55629 & x_55630;
assign x_55632 = x_55628 & x_55631;
assign x_55633 = x_55625 & x_55632;
assign x_55634 = x_24344 & x_24345;
assign x_55635 = x_24343 & x_55634;
assign x_55636 = x_24346 & x_24347;
assign x_55637 = x_24348 & x_24349;
assign x_55638 = x_55636 & x_55637;
assign x_55639 = x_55635 & x_55638;
assign x_55640 = x_24350 & x_24351;
assign x_55641 = x_24352 & x_24353;
assign x_55642 = x_55640 & x_55641;
assign x_55643 = x_24354 & x_24355;
assign x_55644 = x_24356 & x_24357;
assign x_55645 = x_55643 & x_55644;
assign x_55646 = x_55642 & x_55645;
assign x_55647 = x_55639 & x_55646;
assign x_55648 = x_55633 & x_55647;
assign x_55649 = x_24359 & x_24360;
assign x_55650 = x_24358 & x_55649;
assign x_55651 = x_24361 & x_24362;
assign x_55652 = x_24363 & x_24364;
assign x_55653 = x_55651 & x_55652;
assign x_55654 = x_55650 & x_55653;
assign x_55655 = x_24365 & x_24366;
assign x_55656 = x_24367 & x_24368;
assign x_55657 = x_55655 & x_55656;
assign x_55658 = x_24369 & x_24370;
assign x_55659 = x_24371 & x_24372;
assign x_55660 = x_55658 & x_55659;
assign x_55661 = x_55657 & x_55660;
assign x_55662 = x_55654 & x_55661;
assign x_55663 = x_24373 & x_24374;
assign x_55664 = x_24375 & x_24376;
assign x_55665 = x_55663 & x_55664;
assign x_55666 = x_24377 & x_24378;
assign x_55667 = x_24379 & x_24380;
assign x_55668 = x_55666 & x_55667;
assign x_55669 = x_55665 & x_55668;
assign x_55670 = x_24381 & x_24382;
assign x_55671 = x_24383 & x_24384;
assign x_55672 = x_55670 & x_55671;
assign x_55673 = x_24385 & x_24386;
assign x_55674 = x_24387 & x_24388;
assign x_55675 = x_55673 & x_55674;
assign x_55676 = x_55672 & x_55675;
assign x_55677 = x_55669 & x_55676;
assign x_55678 = x_55662 & x_55677;
assign x_55679 = x_55648 & x_55678;
assign x_55680 = x_24390 & x_24391;
assign x_55681 = x_24389 & x_55680;
assign x_55682 = x_24392 & x_24393;
assign x_55683 = x_24394 & x_24395;
assign x_55684 = x_55682 & x_55683;
assign x_55685 = x_55681 & x_55684;
assign x_55686 = x_24396 & x_24397;
assign x_55687 = x_24398 & x_24399;
assign x_55688 = x_55686 & x_55687;
assign x_55689 = x_24400 & x_24401;
assign x_55690 = x_24402 & x_24403;
assign x_55691 = x_55689 & x_55690;
assign x_55692 = x_55688 & x_55691;
assign x_55693 = x_55685 & x_55692;
assign x_55694 = x_24404 & x_24405;
assign x_55695 = x_24406 & x_24407;
assign x_55696 = x_55694 & x_55695;
assign x_55697 = x_24408 & x_24409;
assign x_55698 = x_24410 & x_24411;
assign x_55699 = x_55697 & x_55698;
assign x_55700 = x_55696 & x_55699;
assign x_55701 = x_24412 & x_24413;
assign x_55702 = x_24414 & x_24415;
assign x_55703 = x_55701 & x_55702;
assign x_55704 = x_24416 & x_24417;
assign x_55705 = x_24418 & x_24419;
assign x_55706 = x_55704 & x_55705;
assign x_55707 = x_55703 & x_55706;
assign x_55708 = x_55700 & x_55707;
assign x_55709 = x_55693 & x_55708;
assign x_55710 = x_24421 & x_24422;
assign x_55711 = x_24420 & x_55710;
assign x_55712 = x_24423 & x_24424;
assign x_55713 = x_24425 & x_24426;
assign x_55714 = x_55712 & x_55713;
assign x_55715 = x_55711 & x_55714;
assign x_55716 = x_24427 & x_24428;
assign x_55717 = x_24429 & x_24430;
assign x_55718 = x_55716 & x_55717;
assign x_55719 = x_24431 & x_24432;
assign x_55720 = x_24433 & x_24434;
assign x_55721 = x_55719 & x_55720;
assign x_55722 = x_55718 & x_55721;
assign x_55723 = x_55715 & x_55722;
assign x_55724 = x_24435 & x_24436;
assign x_55725 = x_24437 & x_24438;
assign x_55726 = x_55724 & x_55725;
assign x_55727 = x_24439 & x_24440;
assign x_55728 = x_24441 & x_24442;
assign x_55729 = x_55727 & x_55728;
assign x_55730 = x_55726 & x_55729;
assign x_55731 = x_24443 & x_24444;
assign x_55732 = x_24445 & x_24446;
assign x_55733 = x_55731 & x_55732;
assign x_55734 = x_24447 & x_24448;
assign x_55735 = x_24449 & x_24450;
assign x_55736 = x_55734 & x_55735;
assign x_55737 = x_55733 & x_55736;
assign x_55738 = x_55730 & x_55737;
assign x_55739 = x_55723 & x_55738;
assign x_55740 = x_55709 & x_55739;
assign x_55741 = x_55679 & x_55740;
assign x_55742 = x_55619 & x_55741;
assign x_55743 = x_55498 & x_55742;
assign x_55744 = x_55255 & x_55743;
assign x_55745 = x_24452 & x_24453;
assign x_55746 = x_24451 & x_55745;
assign x_55747 = x_24454 & x_24455;
assign x_55748 = x_24456 & x_24457;
assign x_55749 = x_55747 & x_55748;
assign x_55750 = x_55746 & x_55749;
assign x_55751 = x_24458 & x_24459;
assign x_55752 = x_24460 & x_24461;
assign x_55753 = x_55751 & x_55752;
assign x_55754 = x_24462 & x_24463;
assign x_55755 = x_24464 & x_24465;
assign x_55756 = x_55754 & x_55755;
assign x_55757 = x_55753 & x_55756;
assign x_55758 = x_55750 & x_55757;
assign x_55759 = x_24467 & x_24468;
assign x_55760 = x_24466 & x_55759;
assign x_55761 = x_24469 & x_24470;
assign x_55762 = x_24471 & x_24472;
assign x_55763 = x_55761 & x_55762;
assign x_55764 = x_55760 & x_55763;
assign x_55765 = x_24473 & x_24474;
assign x_55766 = x_24475 & x_24476;
assign x_55767 = x_55765 & x_55766;
assign x_55768 = x_24477 & x_24478;
assign x_55769 = x_24479 & x_24480;
assign x_55770 = x_55768 & x_55769;
assign x_55771 = x_55767 & x_55770;
assign x_55772 = x_55764 & x_55771;
assign x_55773 = x_55758 & x_55772;
assign x_55774 = x_24482 & x_24483;
assign x_55775 = x_24481 & x_55774;
assign x_55776 = x_24484 & x_24485;
assign x_55777 = x_24486 & x_24487;
assign x_55778 = x_55776 & x_55777;
assign x_55779 = x_55775 & x_55778;
assign x_55780 = x_24488 & x_24489;
assign x_55781 = x_24490 & x_24491;
assign x_55782 = x_55780 & x_55781;
assign x_55783 = x_24492 & x_24493;
assign x_55784 = x_24494 & x_24495;
assign x_55785 = x_55783 & x_55784;
assign x_55786 = x_55782 & x_55785;
assign x_55787 = x_55779 & x_55786;
assign x_55788 = x_24496 & x_24497;
assign x_55789 = x_24498 & x_24499;
assign x_55790 = x_55788 & x_55789;
assign x_55791 = x_24500 & x_24501;
assign x_55792 = x_24502 & x_24503;
assign x_55793 = x_55791 & x_55792;
assign x_55794 = x_55790 & x_55793;
assign x_55795 = x_24504 & x_24505;
assign x_55796 = x_24506 & x_24507;
assign x_55797 = x_55795 & x_55796;
assign x_55798 = x_24508 & x_24509;
assign x_55799 = x_24510 & x_24511;
assign x_55800 = x_55798 & x_55799;
assign x_55801 = x_55797 & x_55800;
assign x_55802 = x_55794 & x_55801;
assign x_55803 = x_55787 & x_55802;
assign x_55804 = x_55773 & x_55803;
assign x_55805 = x_24513 & x_24514;
assign x_55806 = x_24512 & x_55805;
assign x_55807 = x_24515 & x_24516;
assign x_55808 = x_24517 & x_24518;
assign x_55809 = x_55807 & x_55808;
assign x_55810 = x_55806 & x_55809;
assign x_55811 = x_24519 & x_24520;
assign x_55812 = x_24521 & x_24522;
assign x_55813 = x_55811 & x_55812;
assign x_55814 = x_24523 & x_24524;
assign x_55815 = x_24525 & x_24526;
assign x_55816 = x_55814 & x_55815;
assign x_55817 = x_55813 & x_55816;
assign x_55818 = x_55810 & x_55817;
assign x_55819 = x_24528 & x_24529;
assign x_55820 = x_24527 & x_55819;
assign x_55821 = x_24530 & x_24531;
assign x_55822 = x_24532 & x_24533;
assign x_55823 = x_55821 & x_55822;
assign x_55824 = x_55820 & x_55823;
assign x_55825 = x_24534 & x_24535;
assign x_55826 = x_24536 & x_24537;
assign x_55827 = x_55825 & x_55826;
assign x_55828 = x_24538 & x_24539;
assign x_55829 = x_24540 & x_24541;
assign x_55830 = x_55828 & x_55829;
assign x_55831 = x_55827 & x_55830;
assign x_55832 = x_55824 & x_55831;
assign x_55833 = x_55818 & x_55832;
assign x_55834 = x_24543 & x_24544;
assign x_55835 = x_24542 & x_55834;
assign x_55836 = x_24545 & x_24546;
assign x_55837 = x_24547 & x_24548;
assign x_55838 = x_55836 & x_55837;
assign x_55839 = x_55835 & x_55838;
assign x_55840 = x_24549 & x_24550;
assign x_55841 = x_24551 & x_24552;
assign x_55842 = x_55840 & x_55841;
assign x_55843 = x_24553 & x_24554;
assign x_55844 = x_24555 & x_24556;
assign x_55845 = x_55843 & x_55844;
assign x_55846 = x_55842 & x_55845;
assign x_55847 = x_55839 & x_55846;
assign x_55848 = x_24557 & x_24558;
assign x_55849 = x_24559 & x_24560;
assign x_55850 = x_55848 & x_55849;
assign x_55851 = x_24561 & x_24562;
assign x_55852 = x_24563 & x_24564;
assign x_55853 = x_55851 & x_55852;
assign x_55854 = x_55850 & x_55853;
assign x_55855 = x_24565 & x_24566;
assign x_55856 = x_24567 & x_24568;
assign x_55857 = x_55855 & x_55856;
assign x_55858 = x_24569 & x_24570;
assign x_55859 = x_24571 & x_24572;
assign x_55860 = x_55858 & x_55859;
assign x_55861 = x_55857 & x_55860;
assign x_55862 = x_55854 & x_55861;
assign x_55863 = x_55847 & x_55862;
assign x_55864 = x_55833 & x_55863;
assign x_55865 = x_55804 & x_55864;
assign x_55866 = x_24574 & x_24575;
assign x_55867 = x_24573 & x_55866;
assign x_55868 = x_24576 & x_24577;
assign x_55869 = x_24578 & x_24579;
assign x_55870 = x_55868 & x_55869;
assign x_55871 = x_55867 & x_55870;
assign x_55872 = x_24580 & x_24581;
assign x_55873 = x_24582 & x_24583;
assign x_55874 = x_55872 & x_55873;
assign x_55875 = x_24584 & x_24585;
assign x_55876 = x_24586 & x_24587;
assign x_55877 = x_55875 & x_55876;
assign x_55878 = x_55874 & x_55877;
assign x_55879 = x_55871 & x_55878;
assign x_55880 = x_24589 & x_24590;
assign x_55881 = x_24588 & x_55880;
assign x_55882 = x_24591 & x_24592;
assign x_55883 = x_24593 & x_24594;
assign x_55884 = x_55882 & x_55883;
assign x_55885 = x_55881 & x_55884;
assign x_55886 = x_24595 & x_24596;
assign x_55887 = x_24597 & x_24598;
assign x_55888 = x_55886 & x_55887;
assign x_55889 = x_24599 & x_24600;
assign x_55890 = x_24601 & x_24602;
assign x_55891 = x_55889 & x_55890;
assign x_55892 = x_55888 & x_55891;
assign x_55893 = x_55885 & x_55892;
assign x_55894 = x_55879 & x_55893;
assign x_55895 = x_24604 & x_24605;
assign x_55896 = x_24603 & x_55895;
assign x_55897 = x_24606 & x_24607;
assign x_55898 = x_24608 & x_24609;
assign x_55899 = x_55897 & x_55898;
assign x_55900 = x_55896 & x_55899;
assign x_55901 = x_24610 & x_24611;
assign x_55902 = x_24612 & x_24613;
assign x_55903 = x_55901 & x_55902;
assign x_55904 = x_24614 & x_24615;
assign x_55905 = x_24616 & x_24617;
assign x_55906 = x_55904 & x_55905;
assign x_55907 = x_55903 & x_55906;
assign x_55908 = x_55900 & x_55907;
assign x_55909 = x_24618 & x_24619;
assign x_55910 = x_24620 & x_24621;
assign x_55911 = x_55909 & x_55910;
assign x_55912 = x_24622 & x_24623;
assign x_55913 = x_24624 & x_24625;
assign x_55914 = x_55912 & x_55913;
assign x_55915 = x_55911 & x_55914;
assign x_55916 = x_24626 & x_24627;
assign x_55917 = x_24628 & x_24629;
assign x_55918 = x_55916 & x_55917;
assign x_55919 = x_24630 & x_24631;
assign x_55920 = x_24632 & x_24633;
assign x_55921 = x_55919 & x_55920;
assign x_55922 = x_55918 & x_55921;
assign x_55923 = x_55915 & x_55922;
assign x_55924 = x_55908 & x_55923;
assign x_55925 = x_55894 & x_55924;
assign x_55926 = x_24635 & x_24636;
assign x_55927 = x_24634 & x_55926;
assign x_55928 = x_24637 & x_24638;
assign x_55929 = x_24639 & x_24640;
assign x_55930 = x_55928 & x_55929;
assign x_55931 = x_55927 & x_55930;
assign x_55932 = x_24641 & x_24642;
assign x_55933 = x_24643 & x_24644;
assign x_55934 = x_55932 & x_55933;
assign x_55935 = x_24645 & x_24646;
assign x_55936 = x_24647 & x_24648;
assign x_55937 = x_55935 & x_55936;
assign x_55938 = x_55934 & x_55937;
assign x_55939 = x_55931 & x_55938;
assign x_55940 = x_24650 & x_24651;
assign x_55941 = x_24649 & x_55940;
assign x_55942 = x_24652 & x_24653;
assign x_55943 = x_24654 & x_24655;
assign x_55944 = x_55942 & x_55943;
assign x_55945 = x_55941 & x_55944;
assign x_55946 = x_24656 & x_24657;
assign x_55947 = x_24658 & x_24659;
assign x_55948 = x_55946 & x_55947;
assign x_55949 = x_24660 & x_24661;
assign x_55950 = x_24662 & x_24663;
assign x_55951 = x_55949 & x_55950;
assign x_55952 = x_55948 & x_55951;
assign x_55953 = x_55945 & x_55952;
assign x_55954 = x_55939 & x_55953;
assign x_55955 = x_24665 & x_24666;
assign x_55956 = x_24664 & x_55955;
assign x_55957 = x_24667 & x_24668;
assign x_55958 = x_24669 & x_24670;
assign x_55959 = x_55957 & x_55958;
assign x_55960 = x_55956 & x_55959;
assign x_55961 = x_24671 & x_24672;
assign x_55962 = x_24673 & x_24674;
assign x_55963 = x_55961 & x_55962;
assign x_55964 = x_24675 & x_24676;
assign x_55965 = x_24677 & x_24678;
assign x_55966 = x_55964 & x_55965;
assign x_55967 = x_55963 & x_55966;
assign x_55968 = x_55960 & x_55967;
assign x_55969 = x_24679 & x_24680;
assign x_55970 = x_24681 & x_24682;
assign x_55971 = x_55969 & x_55970;
assign x_55972 = x_24683 & x_24684;
assign x_55973 = x_24685 & x_24686;
assign x_55974 = x_55972 & x_55973;
assign x_55975 = x_55971 & x_55974;
assign x_55976 = x_24687 & x_24688;
assign x_55977 = x_24689 & x_24690;
assign x_55978 = x_55976 & x_55977;
assign x_55979 = x_24691 & x_24692;
assign x_55980 = x_24693 & x_24694;
assign x_55981 = x_55979 & x_55980;
assign x_55982 = x_55978 & x_55981;
assign x_55983 = x_55975 & x_55982;
assign x_55984 = x_55968 & x_55983;
assign x_55985 = x_55954 & x_55984;
assign x_55986 = x_55925 & x_55985;
assign x_55987 = x_55865 & x_55986;
assign x_55988 = x_24696 & x_24697;
assign x_55989 = x_24695 & x_55988;
assign x_55990 = x_24698 & x_24699;
assign x_55991 = x_24700 & x_24701;
assign x_55992 = x_55990 & x_55991;
assign x_55993 = x_55989 & x_55992;
assign x_55994 = x_24702 & x_24703;
assign x_55995 = x_24704 & x_24705;
assign x_55996 = x_55994 & x_55995;
assign x_55997 = x_24706 & x_24707;
assign x_55998 = x_24708 & x_24709;
assign x_55999 = x_55997 & x_55998;
assign x_56000 = x_55996 & x_55999;
assign x_56001 = x_55993 & x_56000;
assign x_56002 = x_24711 & x_24712;
assign x_56003 = x_24710 & x_56002;
assign x_56004 = x_24713 & x_24714;
assign x_56005 = x_24715 & x_24716;
assign x_56006 = x_56004 & x_56005;
assign x_56007 = x_56003 & x_56006;
assign x_56008 = x_24717 & x_24718;
assign x_56009 = x_24719 & x_24720;
assign x_56010 = x_56008 & x_56009;
assign x_56011 = x_24721 & x_24722;
assign x_56012 = x_24723 & x_24724;
assign x_56013 = x_56011 & x_56012;
assign x_56014 = x_56010 & x_56013;
assign x_56015 = x_56007 & x_56014;
assign x_56016 = x_56001 & x_56015;
assign x_56017 = x_24726 & x_24727;
assign x_56018 = x_24725 & x_56017;
assign x_56019 = x_24728 & x_24729;
assign x_56020 = x_24730 & x_24731;
assign x_56021 = x_56019 & x_56020;
assign x_56022 = x_56018 & x_56021;
assign x_56023 = x_24732 & x_24733;
assign x_56024 = x_24734 & x_24735;
assign x_56025 = x_56023 & x_56024;
assign x_56026 = x_24736 & x_24737;
assign x_56027 = x_24738 & x_24739;
assign x_56028 = x_56026 & x_56027;
assign x_56029 = x_56025 & x_56028;
assign x_56030 = x_56022 & x_56029;
assign x_56031 = x_24740 & x_24741;
assign x_56032 = x_24742 & x_24743;
assign x_56033 = x_56031 & x_56032;
assign x_56034 = x_24744 & x_24745;
assign x_56035 = x_24746 & x_24747;
assign x_56036 = x_56034 & x_56035;
assign x_56037 = x_56033 & x_56036;
assign x_56038 = x_24748 & x_24749;
assign x_56039 = x_24750 & x_24751;
assign x_56040 = x_56038 & x_56039;
assign x_56041 = x_24752 & x_24753;
assign x_56042 = x_24754 & x_24755;
assign x_56043 = x_56041 & x_56042;
assign x_56044 = x_56040 & x_56043;
assign x_56045 = x_56037 & x_56044;
assign x_56046 = x_56030 & x_56045;
assign x_56047 = x_56016 & x_56046;
assign x_56048 = x_24757 & x_24758;
assign x_56049 = x_24756 & x_56048;
assign x_56050 = x_24759 & x_24760;
assign x_56051 = x_24761 & x_24762;
assign x_56052 = x_56050 & x_56051;
assign x_56053 = x_56049 & x_56052;
assign x_56054 = x_24763 & x_24764;
assign x_56055 = x_24765 & x_24766;
assign x_56056 = x_56054 & x_56055;
assign x_56057 = x_24767 & x_24768;
assign x_56058 = x_24769 & x_24770;
assign x_56059 = x_56057 & x_56058;
assign x_56060 = x_56056 & x_56059;
assign x_56061 = x_56053 & x_56060;
assign x_56062 = x_24772 & x_24773;
assign x_56063 = x_24771 & x_56062;
assign x_56064 = x_24774 & x_24775;
assign x_56065 = x_24776 & x_24777;
assign x_56066 = x_56064 & x_56065;
assign x_56067 = x_56063 & x_56066;
assign x_56068 = x_24778 & x_24779;
assign x_56069 = x_24780 & x_24781;
assign x_56070 = x_56068 & x_56069;
assign x_56071 = x_24782 & x_24783;
assign x_56072 = x_24784 & x_24785;
assign x_56073 = x_56071 & x_56072;
assign x_56074 = x_56070 & x_56073;
assign x_56075 = x_56067 & x_56074;
assign x_56076 = x_56061 & x_56075;
assign x_56077 = x_24787 & x_24788;
assign x_56078 = x_24786 & x_56077;
assign x_56079 = x_24789 & x_24790;
assign x_56080 = x_24791 & x_24792;
assign x_56081 = x_56079 & x_56080;
assign x_56082 = x_56078 & x_56081;
assign x_56083 = x_24793 & x_24794;
assign x_56084 = x_24795 & x_24796;
assign x_56085 = x_56083 & x_56084;
assign x_56086 = x_24797 & x_24798;
assign x_56087 = x_24799 & x_24800;
assign x_56088 = x_56086 & x_56087;
assign x_56089 = x_56085 & x_56088;
assign x_56090 = x_56082 & x_56089;
assign x_56091 = x_24801 & x_24802;
assign x_56092 = x_24803 & x_24804;
assign x_56093 = x_56091 & x_56092;
assign x_56094 = x_24805 & x_24806;
assign x_56095 = x_24807 & x_24808;
assign x_56096 = x_56094 & x_56095;
assign x_56097 = x_56093 & x_56096;
assign x_56098 = x_24809 & x_24810;
assign x_56099 = x_24811 & x_24812;
assign x_56100 = x_56098 & x_56099;
assign x_56101 = x_24813 & x_24814;
assign x_56102 = x_24815 & x_24816;
assign x_56103 = x_56101 & x_56102;
assign x_56104 = x_56100 & x_56103;
assign x_56105 = x_56097 & x_56104;
assign x_56106 = x_56090 & x_56105;
assign x_56107 = x_56076 & x_56106;
assign x_56108 = x_56047 & x_56107;
assign x_56109 = x_24818 & x_24819;
assign x_56110 = x_24817 & x_56109;
assign x_56111 = x_24820 & x_24821;
assign x_56112 = x_24822 & x_24823;
assign x_56113 = x_56111 & x_56112;
assign x_56114 = x_56110 & x_56113;
assign x_56115 = x_24824 & x_24825;
assign x_56116 = x_24826 & x_24827;
assign x_56117 = x_56115 & x_56116;
assign x_56118 = x_24828 & x_24829;
assign x_56119 = x_24830 & x_24831;
assign x_56120 = x_56118 & x_56119;
assign x_56121 = x_56117 & x_56120;
assign x_56122 = x_56114 & x_56121;
assign x_56123 = x_24833 & x_24834;
assign x_56124 = x_24832 & x_56123;
assign x_56125 = x_24835 & x_24836;
assign x_56126 = x_24837 & x_24838;
assign x_56127 = x_56125 & x_56126;
assign x_56128 = x_56124 & x_56127;
assign x_56129 = x_24839 & x_24840;
assign x_56130 = x_24841 & x_24842;
assign x_56131 = x_56129 & x_56130;
assign x_56132 = x_24843 & x_24844;
assign x_56133 = x_24845 & x_24846;
assign x_56134 = x_56132 & x_56133;
assign x_56135 = x_56131 & x_56134;
assign x_56136 = x_56128 & x_56135;
assign x_56137 = x_56122 & x_56136;
assign x_56138 = x_24848 & x_24849;
assign x_56139 = x_24847 & x_56138;
assign x_56140 = x_24850 & x_24851;
assign x_56141 = x_24852 & x_24853;
assign x_56142 = x_56140 & x_56141;
assign x_56143 = x_56139 & x_56142;
assign x_56144 = x_24854 & x_24855;
assign x_56145 = x_24856 & x_24857;
assign x_56146 = x_56144 & x_56145;
assign x_56147 = x_24858 & x_24859;
assign x_56148 = x_24860 & x_24861;
assign x_56149 = x_56147 & x_56148;
assign x_56150 = x_56146 & x_56149;
assign x_56151 = x_56143 & x_56150;
assign x_56152 = x_24862 & x_24863;
assign x_56153 = x_24864 & x_24865;
assign x_56154 = x_56152 & x_56153;
assign x_56155 = x_24866 & x_24867;
assign x_56156 = x_24868 & x_24869;
assign x_56157 = x_56155 & x_56156;
assign x_56158 = x_56154 & x_56157;
assign x_56159 = x_24870 & x_24871;
assign x_56160 = x_24872 & x_24873;
assign x_56161 = x_56159 & x_56160;
assign x_56162 = x_24874 & x_24875;
assign x_56163 = x_24876 & x_24877;
assign x_56164 = x_56162 & x_56163;
assign x_56165 = x_56161 & x_56164;
assign x_56166 = x_56158 & x_56165;
assign x_56167 = x_56151 & x_56166;
assign x_56168 = x_56137 & x_56167;
assign x_56169 = x_24879 & x_24880;
assign x_56170 = x_24878 & x_56169;
assign x_56171 = x_24881 & x_24882;
assign x_56172 = x_24883 & x_24884;
assign x_56173 = x_56171 & x_56172;
assign x_56174 = x_56170 & x_56173;
assign x_56175 = x_24885 & x_24886;
assign x_56176 = x_24887 & x_24888;
assign x_56177 = x_56175 & x_56176;
assign x_56178 = x_24889 & x_24890;
assign x_56179 = x_24891 & x_24892;
assign x_56180 = x_56178 & x_56179;
assign x_56181 = x_56177 & x_56180;
assign x_56182 = x_56174 & x_56181;
assign x_56183 = x_24893 & x_24894;
assign x_56184 = x_24895 & x_24896;
assign x_56185 = x_56183 & x_56184;
assign x_56186 = x_24897 & x_24898;
assign x_56187 = x_24899 & x_24900;
assign x_56188 = x_56186 & x_56187;
assign x_56189 = x_56185 & x_56188;
assign x_56190 = x_24901 & x_24902;
assign x_56191 = x_24903 & x_24904;
assign x_56192 = x_56190 & x_56191;
assign x_56193 = x_24905 & x_24906;
assign x_56194 = x_24907 & x_24908;
assign x_56195 = x_56193 & x_56194;
assign x_56196 = x_56192 & x_56195;
assign x_56197 = x_56189 & x_56196;
assign x_56198 = x_56182 & x_56197;
assign x_56199 = x_24910 & x_24911;
assign x_56200 = x_24909 & x_56199;
assign x_56201 = x_24912 & x_24913;
assign x_56202 = x_24914 & x_24915;
assign x_56203 = x_56201 & x_56202;
assign x_56204 = x_56200 & x_56203;
assign x_56205 = x_24916 & x_24917;
assign x_56206 = x_24918 & x_24919;
assign x_56207 = x_56205 & x_56206;
assign x_56208 = x_24920 & x_24921;
assign x_56209 = x_24922 & x_24923;
assign x_56210 = x_56208 & x_56209;
assign x_56211 = x_56207 & x_56210;
assign x_56212 = x_56204 & x_56211;
assign x_56213 = x_24924 & x_24925;
assign x_56214 = x_24926 & x_24927;
assign x_56215 = x_56213 & x_56214;
assign x_56216 = x_24928 & x_24929;
assign x_56217 = x_24930 & x_24931;
assign x_56218 = x_56216 & x_56217;
assign x_56219 = x_56215 & x_56218;
assign x_56220 = x_24932 & x_24933;
assign x_56221 = x_24934 & x_24935;
assign x_56222 = x_56220 & x_56221;
assign x_56223 = x_24936 & x_24937;
assign x_56224 = x_24938 & x_24939;
assign x_56225 = x_56223 & x_56224;
assign x_56226 = x_56222 & x_56225;
assign x_56227 = x_56219 & x_56226;
assign x_56228 = x_56212 & x_56227;
assign x_56229 = x_56198 & x_56228;
assign x_56230 = x_56168 & x_56229;
assign x_56231 = x_56108 & x_56230;
assign x_56232 = x_55987 & x_56231;
assign x_56233 = x_24941 & x_24942;
assign x_56234 = x_24940 & x_56233;
assign x_56235 = x_24943 & x_24944;
assign x_56236 = x_24945 & x_24946;
assign x_56237 = x_56235 & x_56236;
assign x_56238 = x_56234 & x_56237;
assign x_56239 = x_24947 & x_24948;
assign x_56240 = x_24949 & x_24950;
assign x_56241 = x_56239 & x_56240;
assign x_56242 = x_24951 & x_24952;
assign x_56243 = x_24953 & x_24954;
assign x_56244 = x_56242 & x_56243;
assign x_56245 = x_56241 & x_56244;
assign x_56246 = x_56238 & x_56245;
assign x_56247 = x_24956 & x_24957;
assign x_56248 = x_24955 & x_56247;
assign x_56249 = x_24958 & x_24959;
assign x_56250 = x_24960 & x_24961;
assign x_56251 = x_56249 & x_56250;
assign x_56252 = x_56248 & x_56251;
assign x_56253 = x_24962 & x_24963;
assign x_56254 = x_24964 & x_24965;
assign x_56255 = x_56253 & x_56254;
assign x_56256 = x_24966 & x_24967;
assign x_56257 = x_24968 & x_24969;
assign x_56258 = x_56256 & x_56257;
assign x_56259 = x_56255 & x_56258;
assign x_56260 = x_56252 & x_56259;
assign x_56261 = x_56246 & x_56260;
assign x_56262 = x_24971 & x_24972;
assign x_56263 = x_24970 & x_56262;
assign x_56264 = x_24973 & x_24974;
assign x_56265 = x_24975 & x_24976;
assign x_56266 = x_56264 & x_56265;
assign x_56267 = x_56263 & x_56266;
assign x_56268 = x_24977 & x_24978;
assign x_56269 = x_24979 & x_24980;
assign x_56270 = x_56268 & x_56269;
assign x_56271 = x_24981 & x_24982;
assign x_56272 = x_24983 & x_24984;
assign x_56273 = x_56271 & x_56272;
assign x_56274 = x_56270 & x_56273;
assign x_56275 = x_56267 & x_56274;
assign x_56276 = x_24985 & x_24986;
assign x_56277 = x_24987 & x_24988;
assign x_56278 = x_56276 & x_56277;
assign x_56279 = x_24989 & x_24990;
assign x_56280 = x_24991 & x_24992;
assign x_56281 = x_56279 & x_56280;
assign x_56282 = x_56278 & x_56281;
assign x_56283 = x_24993 & x_24994;
assign x_56284 = x_24995 & x_24996;
assign x_56285 = x_56283 & x_56284;
assign x_56286 = x_24997 & x_24998;
assign x_56287 = x_24999 & x_25000;
assign x_56288 = x_56286 & x_56287;
assign x_56289 = x_56285 & x_56288;
assign x_56290 = x_56282 & x_56289;
assign x_56291 = x_56275 & x_56290;
assign x_56292 = x_56261 & x_56291;
assign x_56293 = x_25002 & x_25003;
assign x_56294 = x_25001 & x_56293;
assign x_56295 = x_25004 & x_25005;
assign x_56296 = x_25006 & x_25007;
assign x_56297 = x_56295 & x_56296;
assign x_56298 = x_56294 & x_56297;
assign x_56299 = x_25008 & x_25009;
assign x_56300 = x_25010 & x_25011;
assign x_56301 = x_56299 & x_56300;
assign x_56302 = x_25012 & x_25013;
assign x_56303 = x_25014 & x_25015;
assign x_56304 = x_56302 & x_56303;
assign x_56305 = x_56301 & x_56304;
assign x_56306 = x_56298 & x_56305;
assign x_56307 = x_25017 & x_25018;
assign x_56308 = x_25016 & x_56307;
assign x_56309 = x_25019 & x_25020;
assign x_56310 = x_25021 & x_25022;
assign x_56311 = x_56309 & x_56310;
assign x_56312 = x_56308 & x_56311;
assign x_56313 = x_25023 & x_25024;
assign x_56314 = x_25025 & x_25026;
assign x_56315 = x_56313 & x_56314;
assign x_56316 = x_25027 & x_25028;
assign x_56317 = x_25029 & x_25030;
assign x_56318 = x_56316 & x_56317;
assign x_56319 = x_56315 & x_56318;
assign x_56320 = x_56312 & x_56319;
assign x_56321 = x_56306 & x_56320;
assign x_56322 = x_25032 & x_25033;
assign x_56323 = x_25031 & x_56322;
assign x_56324 = x_25034 & x_25035;
assign x_56325 = x_25036 & x_25037;
assign x_56326 = x_56324 & x_56325;
assign x_56327 = x_56323 & x_56326;
assign x_56328 = x_25038 & x_25039;
assign x_56329 = x_25040 & x_25041;
assign x_56330 = x_56328 & x_56329;
assign x_56331 = x_25042 & x_25043;
assign x_56332 = x_25044 & x_25045;
assign x_56333 = x_56331 & x_56332;
assign x_56334 = x_56330 & x_56333;
assign x_56335 = x_56327 & x_56334;
assign x_56336 = x_25046 & x_25047;
assign x_56337 = x_25048 & x_25049;
assign x_56338 = x_56336 & x_56337;
assign x_56339 = x_25050 & x_25051;
assign x_56340 = x_25052 & x_25053;
assign x_56341 = x_56339 & x_56340;
assign x_56342 = x_56338 & x_56341;
assign x_56343 = x_25054 & x_25055;
assign x_56344 = x_25056 & x_25057;
assign x_56345 = x_56343 & x_56344;
assign x_56346 = x_25058 & x_25059;
assign x_56347 = x_25060 & x_25061;
assign x_56348 = x_56346 & x_56347;
assign x_56349 = x_56345 & x_56348;
assign x_56350 = x_56342 & x_56349;
assign x_56351 = x_56335 & x_56350;
assign x_56352 = x_56321 & x_56351;
assign x_56353 = x_56292 & x_56352;
assign x_56354 = x_25063 & x_25064;
assign x_56355 = x_25062 & x_56354;
assign x_56356 = x_25065 & x_25066;
assign x_56357 = x_25067 & x_25068;
assign x_56358 = x_56356 & x_56357;
assign x_56359 = x_56355 & x_56358;
assign x_56360 = x_25069 & x_25070;
assign x_56361 = x_25071 & x_25072;
assign x_56362 = x_56360 & x_56361;
assign x_56363 = x_25073 & x_25074;
assign x_56364 = x_25075 & x_25076;
assign x_56365 = x_56363 & x_56364;
assign x_56366 = x_56362 & x_56365;
assign x_56367 = x_56359 & x_56366;
assign x_56368 = x_25078 & x_25079;
assign x_56369 = x_25077 & x_56368;
assign x_56370 = x_25080 & x_25081;
assign x_56371 = x_25082 & x_25083;
assign x_56372 = x_56370 & x_56371;
assign x_56373 = x_56369 & x_56372;
assign x_56374 = x_25084 & x_25085;
assign x_56375 = x_25086 & x_25087;
assign x_56376 = x_56374 & x_56375;
assign x_56377 = x_25088 & x_25089;
assign x_56378 = x_25090 & x_25091;
assign x_56379 = x_56377 & x_56378;
assign x_56380 = x_56376 & x_56379;
assign x_56381 = x_56373 & x_56380;
assign x_56382 = x_56367 & x_56381;
assign x_56383 = x_25093 & x_25094;
assign x_56384 = x_25092 & x_56383;
assign x_56385 = x_25095 & x_25096;
assign x_56386 = x_25097 & x_25098;
assign x_56387 = x_56385 & x_56386;
assign x_56388 = x_56384 & x_56387;
assign x_56389 = x_25099 & x_25100;
assign x_56390 = x_25101 & x_25102;
assign x_56391 = x_56389 & x_56390;
assign x_56392 = x_25103 & x_25104;
assign x_56393 = x_25105 & x_25106;
assign x_56394 = x_56392 & x_56393;
assign x_56395 = x_56391 & x_56394;
assign x_56396 = x_56388 & x_56395;
assign x_56397 = x_25107 & x_25108;
assign x_56398 = x_25109 & x_25110;
assign x_56399 = x_56397 & x_56398;
assign x_56400 = x_25111 & x_25112;
assign x_56401 = x_25113 & x_25114;
assign x_56402 = x_56400 & x_56401;
assign x_56403 = x_56399 & x_56402;
assign x_56404 = x_25115 & x_25116;
assign x_56405 = x_25117 & x_25118;
assign x_56406 = x_56404 & x_56405;
assign x_56407 = x_25119 & x_25120;
assign x_56408 = x_25121 & x_25122;
assign x_56409 = x_56407 & x_56408;
assign x_56410 = x_56406 & x_56409;
assign x_56411 = x_56403 & x_56410;
assign x_56412 = x_56396 & x_56411;
assign x_56413 = x_56382 & x_56412;
assign x_56414 = x_25124 & x_25125;
assign x_56415 = x_25123 & x_56414;
assign x_56416 = x_25126 & x_25127;
assign x_56417 = x_25128 & x_25129;
assign x_56418 = x_56416 & x_56417;
assign x_56419 = x_56415 & x_56418;
assign x_56420 = x_25130 & x_25131;
assign x_56421 = x_25132 & x_25133;
assign x_56422 = x_56420 & x_56421;
assign x_56423 = x_25134 & x_25135;
assign x_56424 = x_25136 & x_25137;
assign x_56425 = x_56423 & x_56424;
assign x_56426 = x_56422 & x_56425;
assign x_56427 = x_56419 & x_56426;
assign x_56428 = x_25139 & x_25140;
assign x_56429 = x_25138 & x_56428;
assign x_56430 = x_25141 & x_25142;
assign x_56431 = x_25143 & x_25144;
assign x_56432 = x_56430 & x_56431;
assign x_56433 = x_56429 & x_56432;
assign x_56434 = x_25145 & x_25146;
assign x_56435 = x_25147 & x_25148;
assign x_56436 = x_56434 & x_56435;
assign x_56437 = x_25149 & x_25150;
assign x_56438 = x_25151 & x_25152;
assign x_56439 = x_56437 & x_56438;
assign x_56440 = x_56436 & x_56439;
assign x_56441 = x_56433 & x_56440;
assign x_56442 = x_56427 & x_56441;
assign x_56443 = x_25154 & x_25155;
assign x_56444 = x_25153 & x_56443;
assign x_56445 = x_25156 & x_25157;
assign x_56446 = x_25158 & x_25159;
assign x_56447 = x_56445 & x_56446;
assign x_56448 = x_56444 & x_56447;
assign x_56449 = x_25160 & x_25161;
assign x_56450 = x_25162 & x_25163;
assign x_56451 = x_56449 & x_56450;
assign x_56452 = x_25164 & x_25165;
assign x_56453 = x_25166 & x_25167;
assign x_56454 = x_56452 & x_56453;
assign x_56455 = x_56451 & x_56454;
assign x_56456 = x_56448 & x_56455;
assign x_56457 = x_25168 & x_25169;
assign x_56458 = x_25170 & x_25171;
assign x_56459 = x_56457 & x_56458;
assign x_56460 = x_25172 & x_25173;
assign x_56461 = x_25174 & x_25175;
assign x_56462 = x_56460 & x_56461;
assign x_56463 = x_56459 & x_56462;
assign x_56464 = x_25176 & x_25177;
assign x_56465 = x_25178 & x_25179;
assign x_56466 = x_56464 & x_56465;
assign x_56467 = x_25180 & x_25181;
assign x_56468 = x_25182 & x_25183;
assign x_56469 = x_56467 & x_56468;
assign x_56470 = x_56466 & x_56469;
assign x_56471 = x_56463 & x_56470;
assign x_56472 = x_56456 & x_56471;
assign x_56473 = x_56442 & x_56472;
assign x_56474 = x_56413 & x_56473;
assign x_56475 = x_56353 & x_56474;
assign x_56476 = x_25185 & x_25186;
assign x_56477 = x_25184 & x_56476;
assign x_56478 = x_25187 & x_25188;
assign x_56479 = x_25189 & x_25190;
assign x_56480 = x_56478 & x_56479;
assign x_56481 = x_56477 & x_56480;
assign x_56482 = x_25191 & x_25192;
assign x_56483 = x_25193 & x_25194;
assign x_56484 = x_56482 & x_56483;
assign x_56485 = x_25195 & x_25196;
assign x_56486 = x_25197 & x_25198;
assign x_56487 = x_56485 & x_56486;
assign x_56488 = x_56484 & x_56487;
assign x_56489 = x_56481 & x_56488;
assign x_56490 = x_25200 & x_25201;
assign x_56491 = x_25199 & x_56490;
assign x_56492 = x_25202 & x_25203;
assign x_56493 = x_25204 & x_25205;
assign x_56494 = x_56492 & x_56493;
assign x_56495 = x_56491 & x_56494;
assign x_56496 = x_25206 & x_25207;
assign x_56497 = x_25208 & x_25209;
assign x_56498 = x_56496 & x_56497;
assign x_56499 = x_25210 & x_25211;
assign x_56500 = x_25212 & x_25213;
assign x_56501 = x_56499 & x_56500;
assign x_56502 = x_56498 & x_56501;
assign x_56503 = x_56495 & x_56502;
assign x_56504 = x_56489 & x_56503;
assign x_56505 = x_25215 & x_25216;
assign x_56506 = x_25214 & x_56505;
assign x_56507 = x_25217 & x_25218;
assign x_56508 = x_25219 & x_25220;
assign x_56509 = x_56507 & x_56508;
assign x_56510 = x_56506 & x_56509;
assign x_56511 = x_25221 & x_25222;
assign x_56512 = x_25223 & x_25224;
assign x_56513 = x_56511 & x_56512;
assign x_56514 = x_25225 & x_25226;
assign x_56515 = x_25227 & x_25228;
assign x_56516 = x_56514 & x_56515;
assign x_56517 = x_56513 & x_56516;
assign x_56518 = x_56510 & x_56517;
assign x_56519 = x_25229 & x_25230;
assign x_56520 = x_25231 & x_25232;
assign x_56521 = x_56519 & x_56520;
assign x_56522 = x_25233 & x_25234;
assign x_56523 = x_25235 & x_25236;
assign x_56524 = x_56522 & x_56523;
assign x_56525 = x_56521 & x_56524;
assign x_56526 = x_25237 & x_25238;
assign x_56527 = x_25239 & x_25240;
assign x_56528 = x_56526 & x_56527;
assign x_56529 = x_25241 & x_25242;
assign x_56530 = x_25243 & x_25244;
assign x_56531 = x_56529 & x_56530;
assign x_56532 = x_56528 & x_56531;
assign x_56533 = x_56525 & x_56532;
assign x_56534 = x_56518 & x_56533;
assign x_56535 = x_56504 & x_56534;
assign x_56536 = x_25246 & x_25247;
assign x_56537 = x_25245 & x_56536;
assign x_56538 = x_25248 & x_25249;
assign x_56539 = x_25250 & x_25251;
assign x_56540 = x_56538 & x_56539;
assign x_56541 = x_56537 & x_56540;
assign x_56542 = x_25252 & x_25253;
assign x_56543 = x_25254 & x_25255;
assign x_56544 = x_56542 & x_56543;
assign x_56545 = x_25256 & x_25257;
assign x_56546 = x_25258 & x_25259;
assign x_56547 = x_56545 & x_56546;
assign x_56548 = x_56544 & x_56547;
assign x_56549 = x_56541 & x_56548;
assign x_56550 = x_25261 & x_25262;
assign x_56551 = x_25260 & x_56550;
assign x_56552 = x_25263 & x_25264;
assign x_56553 = x_25265 & x_25266;
assign x_56554 = x_56552 & x_56553;
assign x_56555 = x_56551 & x_56554;
assign x_56556 = x_25267 & x_25268;
assign x_56557 = x_25269 & x_25270;
assign x_56558 = x_56556 & x_56557;
assign x_56559 = x_25271 & x_25272;
assign x_56560 = x_25273 & x_25274;
assign x_56561 = x_56559 & x_56560;
assign x_56562 = x_56558 & x_56561;
assign x_56563 = x_56555 & x_56562;
assign x_56564 = x_56549 & x_56563;
assign x_56565 = x_25276 & x_25277;
assign x_56566 = x_25275 & x_56565;
assign x_56567 = x_25278 & x_25279;
assign x_56568 = x_25280 & x_25281;
assign x_56569 = x_56567 & x_56568;
assign x_56570 = x_56566 & x_56569;
assign x_56571 = x_25282 & x_25283;
assign x_56572 = x_25284 & x_25285;
assign x_56573 = x_56571 & x_56572;
assign x_56574 = x_25286 & x_25287;
assign x_56575 = x_25288 & x_25289;
assign x_56576 = x_56574 & x_56575;
assign x_56577 = x_56573 & x_56576;
assign x_56578 = x_56570 & x_56577;
assign x_56579 = x_25290 & x_25291;
assign x_56580 = x_25292 & x_25293;
assign x_56581 = x_56579 & x_56580;
assign x_56582 = x_25294 & x_25295;
assign x_56583 = x_25296 & x_25297;
assign x_56584 = x_56582 & x_56583;
assign x_56585 = x_56581 & x_56584;
assign x_56586 = x_25298 & x_25299;
assign x_56587 = x_25300 & x_25301;
assign x_56588 = x_56586 & x_56587;
assign x_56589 = x_25302 & x_25303;
assign x_56590 = x_25304 & x_25305;
assign x_56591 = x_56589 & x_56590;
assign x_56592 = x_56588 & x_56591;
assign x_56593 = x_56585 & x_56592;
assign x_56594 = x_56578 & x_56593;
assign x_56595 = x_56564 & x_56594;
assign x_56596 = x_56535 & x_56595;
assign x_56597 = x_25307 & x_25308;
assign x_56598 = x_25306 & x_56597;
assign x_56599 = x_25309 & x_25310;
assign x_56600 = x_25311 & x_25312;
assign x_56601 = x_56599 & x_56600;
assign x_56602 = x_56598 & x_56601;
assign x_56603 = x_25313 & x_25314;
assign x_56604 = x_25315 & x_25316;
assign x_56605 = x_56603 & x_56604;
assign x_56606 = x_25317 & x_25318;
assign x_56607 = x_25319 & x_25320;
assign x_56608 = x_56606 & x_56607;
assign x_56609 = x_56605 & x_56608;
assign x_56610 = x_56602 & x_56609;
assign x_56611 = x_25322 & x_25323;
assign x_56612 = x_25321 & x_56611;
assign x_56613 = x_25324 & x_25325;
assign x_56614 = x_25326 & x_25327;
assign x_56615 = x_56613 & x_56614;
assign x_56616 = x_56612 & x_56615;
assign x_56617 = x_25328 & x_25329;
assign x_56618 = x_25330 & x_25331;
assign x_56619 = x_56617 & x_56618;
assign x_56620 = x_25332 & x_25333;
assign x_56621 = x_25334 & x_25335;
assign x_56622 = x_56620 & x_56621;
assign x_56623 = x_56619 & x_56622;
assign x_56624 = x_56616 & x_56623;
assign x_56625 = x_56610 & x_56624;
assign x_56626 = x_25337 & x_25338;
assign x_56627 = x_25336 & x_56626;
assign x_56628 = x_25339 & x_25340;
assign x_56629 = x_25341 & x_25342;
assign x_56630 = x_56628 & x_56629;
assign x_56631 = x_56627 & x_56630;
assign x_56632 = x_25343 & x_25344;
assign x_56633 = x_25345 & x_25346;
assign x_56634 = x_56632 & x_56633;
assign x_56635 = x_25347 & x_25348;
assign x_56636 = x_25349 & x_25350;
assign x_56637 = x_56635 & x_56636;
assign x_56638 = x_56634 & x_56637;
assign x_56639 = x_56631 & x_56638;
assign x_56640 = x_25351 & x_25352;
assign x_56641 = x_25353 & x_25354;
assign x_56642 = x_56640 & x_56641;
assign x_56643 = x_25355 & x_25356;
assign x_56644 = x_25357 & x_25358;
assign x_56645 = x_56643 & x_56644;
assign x_56646 = x_56642 & x_56645;
assign x_56647 = x_25359 & x_25360;
assign x_56648 = x_25361 & x_25362;
assign x_56649 = x_56647 & x_56648;
assign x_56650 = x_25363 & x_25364;
assign x_56651 = x_25365 & x_25366;
assign x_56652 = x_56650 & x_56651;
assign x_56653 = x_56649 & x_56652;
assign x_56654 = x_56646 & x_56653;
assign x_56655 = x_56639 & x_56654;
assign x_56656 = x_56625 & x_56655;
assign x_56657 = x_25368 & x_25369;
assign x_56658 = x_25367 & x_56657;
assign x_56659 = x_25370 & x_25371;
assign x_56660 = x_25372 & x_25373;
assign x_56661 = x_56659 & x_56660;
assign x_56662 = x_56658 & x_56661;
assign x_56663 = x_25374 & x_25375;
assign x_56664 = x_25376 & x_25377;
assign x_56665 = x_56663 & x_56664;
assign x_56666 = x_25378 & x_25379;
assign x_56667 = x_25380 & x_25381;
assign x_56668 = x_56666 & x_56667;
assign x_56669 = x_56665 & x_56668;
assign x_56670 = x_56662 & x_56669;
assign x_56671 = x_25382 & x_25383;
assign x_56672 = x_25384 & x_25385;
assign x_56673 = x_56671 & x_56672;
assign x_56674 = x_25386 & x_25387;
assign x_56675 = x_25388 & x_25389;
assign x_56676 = x_56674 & x_56675;
assign x_56677 = x_56673 & x_56676;
assign x_56678 = x_25390 & x_25391;
assign x_56679 = x_25392 & x_25393;
assign x_56680 = x_56678 & x_56679;
assign x_56681 = x_25394 & x_25395;
assign x_56682 = x_25396 & x_25397;
assign x_56683 = x_56681 & x_56682;
assign x_56684 = x_56680 & x_56683;
assign x_56685 = x_56677 & x_56684;
assign x_56686 = x_56670 & x_56685;
assign x_56687 = x_25399 & x_25400;
assign x_56688 = x_25398 & x_56687;
assign x_56689 = x_25401 & x_25402;
assign x_56690 = x_25403 & x_25404;
assign x_56691 = x_56689 & x_56690;
assign x_56692 = x_56688 & x_56691;
assign x_56693 = x_25405 & x_25406;
assign x_56694 = x_25407 & x_25408;
assign x_56695 = x_56693 & x_56694;
assign x_56696 = x_25409 & x_25410;
assign x_56697 = x_25411 & x_25412;
assign x_56698 = x_56696 & x_56697;
assign x_56699 = x_56695 & x_56698;
assign x_56700 = x_56692 & x_56699;
assign x_56701 = x_25413 & x_25414;
assign x_56702 = x_25415 & x_25416;
assign x_56703 = x_56701 & x_56702;
assign x_56704 = x_25417 & x_25418;
assign x_56705 = x_25419 & x_25420;
assign x_56706 = x_56704 & x_56705;
assign x_56707 = x_56703 & x_56706;
assign x_56708 = x_25421 & x_25422;
assign x_56709 = x_25423 & x_25424;
assign x_56710 = x_56708 & x_56709;
assign x_56711 = x_25425 & x_25426;
assign x_56712 = x_25427 & x_25428;
assign x_56713 = x_56711 & x_56712;
assign x_56714 = x_56710 & x_56713;
assign x_56715 = x_56707 & x_56714;
assign x_56716 = x_56700 & x_56715;
assign x_56717 = x_56686 & x_56716;
assign x_56718 = x_56656 & x_56717;
assign x_56719 = x_56596 & x_56718;
assign x_56720 = x_56475 & x_56719;
assign x_56721 = x_56232 & x_56720;
assign x_56722 = x_55744 & x_56721;
assign x_56723 = x_25430 & x_25431;
assign x_56724 = x_25429 & x_56723;
assign x_56725 = x_25432 & x_25433;
assign x_56726 = x_25434 & x_25435;
assign x_56727 = x_56725 & x_56726;
assign x_56728 = x_56724 & x_56727;
assign x_56729 = x_25436 & x_25437;
assign x_56730 = x_25438 & x_25439;
assign x_56731 = x_56729 & x_56730;
assign x_56732 = x_25440 & x_25441;
assign x_56733 = x_25442 & x_25443;
assign x_56734 = x_56732 & x_56733;
assign x_56735 = x_56731 & x_56734;
assign x_56736 = x_56728 & x_56735;
assign x_56737 = x_25445 & x_25446;
assign x_56738 = x_25444 & x_56737;
assign x_56739 = x_25447 & x_25448;
assign x_56740 = x_25449 & x_25450;
assign x_56741 = x_56739 & x_56740;
assign x_56742 = x_56738 & x_56741;
assign x_56743 = x_25451 & x_25452;
assign x_56744 = x_25453 & x_25454;
assign x_56745 = x_56743 & x_56744;
assign x_56746 = x_25455 & x_25456;
assign x_56747 = x_25457 & x_25458;
assign x_56748 = x_56746 & x_56747;
assign x_56749 = x_56745 & x_56748;
assign x_56750 = x_56742 & x_56749;
assign x_56751 = x_56736 & x_56750;
assign x_56752 = x_25460 & x_25461;
assign x_56753 = x_25459 & x_56752;
assign x_56754 = x_25462 & x_25463;
assign x_56755 = x_25464 & x_25465;
assign x_56756 = x_56754 & x_56755;
assign x_56757 = x_56753 & x_56756;
assign x_56758 = x_25466 & x_25467;
assign x_56759 = x_25468 & x_25469;
assign x_56760 = x_56758 & x_56759;
assign x_56761 = x_25470 & x_25471;
assign x_56762 = x_25472 & x_25473;
assign x_56763 = x_56761 & x_56762;
assign x_56764 = x_56760 & x_56763;
assign x_56765 = x_56757 & x_56764;
assign x_56766 = x_25474 & x_25475;
assign x_56767 = x_25476 & x_25477;
assign x_56768 = x_56766 & x_56767;
assign x_56769 = x_25478 & x_25479;
assign x_56770 = x_25480 & x_25481;
assign x_56771 = x_56769 & x_56770;
assign x_56772 = x_56768 & x_56771;
assign x_56773 = x_25482 & x_25483;
assign x_56774 = x_25484 & x_25485;
assign x_56775 = x_56773 & x_56774;
assign x_56776 = x_25486 & x_25487;
assign x_56777 = x_25488 & x_25489;
assign x_56778 = x_56776 & x_56777;
assign x_56779 = x_56775 & x_56778;
assign x_56780 = x_56772 & x_56779;
assign x_56781 = x_56765 & x_56780;
assign x_56782 = x_56751 & x_56781;
assign x_56783 = x_25491 & x_25492;
assign x_56784 = x_25490 & x_56783;
assign x_56785 = x_25493 & x_25494;
assign x_56786 = x_25495 & x_25496;
assign x_56787 = x_56785 & x_56786;
assign x_56788 = x_56784 & x_56787;
assign x_56789 = x_25497 & x_25498;
assign x_56790 = x_25499 & x_25500;
assign x_56791 = x_56789 & x_56790;
assign x_56792 = x_25501 & x_25502;
assign x_56793 = x_25503 & x_25504;
assign x_56794 = x_56792 & x_56793;
assign x_56795 = x_56791 & x_56794;
assign x_56796 = x_56788 & x_56795;
assign x_56797 = x_25506 & x_25507;
assign x_56798 = x_25505 & x_56797;
assign x_56799 = x_25508 & x_25509;
assign x_56800 = x_25510 & x_25511;
assign x_56801 = x_56799 & x_56800;
assign x_56802 = x_56798 & x_56801;
assign x_56803 = x_25512 & x_25513;
assign x_56804 = x_25514 & x_25515;
assign x_56805 = x_56803 & x_56804;
assign x_56806 = x_25516 & x_25517;
assign x_56807 = x_25518 & x_25519;
assign x_56808 = x_56806 & x_56807;
assign x_56809 = x_56805 & x_56808;
assign x_56810 = x_56802 & x_56809;
assign x_56811 = x_56796 & x_56810;
assign x_56812 = x_25521 & x_25522;
assign x_56813 = x_25520 & x_56812;
assign x_56814 = x_25523 & x_25524;
assign x_56815 = x_25525 & x_25526;
assign x_56816 = x_56814 & x_56815;
assign x_56817 = x_56813 & x_56816;
assign x_56818 = x_25527 & x_25528;
assign x_56819 = x_25529 & x_25530;
assign x_56820 = x_56818 & x_56819;
assign x_56821 = x_25531 & x_25532;
assign x_56822 = x_25533 & x_25534;
assign x_56823 = x_56821 & x_56822;
assign x_56824 = x_56820 & x_56823;
assign x_56825 = x_56817 & x_56824;
assign x_56826 = x_25535 & x_25536;
assign x_56827 = x_25537 & x_25538;
assign x_56828 = x_56826 & x_56827;
assign x_56829 = x_25539 & x_25540;
assign x_56830 = x_25541 & x_25542;
assign x_56831 = x_56829 & x_56830;
assign x_56832 = x_56828 & x_56831;
assign x_56833 = x_25543 & x_25544;
assign x_56834 = x_25545 & x_25546;
assign x_56835 = x_56833 & x_56834;
assign x_56836 = x_25547 & x_25548;
assign x_56837 = x_25549 & x_25550;
assign x_56838 = x_56836 & x_56837;
assign x_56839 = x_56835 & x_56838;
assign x_56840 = x_56832 & x_56839;
assign x_56841 = x_56825 & x_56840;
assign x_56842 = x_56811 & x_56841;
assign x_56843 = x_56782 & x_56842;
assign x_56844 = x_25552 & x_25553;
assign x_56845 = x_25551 & x_56844;
assign x_56846 = x_25554 & x_25555;
assign x_56847 = x_25556 & x_25557;
assign x_56848 = x_56846 & x_56847;
assign x_56849 = x_56845 & x_56848;
assign x_56850 = x_25558 & x_25559;
assign x_56851 = x_25560 & x_25561;
assign x_56852 = x_56850 & x_56851;
assign x_56853 = x_25562 & x_25563;
assign x_56854 = x_25564 & x_25565;
assign x_56855 = x_56853 & x_56854;
assign x_56856 = x_56852 & x_56855;
assign x_56857 = x_56849 & x_56856;
assign x_56858 = x_25567 & x_25568;
assign x_56859 = x_25566 & x_56858;
assign x_56860 = x_25569 & x_25570;
assign x_56861 = x_25571 & x_25572;
assign x_56862 = x_56860 & x_56861;
assign x_56863 = x_56859 & x_56862;
assign x_56864 = x_25573 & x_25574;
assign x_56865 = x_25575 & x_25576;
assign x_56866 = x_56864 & x_56865;
assign x_56867 = x_25577 & x_25578;
assign x_56868 = x_25579 & x_25580;
assign x_56869 = x_56867 & x_56868;
assign x_56870 = x_56866 & x_56869;
assign x_56871 = x_56863 & x_56870;
assign x_56872 = x_56857 & x_56871;
assign x_56873 = x_25582 & x_25583;
assign x_56874 = x_25581 & x_56873;
assign x_56875 = x_25584 & x_25585;
assign x_56876 = x_25586 & x_25587;
assign x_56877 = x_56875 & x_56876;
assign x_56878 = x_56874 & x_56877;
assign x_56879 = x_25588 & x_25589;
assign x_56880 = x_25590 & x_25591;
assign x_56881 = x_56879 & x_56880;
assign x_56882 = x_25592 & x_25593;
assign x_56883 = x_25594 & x_25595;
assign x_56884 = x_56882 & x_56883;
assign x_56885 = x_56881 & x_56884;
assign x_56886 = x_56878 & x_56885;
assign x_56887 = x_25596 & x_25597;
assign x_56888 = x_25598 & x_25599;
assign x_56889 = x_56887 & x_56888;
assign x_56890 = x_25600 & x_25601;
assign x_56891 = x_25602 & x_25603;
assign x_56892 = x_56890 & x_56891;
assign x_56893 = x_56889 & x_56892;
assign x_56894 = x_25604 & x_25605;
assign x_56895 = x_25606 & x_25607;
assign x_56896 = x_56894 & x_56895;
assign x_56897 = x_25608 & x_25609;
assign x_56898 = x_25610 & x_25611;
assign x_56899 = x_56897 & x_56898;
assign x_56900 = x_56896 & x_56899;
assign x_56901 = x_56893 & x_56900;
assign x_56902 = x_56886 & x_56901;
assign x_56903 = x_56872 & x_56902;
assign x_56904 = x_25613 & x_25614;
assign x_56905 = x_25612 & x_56904;
assign x_56906 = x_25615 & x_25616;
assign x_56907 = x_25617 & x_25618;
assign x_56908 = x_56906 & x_56907;
assign x_56909 = x_56905 & x_56908;
assign x_56910 = x_25619 & x_25620;
assign x_56911 = x_25621 & x_25622;
assign x_56912 = x_56910 & x_56911;
assign x_56913 = x_25623 & x_25624;
assign x_56914 = x_25625 & x_25626;
assign x_56915 = x_56913 & x_56914;
assign x_56916 = x_56912 & x_56915;
assign x_56917 = x_56909 & x_56916;
assign x_56918 = x_25628 & x_25629;
assign x_56919 = x_25627 & x_56918;
assign x_56920 = x_25630 & x_25631;
assign x_56921 = x_25632 & x_25633;
assign x_56922 = x_56920 & x_56921;
assign x_56923 = x_56919 & x_56922;
assign x_56924 = x_25634 & x_25635;
assign x_56925 = x_25636 & x_25637;
assign x_56926 = x_56924 & x_56925;
assign x_56927 = x_25638 & x_25639;
assign x_56928 = x_25640 & x_25641;
assign x_56929 = x_56927 & x_56928;
assign x_56930 = x_56926 & x_56929;
assign x_56931 = x_56923 & x_56930;
assign x_56932 = x_56917 & x_56931;
assign x_56933 = x_25643 & x_25644;
assign x_56934 = x_25642 & x_56933;
assign x_56935 = x_25645 & x_25646;
assign x_56936 = x_25647 & x_25648;
assign x_56937 = x_56935 & x_56936;
assign x_56938 = x_56934 & x_56937;
assign x_56939 = x_25649 & x_25650;
assign x_56940 = x_25651 & x_25652;
assign x_56941 = x_56939 & x_56940;
assign x_56942 = x_25653 & x_25654;
assign x_56943 = x_25655 & x_25656;
assign x_56944 = x_56942 & x_56943;
assign x_56945 = x_56941 & x_56944;
assign x_56946 = x_56938 & x_56945;
assign x_56947 = x_25657 & x_25658;
assign x_56948 = x_25659 & x_25660;
assign x_56949 = x_56947 & x_56948;
assign x_56950 = x_25661 & x_25662;
assign x_56951 = x_25663 & x_25664;
assign x_56952 = x_56950 & x_56951;
assign x_56953 = x_56949 & x_56952;
assign x_56954 = x_25665 & x_25666;
assign x_56955 = x_25667 & x_25668;
assign x_56956 = x_56954 & x_56955;
assign x_56957 = x_25669 & x_25670;
assign x_56958 = x_25671 & x_25672;
assign x_56959 = x_56957 & x_56958;
assign x_56960 = x_56956 & x_56959;
assign x_56961 = x_56953 & x_56960;
assign x_56962 = x_56946 & x_56961;
assign x_56963 = x_56932 & x_56962;
assign x_56964 = x_56903 & x_56963;
assign x_56965 = x_56843 & x_56964;
assign x_56966 = x_25674 & x_25675;
assign x_56967 = x_25673 & x_56966;
assign x_56968 = x_25676 & x_25677;
assign x_56969 = x_25678 & x_25679;
assign x_56970 = x_56968 & x_56969;
assign x_56971 = x_56967 & x_56970;
assign x_56972 = x_25680 & x_25681;
assign x_56973 = x_25682 & x_25683;
assign x_56974 = x_56972 & x_56973;
assign x_56975 = x_25684 & x_25685;
assign x_56976 = x_25686 & x_25687;
assign x_56977 = x_56975 & x_56976;
assign x_56978 = x_56974 & x_56977;
assign x_56979 = x_56971 & x_56978;
assign x_56980 = x_25689 & x_25690;
assign x_56981 = x_25688 & x_56980;
assign x_56982 = x_25691 & x_25692;
assign x_56983 = x_25693 & x_25694;
assign x_56984 = x_56982 & x_56983;
assign x_56985 = x_56981 & x_56984;
assign x_56986 = x_25695 & x_25696;
assign x_56987 = x_25697 & x_25698;
assign x_56988 = x_56986 & x_56987;
assign x_56989 = x_25699 & x_25700;
assign x_56990 = x_25701 & x_25702;
assign x_56991 = x_56989 & x_56990;
assign x_56992 = x_56988 & x_56991;
assign x_56993 = x_56985 & x_56992;
assign x_56994 = x_56979 & x_56993;
assign x_56995 = x_25704 & x_25705;
assign x_56996 = x_25703 & x_56995;
assign x_56997 = x_25706 & x_25707;
assign x_56998 = x_25708 & x_25709;
assign x_56999 = x_56997 & x_56998;
assign x_57000 = x_56996 & x_56999;
assign x_57001 = x_25710 & x_25711;
assign x_57002 = x_25712 & x_25713;
assign x_57003 = x_57001 & x_57002;
assign x_57004 = x_25714 & x_25715;
assign x_57005 = x_25716 & x_25717;
assign x_57006 = x_57004 & x_57005;
assign x_57007 = x_57003 & x_57006;
assign x_57008 = x_57000 & x_57007;
assign x_57009 = x_25718 & x_25719;
assign x_57010 = x_25720 & x_25721;
assign x_57011 = x_57009 & x_57010;
assign x_57012 = x_25722 & x_25723;
assign x_57013 = x_25724 & x_25725;
assign x_57014 = x_57012 & x_57013;
assign x_57015 = x_57011 & x_57014;
assign x_57016 = x_25726 & x_25727;
assign x_57017 = x_25728 & x_25729;
assign x_57018 = x_57016 & x_57017;
assign x_57019 = x_25730 & x_25731;
assign x_57020 = x_25732 & x_25733;
assign x_57021 = x_57019 & x_57020;
assign x_57022 = x_57018 & x_57021;
assign x_57023 = x_57015 & x_57022;
assign x_57024 = x_57008 & x_57023;
assign x_57025 = x_56994 & x_57024;
assign x_57026 = x_25735 & x_25736;
assign x_57027 = x_25734 & x_57026;
assign x_57028 = x_25737 & x_25738;
assign x_57029 = x_25739 & x_25740;
assign x_57030 = x_57028 & x_57029;
assign x_57031 = x_57027 & x_57030;
assign x_57032 = x_25741 & x_25742;
assign x_57033 = x_25743 & x_25744;
assign x_57034 = x_57032 & x_57033;
assign x_57035 = x_25745 & x_25746;
assign x_57036 = x_25747 & x_25748;
assign x_57037 = x_57035 & x_57036;
assign x_57038 = x_57034 & x_57037;
assign x_57039 = x_57031 & x_57038;
assign x_57040 = x_25750 & x_25751;
assign x_57041 = x_25749 & x_57040;
assign x_57042 = x_25752 & x_25753;
assign x_57043 = x_25754 & x_25755;
assign x_57044 = x_57042 & x_57043;
assign x_57045 = x_57041 & x_57044;
assign x_57046 = x_25756 & x_25757;
assign x_57047 = x_25758 & x_25759;
assign x_57048 = x_57046 & x_57047;
assign x_57049 = x_25760 & x_25761;
assign x_57050 = x_25762 & x_25763;
assign x_57051 = x_57049 & x_57050;
assign x_57052 = x_57048 & x_57051;
assign x_57053 = x_57045 & x_57052;
assign x_57054 = x_57039 & x_57053;
assign x_57055 = x_25765 & x_25766;
assign x_57056 = x_25764 & x_57055;
assign x_57057 = x_25767 & x_25768;
assign x_57058 = x_25769 & x_25770;
assign x_57059 = x_57057 & x_57058;
assign x_57060 = x_57056 & x_57059;
assign x_57061 = x_25771 & x_25772;
assign x_57062 = x_25773 & x_25774;
assign x_57063 = x_57061 & x_57062;
assign x_57064 = x_25775 & x_25776;
assign x_57065 = x_25777 & x_25778;
assign x_57066 = x_57064 & x_57065;
assign x_57067 = x_57063 & x_57066;
assign x_57068 = x_57060 & x_57067;
assign x_57069 = x_25779 & x_25780;
assign x_57070 = x_25781 & x_25782;
assign x_57071 = x_57069 & x_57070;
assign x_57072 = x_25783 & x_25784;
assign x_57073 = x_25785 & x_25786;
assign x_57074 = x_57072 & x_57073;
assign x_57075 = x_57071 & x_57074;
assign x_57076 = x_25787 & x_25788;
assign x_57077 = x_25789 & x_25790;
assign x_57078 = x_57076 & x_57077;
assign x_57079 = x_25791 & x_25792;
assign x_57080 = x_25793 & x_25794;
assign x_57081 = x_57079 & x_57080;
assign x_57082 = x_57078 & x_57081;
assign x_57083 = x_57075 & x_57082;
assign x_57084 = x_57068 & x_57083;
assign x_57085 = x_57054 & x_57084;
assign x_57086 = x_57025 & x_57085;
assign x_57087 = x_25796 & x_25797;
assign x_57088 = x_25795 & x_57087;
assign x_57089 = x_25798 & x_25799;
assign x_57090 = x_25800 & x_25801;
assign x_57091 = x_57089 & x_57090;
assign x_57092 = x_57088 & x_57091;
assign x_57093 = x_25802 & x_25803;
assign x_57094 = x_25804 & x_25805;
assign x_57095 = x_57093 & x_57094;
assign x_57096 = x_25806 & x_25807;
assign x_57097 = x_25808 & x_25809;
assign x_57098 = x_57096 & x_57097;
assign x_57099 = x_57095 & x_57098;
assign x_57100 = x_57092 & x_57099;
assign x_57101 = x_25811 & x_25812;
assign x_57102 = x_25810 & x_57101;
assign x_57103 = x_25813 & x_25814;
assign x_57104 = x_25815 & x_25816;
assign x_57105 = x_57103 & x_57104;
assign x_57106 = x_57102 & x_57105;
assign x_57107 = x_25817 & x_25818;
assign x_57108 = x_25819 & x_25820;
assign x_57109 = x_57107 & x_57108;
assign x_57110 = x_25821 & x_25822;
assign x_57111 = x_25823 & x_25824;
assign x_57112 = x_57110 & x_57111;
assign x_57113 = x_57109 & x_57112;
assign x_57114 = x_57106 & x_57113;
assign x_57115 = x_57100 & x_57114;
assign x_57116 = x_25826 & x_25827;
assign x_57117 = x_25825 & x_57116;
assign x_57118 = x_25828 & x_25829;
assign x_57119 = x_25830 & x_25831;
assign x_57120 = x_57118 & x_57119;
assign x_57121 = x_57117 & x_57120;
assign x_57122 = x_25832 & x_25833;
assign x_57123 = x_25834 & x_25835;
assign x_57124 = x_57122 & x_57123;
assign x_57125 = x_25836 & x_25837;
assign x_57126 = x_25838 & x_25839;
assign x_57127 = x_57125 & x_57126;
assign x_57128 = x_57124 & x_57127;
assign x_57129 = x_57121 & x_57128;
assign x_57130 = x_25840 & x_25841;
assign x_57131 = x_25842 & x_25843;
assign x_57132 = x_57130 & x_57131;
assign x_57133 = x_25844 & x_25845;
assign x_57134 = x_25846 & x_25847;
assign x_57135 = x_57133 & x_57134;
assign x_57136 = x_57132 & x_57135;
assign x_57137 = x_25848 & x_25849;
assign x_57138 = x_25850 & x_25851;
assign x_57139 = x_57137 & x_57138;
assign x_57140 = x_25852 & x_25853;
assign x_57141 = x_25854 & x_25855;
assign x_57142 = x_57140 & x_57141;
assign x_57143 = x_57139 & x_57142;
assign x_57144 = x_57136 & x_57143;
assign x_57145 = x_57129 & x_57144;
assign x_57146 = x_57115 & x_57145;
assign x_57147 = x_25857 & x_25858;
assign x_57148 = x_25856 & x_57147;
assign x_57149 = x_25859 & x_25860;
assign x_57150 = x_25861 & x_25862;
assign x_57151 = x_57149 & x_57150;
assign x_57152 = x_57148 & x_57151;
assign x_57153 = x_25863 & x_25864;
assign x_57154 = x_25865 & x_25866;
assign x_57155 = x_57153 & x_57154;
assign x_57156 = x_25867 & x_25868;
assign x_57157 = x_25869 & x_25870;
assign x_57158 = x_57156 & x_57157;
assign x_57159 = x_57155 & x_57158;
assign x_57160 = x_57152 & x_57159;
assign x_57161 = x_25871 & x_25872;
assign x_57162 = x_25873 & x_25874;
assign x_57163 = x_57161 & x_57162;
assign x_57164 = x_25875 & x_25876;
assign x_57165 = x_25877 & x_25878;
assign x_57166 = x_57164 & x_57165;
assign x_57167 = x_57163 & x_57166;
assign x_57168 = x_25879 & x_25880;
assign x_57169 = x_25881 & x_25882;
assign x_57170 = x_57168 & x_57169;
assign x_57171 = x_25883 & x_25884;
assign x_57172 = x_25885 & x_25886;
assign x_57173 = x_57171 & x_57172;
assign x_57174 = x_57170 & x_57173;
assign x_57175 = x_57167 & x_57174;
assign x_57176 = x_57160 & x_57175;
assign x_57177 = x_25888 & x_25889;
assign x_57178 = x_25887 & x_57177;
assign x_57179 = x_25890 & x_25891;
assign x_57180 = x_25892 & x_25893;
assign x_57181 = x_57179 & x_57180;
assign x_57182 = x_57178 & x_57181;
assign x_57183 = x_25894 & x_25895;
assign x_57184 = x_25896 & x_25897;
assign x_57185 = x_57183 & x_57184;
assign x_57186 = x_25898 & x_25899;
assign x_57187 = x_25900 & x_25901;
assign x_57188 = x_57186 & x_57187;
assign x_57189 = x_57185 & x_57188;
assign x_57190 = x_57182 & x_57189;
assign x_57191 = x_25902 & x_25903;
assign x_57192 = x_25904 & x_25905;
assign x_57193 = x_57191 & x_57192;
assign x_57194 = x_25906 & x_25907;
assign x_57195 = x_25908 & x_25909;
assign x_57196 = x_57194 & x_57195;
assign x_57197 = x_57193 & x_57196;
assign x_57198 = x_25910 & x_25911;
assign x_57199 = x_25912 & x_25913;
assign x_57200 = x_57198 & x_57199;
assign x_57201 = x_25914 & x_25915;
assign x_57202 = x_25916 & x_25917;
assign x_57203 = x_57201 & x_57202;
assign x_57204 = x_57200 & x_57203;
assign x_57205 = x_57197 & x_57204;
assign x_57206 = x_57190 & x_57205;
assign x_57207 = x_57176 & x_57206;
assign x_57208 = x_57146 & x_57207;
assign x_57209 = x_57086 & x_57208;
assign x_57210 = x_56965 & x_57209;
assign x_57211 = x_25919 & x_25920;
assign x_57212 = x_25918 & x_57211;
assign x_57213 = x_25921 & x_25922;
assign x_57214 = x_25923 & x_25924;
assign x_57215 = x_57213 & x_57214;
assign x_57216 = x_57212 & x_57215;
assign x_57217 = x_25925 & x_25926;
assign x_57218 = x_25927 & x_25928;
assign x_57219 = x_57217 & x_57218;
assign x_57220 = x_25929 & x_25930;
assign x_57221 = x_25931 & x_25932;
assign x_57222 = x_57220 & x_57221;
assign x_57223 = x_57219 & x_57222;
assign x_57224 = x_57216 & x_57223;
assign x_57225 = x_25934 & x_25935;
assign x_57226 = x_25933 & x_57225;
assign x_57227 = x_25936 & x_25937;
assign x_57228 = x_25938 & x_25939;
assign x_57229 = x_57227 & x_57228;
assign x_57230 = x_57226 & x_57229;
assign x_57231 = x_25940 & x_25941;
assign x_57232 = x_25942 & x_25943;
assign x_57233 = x_57231 & x_57232;
assign x_57234 = x_25944 & x_25945;
assign x_57235 = x_25946 & x_25947;
assign x_57236 = x_57234 & x_57235;
assign x_57237 = x_57233 & x_57236;
assign x_57238 = x_57230 & x_57237;
assign x_57239 = x_57224 & x_57238;
assign x_57240 = x_25949 & x_25950;
assign x_57241 = x_25948 & x_57240;
assign x_57242 = x_25951 & x_25952;
assign x_57243 = x_25953 & x_25954;
assign x_57244 = x_57242 & x_57243;
assign x_57245 = x_57241 & x_57244;
assign x_57246 = x_25955 & x_25956;
assign x_57247 = x_25957 & x_25958;
assign x_57248 = x_57246 & x_57247;
assign x_57249 = x_25959 & x_25960;
assign x_57250 = x_25961 & x_25962;
assign x_57251 = x_57249 & x_57250;
assign x_57252 = x_57248 & x_57251;
assign x_57253 = x_57245 & x_57252;
assign x_57254 = x_25963 & x_25964;
assign x_57255 = x_25965 & x_25966;
assign x_57256 = x_57254 & x_57255;
assign x_57257 = x_25967 & x_25968;
assign x_57258 = x_25969 & x_25970;
assign x_57259 = x_57257 & x_57258;
assign x_57260 = x_57256 & x_57259;
assign x_57261 = x_25971 & x_25972;
assign x_57262 = x_25973 & x_25974;
assign x_57263 = x_57261 & x_57262;
assign x_57264 = x_25975 & x_25976;
assign x_57265 = x_25977 & x_25978;
assign x_57266 = x_57264 & x_57265;
assign x_57267 = x_57263 & x_57266;
assign x_57268 = x_57260 & x_57267;
assign x_57269 = x_57253 & x_57268;
assign x_57270 = x_57239 & x_57269;
assign x_57271 = x_25980 & x_25981;
assign x_57272 = x_25979 & x_57271;
assign x_57273 = x_25982 & x_25983;
assign x_57274 = x_25984 & x_25985;
assign x_57275 = x_57273 & x_57274;
assign x_57276 = x_57272 & x_57275;
assign x_57277 = x_25986 & x_25987;
assign x_57278 = x_25988 & x_25989;
assign x_57279 = x_57277 & x_57278;
assign x_57280 = x_25990 & x_25991;
assign x_57281 = x_25992 & x_25993;
assign x_57282 = x_57280 & x_57281;
assign x_57283 = x_57279 & x_57282;
assign x_57284 = x_57276 & x_57283;
assign x_57285 = x_25995 & x_25996;
assign x_57286 = x_25994 & x_57285;
assign x_57287 = x_25997 & x_25998;
assign x_57288 = x_25999 & x_26000;
assign x_57289 = x_57287 & x_57288;
assign x_57290 = x_57286 & x_57289;
assign x_57291 = x_26001 & x_26002;
assign x_57292 = x_26003 & x_26004;
assign x_57293 = x_57291 & x_57292;
assign x_57294 = x_26005 & x_26006;
assign x_57295 = x_26007 & x_26008;
assign x_57296 = x_57294 & x_57295;
assign x_57297 = x_57293 & x_57296;
assign x_57298 = x_57290 & x_57297;
assign x_57299 = x_57284 & x_57298;
assign x_57300 = x_26010 & x_26011;
assign x_57301 = x_26009 & x_57300;
assign x_57302 = x_26012 & x_26013;
assign x_57303 = x_26014 & x_26015;
assign x_57304 = x_57302 & x_57303;
assign x_57305 = x_57301 & x_57304;
assign x_57306 = x_26016 & x_26017;
assign x_57307 = x_26018 & x_26019;
assign x_57308 = x_57306 & x_57307;
assign x_57309 = x_26020 & x_26021;
assign x_57310 = x_26022 & x_26023;
assign x_57311 = x_57309 & x_57310;
assign x_57312 = x_57308 & x_57311;
assign x_57313 = x_57305 & x_57312;
assign x_57314 = x_26024 & x_26025;
assign x_57315 = x_26026 & x_26027;
assign x_57316 = x_57314 & x_57315;
assign x_57317 = x_26028 & x_26029;
assign x_57318 = x_26030 & x_26031;
assign x_57319 = x_57317 & x_57318;
assign x_57320 = x_57316 & x_57319;
assign x_57321 = x_26032 & x_26033;
assign x_57322 = x_26034 & x_26035;
assign x_57323 = x_57321 & x_57322;
assign x_57324 = x_26036 & x_26037;
assign x_57325 = x_26038 & x_26039;
assign x_57326 = x_57324 & x_57325;
assign x_57327 = x_57323 & x_57326;
assign x_57328 = x_57320 & x_57327;
assign x_57329 = x_57313 & x_57328;
assign x_57330 = x_57299 & x_57329;
assign x_57331 = x_57270 & x_57330;
assign x_57332 = x_26041 & x_26042;
assign x_57333 = x_26040 & x_57332;
assign x_57334 = x_26043 & x_26044;
assign x_57335 = x_26045 & x_26046;
assign x_57336 = x_57334 & x_57335;
assign x_57337 = x_57333 & x_57336;
assign x_57338 = x_26047 & x_26048;
assign x_57339 = x_26049 & x_26050;
assign x_57340 = x_57338 & x_57339;
assign x_57341 = x_26051 & x_26052;
assign x_57342 = x_26053 & x_26054;
assign x_57343 = x_57341 & x_57342;
assign x_57344 = x_57340 & x_57343;
assign x_57345 = x_57337 & x_57344;
assign x_57346 = x_26056 & x_26057;
assign x_57347 = x_26055 & x_57346;
assign x_57348 = x_26058 & x_26059;
assign x_57349 = x_26060 & x_26061;
assign x_57350 = x_57348 & x_57349;
assign x_57351 = x_57347 & x_57350;
assign x_57352 = x_26062 & x_26063;
assign x_57353 = x_26064 & x_26065;
assign x_57354 = x_57352 & x_57353;
assign x_57355 = x_26066 & x_26067;
assign x_57356 = x_26068 & x_26069;
assign x_57357 = x_57355 & x_57356;
assign x_57358 = x_57354 & x_57357;
assign x_57359 = x_57351 & x_57358;
assign x_57360 = x_57345 & x_57359;
assign x_57361 = x_26071 & x_26072;
assign x_57362 = x_26070 & x_57361;
assign x_57363 = x_26073 & x_26074;
assign x_57364 = x_26075 & x_26076;
assign x_57365 = x_57363 & x_57364;
assign x_57366 = x_57362 & x_57365;
assign x_57367 = x_26077 & x_26078;
assign x_57368 = x_26079 & x_26080;
assign x_57369 = x_57367 & x_57368;
assign x_57370 = x_26081 & x_26082;
assign x_57371 = x_26083 & x_26084;
assign x_57372 = x_57370 & x_57371;
assign x_57373 = x_57369 & x_57372;
assign x_57374 = x_57366 & x_57373;
assign x_57375 = x_26085 & x_26086;
assign x_57376 = x_26087 & x_26088;
assign x_57377 = x_57375 & x_57376;
assign x_57378 = x_26089 & x_26090;
assign x_57379 = x_26091 & x_26092;
assign x_57380 = x_57378 & x_57379;
assign x_57381 = x_57377 & x_57380;
assign x_57382 = x_26093 & x_26094;
assign x_57383 = x_26095 & x_26096;
assign x_57384 = x_57382 & x_57383;
assign x_57385 = x_26097 & x_26098;
assign x_57386 = x_26099 & x_26100;
assign x_57387 = x_57385 & x_57386;
assign x_57388 = x_57384 & x_57387;
assign x_57389 = x_57381 & x_57388;
assign x_57390 = x_57374 & x_57389;
assign x_57391 = x_57360 & x_57390;
assign x_57392 = x_26102 & x_26103;
assign x_57393 = x_26101 & x_57392;
assign x_57394 = x_26104 & x_26105;
assign x_57395 = x_26106 & x_26107;
assign x_57396 = x_57394 & x_57395;
assign x_57397 = x_57393 & x_57396;
assign x_57398 = x_26108 & x_26109;
assign x_57399 = x_26110 & x_26111;
assign x_57400 = x_57398 & x_57399;
assign x_57401 = x_26112 & x_26113;
assign x_57402 = x_26114 & x_26115;
assign x_57403 = x_57401 & x_57402;
assign x_57404 = x_57400 & x_57403;
assign x_57405 = x_57397 & x_57404;
assign x_57406 = x_26117 & x_26118;
assign x_57407 = x_26116 & x_57406;
assign x_57408 = x_26119 & x_26120;
assign x_57409 = x_26121 & x_26122;
assign x_57410 = x_57408 & x_57409;
assign x_57411 = x_57407 & x_57410;
assign x_57412 = x_26123 & x_26124;
assign x_57413 = x_26125 & x_26126;
assign x_57414 = x_57412 & x_57413;
assign x_57415 = x_26127 & x_26128;
assign x_57416 = x_26129 & x_26130;
assign x_57417 = x_57415 & x_57416;
assign x_57418 = x_57414 & x_57417;
assign x_57419 = x_57411 & x_57418;
assign x_57420 = x_57405 & x_57419;
assign x_57421 = x_26132 & x_26133;
assign x_57422 = x_26131 & x_57421;
assign x_57423 = x_26134 & x_26135;
assign x_57424 = x_26136 & x_26137;
assign x_57425 = x_57423 & x_57424;
assign x_57426 = x_57422 & x_57425;
assign x_57427 = x_26138 & x_26139;
assign x_57428 = x_26140 & x_26141;
assign x_57429 = x_57427 & x_57428;
assign x_57430 = x_26142 & x_26143;
assign x_57431 = x_26144 & x_26145;
assign x_57432 = x_57430 & x_57431;
assign x_57433 = x_57429 & x_57432;
assign x_57434 = x_57426 & x_57433;
assign x_57435 = x_26146 & x_26147;
assign x_57436 = x_26148 & x_26149;
assign x_57437 = x_57435 & x_57436;
assign x_57438 = x_26150 & x_26151;
assign x_57439 = x_26152 & x_26153;
assign x_57440 = x_57438 & x_57439;
assign x_57441 = x_57437 & x_57440;
assign x_57442 = x_26154 & x_26155;
assign x_57443 = x_26156 & x_26157;
assign x_57444 = x_57442 & x_57443;
assign x_57445 = x_26158 & x_26159;
assign x_57446 = x_26160 & x_26161;
assign x_57447 = x_57445 & x_57446;
assign x_57448 = x_57444 & x_57447;
assign x_57449 = x_57441 & x_57448;
assign x_57450 = x_57434 & x_57449;
assign x_57451 = x_57420 & x_57450;
assign x_57452 = x_57391 & x_57451;
assign x_57453 = x_57331 & x_57452;
assign x_57454 = x_26163 & x_26164;
assign x_57455 = x_26162 & x_57454;
assign x_57456 = x_26165 & x_26166;
assign x_57457 = x_26167 & x_26168;
assign x_57458 = x_57456 & x_57457;
assign x_57459 = x_57455 & x_57458;
assign x_57460 = x_26169 & x_26170;
assign x_57461 = x_26171 & x_26172;
assign x_57462 = x_57460 & x_57461;
assign x_57463 = x_26173 & x_26174;
assign x_57464 = x_26175 & x_26176;
assign x_57465 = x_57463 & x_57464;
assign x_57466 = x_57462 & x_57465;
assign x_57467 = x_57459 & x_57466;
assign x_57468 = x_26178 & x_26179;
assign x_57469 = x_26177 & x_57468;
assign x_57470 = x_26180 & x_26181;
assign x_57471 = x_26182 & x_26183;
assign x_57472 = x_57470 & x_57471;
assign x_57473 = x_57469 & x_57472;
assign x_57474 = x_26184 & x_26185;
assign x_57475 = x_26186 & x_26187;
assign x_57476 = x_57474 & x_57475;
assign x_57477 = x_26188 & x_26189;
assign x_57478 = x_26190 & x_26191;
assign x_57479 = x_57477 & x_57478;
assign x_57480 = x_57476 & x_57479;
assign x_57481 = x_57473 & x_57480;
assign x_57482 = x_57467 & x_57481;
assign x_57483 = x_26193 & x_26194;
assign x_57484 = x_26192 & x_57483;
assign x_57485 = x_26195 & x_26196;
assign x_57486 = x_26197 & x_26198;
assign x_57487 = x_57485 & x_57486;
assign x_57488 = x_57484 & x_57487;
assign x_57489 = x_26199 & x_26200;
assign x_57490 = x_26201 & x_26202;
assign x_57491 = x_57489 & x_57490;
assign x_57492 = x_26203 & x_26204;
assign x_57493 = x_26205 & x_26206;
assign x_57494 = x_57492 & x_57493;
assign x_57495 = x_57491 & x_57494;
assign x_57496 = x_57488 & x_57495;
assign x_57497 = x_26207 & x_26208;
assign x_57498 = x_26209 & x_26210;
assign x_57499 = x_57497 & x_57498;
assign x_57500 = x_26211 & x_26212;
assign x_57501 = x_26213 & x_26214;
assign x_57502 = x_57500 & x_57501;
assign x_57503 = x_57499 & x_57502;
assign x_57504 = x_26215 & x_26216;
assign x_57505 = x_26217 & x_26218;
assign x_57506 = x_57504 & x_57505;
assign x_57507 = x_26219 & x_26220;
assign x_57508 = x_26221 & x_26222;
assign x_57509 = x_57507 & x_57508;
assign x_57510 = x_57506 & x_57509;
assign x_57511 = x_57503 & x_57510;
assign x_57512 = x_57496 & x_57511;
assign x_57513 = x_57482 & x_57512;
assign x_57514 = x_26224 & x_26225;
assign x_57515 = x_26223 & x_57514;
assign x_57516 = x_26226 & x_26227;
assign x_57517 = x_26228 & x_26229;
assign x_57518 = x_57516 & x_57517;
assign x_57519 = x_57515 & x_57518;
assign x_57520 = x_26230 & x_26231;
assign x_57521 = x_26232 & x_26233;
assign x_57522 = x_57520 & x_57521;
assign x_57523 = x_26234 & x_26235;
assign x_57524 = x_26236 & x_26237;
assign x_57525 = x_57523 & x_57524;
assign x_57526 = x_57522 & x_57525;
assign x_57527 = x_57519 & x_57526;
assign x_57528 = x_26239 & x_26240;
assign x_57529 = x_26238 & x_57528;
assign x_57530 = x_26241 & x_26242;
assign x_57531 = x_26243 & x_26244;
assign x_57532 = x_57530 & x_57531;
assign x_57533 = x_57529 & x_57532;
assign x_57534 = x_26245 & x_26246;
assign x_57535 = x_26247 & x_26248;
assign x_57536 = x_57534 & x_57535;
assign x_57537 = x_26249 & x_26250;
assign x_57538 = x_26251 & x_26252;
assign x_57539 = x_57537 & x_57538;
assign x_57540 = x_57536 & x_57539;
assign x_57541 = x_57533 & x_57540;
assign x_57542 = x_57527 & x_57541;
assign x_57543 = x_26254 & x_26255;
assign x_57544 = x_26253 & x_57543;
assign x_57545 = x_26256 & x_26257;
assign x_57546 = x_26258 & x_26259;
assign x_57547 = x_57545 & x_57546;
assign x_57548 = x_57544 & x_57547;
assign x_57549 = x_26260 & x_26261;
assign x_57550 = x_26262 & x_26263;
assign x_57551 = x_57549 & x_57550;
assign x_57552 = x_26264 & x_26265;
assign x_57553 = x_26266 & x_26267;
assign x_57554 = x_57552 & x_57553;
assign x_57555 = x_57551 & x_57554;
assign x_57556 = x_57548 & x_57555;
assign x_57557 = x_26268 & x_26269;
assign x_57558 = x_26270 & x_26271;
assign x_57559 = x_57557 & x_57558;
assign x_57560 = x_26272 & x_26273;
assign x_57561 = x_26274 & x_26275;
assign x_57562 = x_57560 & x_57561;
assign x_57563 = x_57559 & x_57562;
assign x_57564 = x_26276 & x_26277;
assign x_57565 = x_26278 & x_26279;
assign x_57566 = x_57564 & x_57565;
assign x_57567 = x_26280 & x_26281;
assign x_57568 = x_26282 & x_26283;
assign x_57569 = x_57567 & x_57568;
assign x_57570 = x_57566 & x_57569;
assign x_57571 = x_57563 & x_57570;
assign x_57572 = x_57556 & x_57571;
assign x_57573 = x_57542 & x_57572;
assign x_57574 = x_57513 & x_57573;
assign x_57575 = x_26285 & x_26286;
assign x_57576 = x_26284 & x_57575;
assign x_57577 = x_26287 & x_26288;
assign x_57578 = x_26289 & x_26290;
assign x_57579 = x_57577 & x_57578;
assign x_57580 = x_57576 & x_57579;
assign x_57581 = x_26291 & x_26292;
assign x_57582 = x_26293 & x_26294;
assign x_57583 = x_57581 & x_57582;
assign x_57584 = x_26295 & x_26296;
assign x_57585 = x_26297 & x_26298;
assign x_57586 = x_57584 & x_57585;
assign x_57587 = x_57583 & x_57586;
assign x_57588 = x_57580 & x_57587;
assign x_57589 = x_26300 & x_26301;
assign x_57590 = x_26299 & x_57589;
assign x_57591 = x_26302 & x_26303;
assign x_57592 = x_26304 & x_26305;
assign x_57593 = x_57591 & x_57592;
assign x_57594 = x_57590 & x_57593;
assign x_57595 = x_26306 & x_26307;
assign x_57596 = x_26308 & x_26309;
assign x_57597 = x_57595 & x_57596;
assign x_57598 = x_26310 & x_26311;
assign x_57599 = x_26312 & x_26313;
assign x_57600 = x_57598 & x_57599;
assign x_57601 = x_57597 & x_57600;
assign x_57602 = x_57594 & x_57601;
assign x_57603 = x_57588 & x_57602;
assign x_57604 = x_26315 & x_26316;
assign x_57605 = x_26314 & x_57604;
assign x_57606 = x_26317 & x_26318;
assign x_57607 = x_26319 & x_26320;
assign x_57608 = x_57606 & x_57607;
assign x_57609 = x_57605 & x_57608;
assign x_57610 = x_26321 & x_26322;
assign x_57611 = x_26323 & x_26324;
assign x_57612 = x_57610 & x_57611;
assign x_57613 = x_26325 & x_26326;
assign x_57614 = x_26327 & x_26328;
assign x_57615 = x_57613 & x_57614;
assign x_57616 = x_57612 & x_57615;
assign x_57617 = x_57609 & x_57616;
assign x_57618 = x_26329 & x_26330;
assign x_57619 = x_26331 & x_26332;
assign x_57620 = x_57618 & x_57619;
assign x_57621 = x_26333 & x_26334;
assign x_57622 = x_26335 & x_26336;
assign x_57623 = x_57621 & x_57622;
assign x_57624 = x_57620 & x_57623;
assign x_57625 = x_26337 & x_26338;
assign x_57626 = x_26339 & x_26340;
assign x_57627 = x_57625 & x_57626;
assign x_57628 = x_26341 & x_26342;
assign x_57629 = x_26343 & x_26344;
assign x_57630 = x_57628 & x_57629;
assign x_57631 = x_57627 & x_57630;
assign x_57632 = x_57624 & x_57631;
assign x_57633 = x_57617 & x_57632;
assign x_57634 = x_57603 & x_57633;
assign x_57635 = x_26346 & x_26347;
assign x_57636 = x_26345 & x_57635;
assign x_57637 = x_26348 & x_26349;
assign x_57638 = x_26350 & x_26351;
assign x_57639 = x_57637 & x_57638;
assign x_57640 = x_57636 & x_57639;
assign x_57641 = x_26352 & x_26353;
assign x_57642 = x_26354 & x_26355;
assign x_57643 = x_57641 & x_57642;
assign x_57644 = x_26356 & x_26357;
assign x_57645 = x_26358 & x_26359;
assign x_57646 = x_57644 & x_57645;
assign x_57647 = x_57643 & x_57646;
assign x_57648 = x_57640 & x_57647;
assign x_57649 = x_26360 & x_26361;
assign x_57650 = x_26362 & x_26363;
assign x_57651 = x_57649 & x_57650;
assign x_57652 = x_26364 & x_26365;
assign x_57653 = x_26366 & x_26367;
assign x_57654 = x_57652 & x_57653;
assign x_57655 = x_57651 & x_57654;
assign x_57656 = x_26368 & x_26369;
assign x_57657 = x_26370 & x_26371;
assign x_57658 = x_57656 & x_57657;
assign x_57659 = x_26372 & x_26373;
assign x_57660 = x_26374 & x_26375;
assign x_57661 = x_57659 & x_57660;
assign x_57662 = x_57658 & x_57661;
assign x_57663 = x_57655 & x_57662;
assign x_57664 = x_57648 & x_57663;
assign x_57665 = x_26377 & x_26378;
assign x_57666 = x_26376 & x_57665;
assign x_57667 = x_26379 & x_26380;
assign x_57668 = x_26381 & x_26382;
assign x_57669 = x_57667 & x_57668;
assign x_57670 = x_57666 & x_57669;
assign x_57671 = x_26383 & x_26384;
assign x_57672 = x_26385 & x_26386;
assign x_57673 = x_57671 & x_57672;
assign x_57674 = x_26387 & x_26388;
assign x_57675 = x_26389 & x_26390;
assign x_57676 = x_57674 & x_57675;
assign x_57677 = x_57673 & x_57676;
assign x_57678 = x_57670 & x_57677;
assign x_57679 = x_26391 & x_26392;
assign x_57680 = x_26393 & x_26394;
assign x_57681 = x_57679 & x_57680;
assign x_57682 = x_26395 & x_26396;
assign x_57683 = x_26397 & x_26398;
assign x_57684 = x_57682 & x_57683;
assign x_57685 = x_57681 & x_57684;
assign x_57686 = x_26399 & x_26400;
assign x_57687 = x_26401 & x_26402;
assign x_57688 = x_57686 & x_57687;
assign x_57689 = x_26403 & x_26404;
assign x_57690 = x_26405 & x_26406;
assign x_57691 = x_57689 & x_57690;
assign x_57692 = x_57688 & x_57691;
assign x_57693 = x_57685 & x_57692;
assign x_57694 = x_57678 & x_57693;
assign x_57695 = x_57664 & x_57694;
assign x_57696 = x_57634 & x_57695;
assign x_57697 = x_57574 & x_57696;
assign x_57698 = x_57453 & x_57697;
assign x_57699 = x_57210 & x_57698;
assign x_57700 = x_26408 & x_26409;
assign x_57701 = x_26407 & x_57700;
assign x_57702 = x_26410 & x_26411;
assign x_57703 = x_26412 & x_26413;
assign x_57704 = x_57702 & x_57703;
assign x_57705 = x_57701 & x_57704;
assign x_57706 = x_26414 & x_26415;
assign x_57707 = x_26416 & x_26417;
assign x_57708 = x_57706 & x_57707;
assign x_57709 = x_26418 & x_26419;
assign x_57710 = x_26420 & x_26421;
assign x_57711 = x_57709 & x_57710;
assign x_57712 = x_57708 & x_57711;
assign x_57713 = x_57705 & x_57712;
assign x_57714 = x_26423 & x_26424;
assign x_57715 = x_26422 & x_57714;
assign x_57716 = x_26425 & x_26426;
assign x_57717 = x_26427 & x_26428;
assign x_57718 = x_57716 & x_57717;
assign x_57719 = x_57715 & x_57718;
assign x_57720 = x_26429 & x_26430;
assign x_57721 = x_26431 & x_26432;
assign x_57722 = x_57720 & x_57721;
assign x_57723 = x_26433 & x_26434;
assign x_57724 = x_26435 & x_26436;
assign x_57725 = x_57723 & x_57724;
assign x_57726 = x_57722 & x_57725;
assign x_57727 = x_57719 & x_57726;
assign x_57728 = x_57713 & x_57727;
assign x_57729 = x_26438 & x_26439;
assign x_57730 = x_26437 & x_57729;
assign x_57731 = x_26440 & x_26441;
assign x_57732 = x_26442 & x_26443;
assign x_57733 = x_57731 & x_57732;
assign x_57734 = x_57730 & x_57733;
assign x_57735 = x_26444 & x_26445;
assign x_57736 = x_26446 & x_26447;
assign x_57737 = x_57735 & x_57736;
assign x_57738 = x_26448 & x_26449;
assign x_57739 = x_26450 & x_26451;
assign x_57740 = x_57738 & x_57739;
assign x_57741 = x_57737 & x_57740;
assign x_57742 = x_57734 & x_57741;
assign x_57743 = x_26452 & x_26453;
assign x_57744 = x_26454 & x_26455;
assign x_57745 = x_57743 & x_57744;
assign x_57746 = x_26456 & x_26457;
assign x_57747 = x_26458 & x_26459;
assign x_57748 = x_57746 & x_57747;
assign x_57749 = x_57745 & x_57748;
assign x_57750 = x_26460 & x_26461;
assign x_57751 = x_26462 & x_26463;
assign x_57752 = x_57750 & x_57751;
assign x_57753 = x_26464 & x_26465;
assign x_57754 = x_26466 & x_26467;
assign x_57755 = x_57753 & x_57754;
assign x_57756 = x_57752 & x_57755;
assign x_57757 = x_57749 & x_57756;
assign x_57758 = x_57742 & x_57757;
assign x_57759 = x_57728 & x_57758;
assign x_57760 = x_26469 & x_26470;
assign x_57761 = x_26468 & x_57760;
assign x_57762 = x_26471 & x_26472;
assign x_57763 = x_26473 & x_26474;
assign x_57764 = x_57762 & x_57763;
assign x_57765 = x_57761 & x_57764;
assign x_57766 = x_26475 & x_26476;
assign x_57767 = x_26477 & x_26478;
assign x_57768 = x_57766 & x_57767;
assign x_57769 = x_26479 & x_26480;
assign x_57770 = x_26481 & x_26482;
assign x_57771 = x_57769 & x_57770;
assign x_57772 = x_57768 & x_57771;
assign x_57773 = x_57765 & x_57772;
assign x_57774 = x_26484 & x_26485;
assign x_57775 = x_26483 & x_57774;
assign x_57776 = x_26486 & x_26487;
assign x_57777 = x_26488 & x_26489;
assign x_57778 = x_57776 & x_57777;
assign x_57779 = x_57775 & x_57778;
assign x_57780 = x_26490 & x_26491;
assign x_57781 = x_26492 & x_26493;
assign x_57782 = x_57780 & x_57781;
assign x_57783 = x_26494 & x_26495;
assign x_57784 = x_26496 & x_26497;
assign x_57785 = x_57783 & x_57784;
assign x_57786 = x_57782 & x_57785;
assign x_57787 = x_57779 & x_57786;
assign x_57788 = x_57773 & x_57787;
assign x_57789 = x_26499 & x_26500;
assign x_57790 = x_26498 & x_57789;
assign x_57791 = x_26501 & x_26502;
assign x_57792 = x_26503 & x_26504;
assign x_57793 = x_57791 & x_57792;
assign x_57794 = x_57790 & x_57793;
assign x_57795 = x_26505 & x_26506;
assign x_57796 = x_26507 & x_26508;
assign x_57797 = x_57795 & x_57796;
assign x_57798 = x_26509 & x_26510;
assign x_57799 = x_26511 & x_26512;
assign x_57800 = x_57798 & x_57799;
assign x_57801 = x_57797 & x_57800;
assign x_57802 = x_57794 & x_57801;
assign x_57803 = x_26513 & x_26514;
assign x_57804 = x_26515 & x_26516;
assign x_57805 = x_57803 & x_57804;
assign x_57806 = x_26517 & x_26518;
assign x_57807 = x_26519 & x_26520;
assign x_57808 = x_57806 & x_57807;
assign x_57809 = x_57805 & x_57808;
assign x_57810 = x_26521 & x_26522;
assign x_57811 = x_26523 & x_26524;
assign x_57812 = x_57810 & x_57811;
assign x_57813 = x_26525 & x_26526;
assign x_57814 = x_26527 & x_26528;
assign x_57815 = x_57813 & x_57814;
assign x_57816 = x_57812 & x_57815;
assign x_57817 = x_57809 & x_57816;
assign x_57818 = x_57802 & x_57817;
assign x_57819 = x_57788 & x_57818;
assign x_57820 = x_57759 & x_57819;
assign x_57821 = x_26530 & x_26531;
assign x_57822 = x_26529 & x_57821;
assign x_57823 = x_26532 & x_26533;
assign x_57824 = x_26534 & x_26535;
assign x_57825 = x_57823 & x_57824;
assign x_57826 = x_57822 & x_57825;
assign x_57827 = x_26536 & x_26537;
assign x_57828 = x_26538 & x_26539;
assign x_57829 = x_57827 & x_57828;
assign x_57830 = x_26540 & x_26541;
assign x_57831 = x_26542 & x_26543;
assign x_57832 = x_57830 & x_57831;
assign x_57833 = x_57829 & x_57832;
assign x_57834 = x_57826 & x_57833;
assign x_57835 = x_26545 & x_26546;
assign x_57836 = x_26544 & x_57835;
assign x_57837 = x_26547 & x_26548;
assign x_57838 = x_26549 & x_26550;
assign x_57839 = x_57837 & x_57838;
assign x_57840 = x_57836 & x_57839;
assign x_57841 = x_26551 & x_26552;
assign x_57842 = x_26553 & x_26554;
assign x_57843 = x_57841 & x_57842;
assign x_57844 = x_26555 & x_26556;
assign x_57845 = x_26557 & x_26558;
assign x_57846 = x_57844 & x_57845;
assign x_57847 = x_57843 & x_57846;
assign x_57848 = x_57840 & x_57847;
assign x_57849 = x_57834 & x_57848;
assign x_57850 = x_26560 & x_26561;
assign x_57851 = x_26559 & x_57850;
assign x_57852 = x_26562 & x_26563;
assign x_57853 = x_26564 & x_26565;
assign x_57854 = x_57852 & x_57853;
assign x_57855 = x_57851 & x_57854;
assign x_57856 = x_26566 & x_26567;
assign x_57857 = x_26568 & x_26569;
assign x_57858 = x_57856 & x_57857;
assign x_57859 = x_26570 & x_26571;
assign x_57860 = x_26572 & x_26573;
assign x_57861 = x_57859 & x_57860;
assign x_57862 = x_57858 & x_57861;
assign x_57863 = x_57855 & x_57862;
assign x_57864 = x_26574 & x_26575;
assign x_57865 = x_26576 & x_26577;
assign x_57866 = x_57864 & x_57865;
assign x_57867 = x_26578 & x_26579;
assign x_57868 = x_26580 & x_26581;
assign x_57869 = x_57867 & x_57868;
assign x_57870 = x_57866 & x_57869;
assign x_57871 = x_26582 & x_26583;
assign x_57872 = x_26584 & x_26585;
assign x_57873 = x_57871 & x_57872;
assign x_57874 = x_26586 & x_26587;
assign x_57875 = x_26588 & x_26589;
assign x_57876 = x_57874 & x_57875;
assign x_57877 = x_57873 & x_57876;
assign x_57878 = x_57870 & x_57877;
assign x_57879 = x_57863 & x_57878;
assign x_57880 = x_57849 & x_57879;
assign x_57881 = x_26591 & x_26592;
assign x_57882 = x_26590 & x_57881;
assign x_57883 = x_26593 & x_26594;
assign x_57884 = x_26595 & x_26596;
assign x_57885 = x_57883 & x_57884;
assign x_57886 = x_57882 & x_57885;
assign x_57887 = x_26597 & x_26598;
assign x_57888 = x_26599 & x_26600;
assign x_57889 = x_57887 & x_57888;
assign x_57890 = x_26601 & x_26602;
assign x_57891 = x_26603 & x_26604;
assign x_57892 = x_57890 & x_57891;
assign x_57893 = x_57889 & x_57892;
assign x_57894 = x_57886 & x_57893;
assign x_57895 = x_26606 & x_26607;
assign x_57896 = x_26605 & x_57895;
assign x_57897 = x_26608 & x_26609;
assign x_57898 = x_26610 & x_26611;
assign x_57899 = x_57897 & x_57898;
assign x_57900 = x_57896 & x_57899;
assign x_57901 = x_26612 & x_26613;
assign x_57902 = x_26614 & x_26615;
assign x_57903 = x_57901 & x_57902;
assign x_57904 = x_26616 & x_26617;
assign x_57905 = x_26618 & x_26619;
assign x_57906 = x_57904 & x_57905;
assign x_57907 = x_57903 & x_57906;
assign x_57908 = x_57900 & x_57907;
assign x_57909 = x_57894 & x_57908;
assign x_57910 = x_26621 & x_26622;
assign x_57911 = x_26620 & x_57910;
assign x_57912 = x_26623 & x_26624;
assign x_57913 = x_26625 & x_26626;
assign x_57914 = x_57912 & x_57913;
assign x_57915 = x_57911 & x_57914;
assign x_57916 = x_26627 & x_26628;
assign x_57917 = x_26629 & x_26630;
assign x_57918 = x_57916 & x_57917;
assign x_57919 = x_26631 & x_26632;
assign x_57920 = x_26633 & x_26634;
assign x_57921 = x_57919 & x_57920;
assign x_57922 = x_57918 & x_57921;
assign x_57923 = x_57915 & x_57922;
assign x_57924 = x_26635 & x_26636;
assign x_57925 = x_26637 & x_26638;
assign x_57926 = x_57924 & x_57925;
assign x_57927 = x_26639 & x_26640;
assign x_57928 = x_26641 & x_26642;
assign x_57929 = x_57927 & x_57928;
assign x_57930 = x_57926 & x_57929;
assign x_57931 = x_26643 & x_26644;
assign x_57932 = x_26645 & x_26646;
assign x_57933 = x_57931 & x_57932;
assign x_57934 = x_26647 & x_26648;
assign x_57935 = x_26649 & x_26650;
assign x_57936 = x_57934 & x_57935;
assign x_57937 = x_57933 & x_57936;
assign x_57938 = x_57930 & x_57937;
assign x_57939 = x_57923 & x_57938;
assign x_57940 = x_57909 & x_57939;
assign x_57941 = x_57880 & x_57940;
assign x_57942 = x_57820 & x_57941;
assign x_57943 = x_26652 & x_26653;
assign x_57944 = x_26651 & x_57943;
assign x_57945 = x_26654 & x_26655;
assign x_57946 = x_26656 & x_26657;
assign x_57947 = x_57945 & x_57946;
assign x_57948 = x_57944 & x_57947;
assign x_57949 = x_26658 & x_26659;
assign x_57950 = x_26660 & x_26661;
assign x_57951 = x_57949 & x_57950;
assign x_57952 = x_26662 & x_26663;
assign x_57953 = x_26664 & x_26665;
assign x_57954 = x_57952 & x_57953;
assign x_57955 = x_57951 & x_57954;
assign x_57956 = x_57948 & x_57955;
assign x_57957 = x_26667 & x_26668;
assign x_57958 = x_26666 & x_57957;
assign x_57959 = x_26669 & x_26670;
assign x_57960 = x_26671 & x_26672;
assign x_57961 = x_57959 & x_57960;
assign x_57962 = x_57958 & x_57961;
assign x_57963 = x_26673 & x_26674;
assign x_57964 = x_26675 & x_26676;
assign x_57965 = x_57963 & x_57964;
assign x_57966 = x_26677 & x_26678;
assign x_57967 = x_26679 & x_26680;
assign x_57968 = x_57966 & x_57967;
assign x_57969 = x_57965 & x_57968;
assign x_57970 = x_57962 & x_57969;
assign x_57971 = x_57956 & x_57970;
assign x_57972 = x_26682 & x_26683;
assign x_57973 = x_26681 & x_57972;
assign x_57974 = x_26684 & x_26685;
assign x_57975 = x_26686 & x_26687;
assign x_57976 = x_57974 & x_57975;
assign x_57977 = x_57973 & x_57976;
assign x_57978 = x_26688 & x_26689;
assign x_57979 = x_26690 & x_26691;
assign x_57980 = x_57978 & x_57979;
assign x_57981 = x_26692 & x_26693;
assign x_57982 = x_26694 & x_26695;
assign x_57983 = x_57981 & x_57982;
assign x_57984 = x_57980 & x_57983;
assign x_57985 = x_57977 & x_57984;
assign x_57986 = x_26696 & x_26697;
assign x_57987 = x_26698 & x_26699;
assign x_57988 = x_57986 & x_57987;
assign x_57989 = x_26700 & x_26701;
assign x_57990 = x_26702 & x_26703;
assign x_57991 = x_57989 & x_57990;
assign x_57992 = x_57988 & x_57991;
assign x_57993 = x_26704 & x_26705;
assign x_57994 = x_26706 & x_26707;
assign x_57995 = x_57993 & x_57994;
assign x_57996 = x_26708 & x_26709;
assign x_57997 = x_26710 & x_26711;
assign x_57998 = x_57996 & x_57997;
assign x_57999 = x_57995 & x_57998;
assign x_58000 = x_57992 & x_57999;
assign x_58001 = x_57985 & x_58000;
assign x_58002 = x_57971 & x_58001;
assign x_58003 = x_26713 & x_26714;
assign x_58004 = x_26712 & x_58003;
assign x_58005 = x_26715 & x_26716;
assign x_58006 = x_26717 & x_26718;
assign x_58007 = x_58005 & x_58006;
assign x_58008 = x_58004 & x_58007;
assign x_58009 = x_26719 & x_26720;
assign x_58010 = x_26721 & x_26722;
assign x_58011 = x_58009 & x_58010;
assign x_58012 = x_26723 & x_26724;
assign x_58013 = x_26725 & x_26726;
assign x_58014 = x_58012 & x_58013;
assign x_58015 = x_58011 & x_58014;
assign x_58016 = x_58008 & x_58015;
assign x_58017 = x_26728 & x_26729;
assign x_58018 = x_26727 & x_58017;
assign x_58019 = x_26730 & x_26731;
assign x_58020 = x_26732 & x_26733;
assign x_58021 = x_58019 & x_58020;
assign x_58022 = x_58018 & x_58021;
assign x_58023 = x_26734 & x_26735;
assign x_58024 = x_26736 & x_26737;
assign x_58025 = x_58023 & x_58024;
assign x_58026 = x_26738 & x_26739;
assign x_58027 = x_26740 & x_26741;
assign x_58028 = x_58026 & x_58027;
assign x_58029 = x_58025 & x_58028;
assign x_58030 = x_58022 & x_58029;
assign x_58031 = x_58016 & x_58030;
assign x_58032 = x_26743 & x_26744;
assign x_58033 = x_26742 & x_58032;
assign x_58034 = x_26745 & x_26746;
assign x_58035 = x_26747 & x_26748;
assign x_58036 = x_58034 & x_58035;
assign x_58037 = x_58033 & x_58036;
assign x_58038 = x_26749 & x_26750;
assign x_58039 = x_26751 & x_26752;
assign x_58040 = x_58038 & x_58039;
assign x_58041 = x_26753 & x_26754;
assign x_58042 = x_26755 & x_26756;
assign x_58043 = x_58041 & x_58042;
assign x_58044 = x_58040 & x_58043;
assign x_58045 = x_58037 & x_58044;
assign x_58046 = x_26757 & x_26758;
assign x_58047 = x_26759 & x_26760;
assign x_58048 = x_58046 & x_58047;
assign x_58049 = x_26761 & x_26762;
assign x_58050 = x_26763 & x_26764;
assign x_58051 = x_58049 & x_58050;
assign x_58052 = x_58048 & x_58051;
assign x_58053 = x_26765 & x_26766;
assign x_58054 = x_26767 & x_26768;
assign x_58055 = x_58053 & x_58054;
assign x_58056 = x_26769 & x_26770;
assign x_58057 = x_26771 & x_26772;
assign x_58058 = x_58056 & x_58057;
assign x_58059 = x_58055 & x_58058;
assign x_58060 = x_58052 & x_58059;
assign x_58061 = x_58045 & x_58060;
assign x_58062 = x_58031 & x_58061;
assign x_58063 = x_58002 & x_58062;
assign x_58064 = x_26774 & x_26775;
assign x_58065 = x_26773 & x_58064;
assign x_58066 = x_26776 & x_26777;
assign x_58067 = x_26778 & x_26779;
assign x_58068 = x_58066 & x_58067;
assign x_58069 = x_58065 & x_58068;
assign x_58070 = x_26780 & x_26781;
assign x_58071 = x_26782 & x_26783;
assign x_58072 = x_58070 & x_58071;
assign x_58073 = x_26784 & x_26785;
assign x_58074 = x_26786 & x_26787;
assign x_58075 = x_58073 & x_58074;
assign x_58076 = x_58072 & x_58075;
assign x_58077 = x_58069 & x_58076;
assign x_58078 = x_26789 & x_26790;
assign x_58079 = x_26788 & x_58078;
assign x_58080 = x_26791 & x_26792;
assign x_58081 = x_26793 & x_26794;
assign x_58082 = x_58080 & x_58081;
assign x_58083 = x_58079 & x_58082;
assign x_58084 = x_26795 & x_26796;
assign x_58085 = x_26797 & x_26798;
assign x_58086 = x_58084 & x_58085;
assign x_58087 = x_26799 & x_26800;
assign x_58088 = x_26801 & x_26802;
assign x_58089 = x_58087 & x_58088;
assign x_58090 = x_58086 & x_58089;
assign x_58091 = x_58083 & x_58090;
assign x_58092 = x_58077 & x_58091;
assign x_58093 = x_26804 & x_26805;
assign x_58094 = x_26803 & x_58093;
assign x_58095 = x_26806 & x_26807;
assign x_58096 = x_26808 & x_26809;
assign x_58097 = x_58095 & x_58096;
assign x_58098 = x_58094 & x_58097;
assign x_58099 = x_26810 & x_26811;
assign x_58100 = x_26812 & x_26813;
assign x_58101 = x_58099 & x_58100;
assign x_58102 = x_26814 & x_26815;
assign x_58103 = x_26816 & x_26817;
assign x_58104 = x_58102 & x_58103;
assign x_58105 = x_58101 & x_58104;
assign x_58106 = x_58098 & x_58105;
assign x_58107 = x_26818 & x_26819;
assign x_58108 = x_26820 & x_26821;
assign x_58109 = x_58107 & x_58108;
assign x_58110 = x_26822 & x_26823;
assign x_58111 = x_26824 & x_26825;
assign x_58112 = x_58110 & x_58111;
assign x_58113 = x_58109 & x_58112;
assign x_58114 = x_26826 & x_26827;
assign x_58115 = x_26828 & x_26829;
assign x_58116 = x_58114 & x_58115;
assign x_58117 = x_26830 & x_26831;
assign x_58118 = x_26832 & x_26833;
assign x_58119 = x_58117 & x_58118;
assign x_58120 = x_58116 & x_58119;
assign x_58121 = x_58113 & x_58120;
assign x_58122 = x_58106 & x_58121;
assign x_58123 = x_58092 & x_58122;
assign x_58124 = x_26835 & x_26836;
assign x_58125 = x_26834 & x_58124;
assign x_58126 = x_26837 & x_26838;
assign x_58127 = x_26839 & x_26840;
assign x_58128 = x_58126 & x_58127;
assign x_58129 = x_58125 & x_58128;
assign x_58130 = x_26841 & x_26842;
assign x_58131 = x_26843 & x_26844;
assign x_58132 = x_58130 & x_58131;
assign x_58133 = x_26845 & x_26846;
assign x_58134 = x_26847 & x_26848;
assign x_58135 = x_58133 & x_58134;
assign x_58136 = x_58132 & x_58135;
assign x_58137 = x_58129 & x_58136;
assign x_58138 = x_26849 & x_26850;
assign x_58139 = x_26851 & x_26852;
assign x_58140 = x_58138 & x_58139;
assign x_58141 = x_26853 & x_26854;
assign x_58142 = x_26855 & x_26856;
assign x_58143 = x_58141 & x_58142;
assign x_58144 = x_58140 & x_58143;
assign x_58145 = x_26857 & x_26858;
assign x_58146 = x_26859 & x_26860;
assign x_58147 = x_58145 & x_58146;
assign x_58148 = x_26861 & x_26862;
assign x_58149 = x_26863 & x_26864;
assign x_58150 = x_58148 & x_58149;
assign x_58151 = x_58147 & x_58150;
assign x_58152 = x_58144 & x_58151;
assign x_58153 = x_58137 & x_58152;
assign x_58154 = x_26866 & x_26867;
assign x_58155 = x_26865 & x_58154;
assign x_58156 = x_26868 & x_26869;
assign x_58157 = x_26870 & x_26871;
assign x_58158 = x_58156 & x_58157;
assign x_58159 = x_58155 & x_58158;
assign x_58160 = x_26872 & x_26873;
assign x_58161 = x_26874 & x_26875;
assign x_58162 = x_58160 & x_58161;
assign x_58163 = x_26876 & x_26877;
assign x_58164 = x_26878 & x_26879;
assign x_58165 = x_58163 & x_58164;
assign x_58166 = x_58162 & x_58165;
assign x_58167 = x_58159 & x_58166;
assign x_58168 = x_26880 & x_26881;
assign x_58169 = x_26882 & x_26883;
assign x_58170 = x_58168 & x_58169;
assign x_58171 = x_26884 & x_26885;
assign x_58172 = x_26886 & x_26887;
assign x_58173 = x_58171 & x_58172;
assign x_58174 = x_58170 & x_58173;
assign x_58175 = x_26888 & x_26889;
assign x_58176 = x_26890 & x_26891;
assign x_58177 = x_58175 & x_58176;
assign x_58178 = x_26892 & x_26893;
assign x_58179 = x_26894 & x_26895;
assign x_58180 = x_58178 & x_58179;
assign x_58181 = x_58177 & x_58180;
assign x_58182 = x_58174 & x_58181;
assign x_58183 = x_58167 & x_58182;
assign x_58184 = x_58153 & x_58183;
assign x_58185 = x_58123 & x_58184;
assign x_58186 = x_58063 & x_58185;
assign x_58187 = x_57942 & x_58186;
assign x_58188 = x_26897 & x_26898;
assign x_58189 = x_26896 & x_58188;
assign x_58190 = x_26899 & x_26900;
assign x_58191 = x_26901 & x_26902;
assign x_58192 = x_58190 & x_58191;
assign x_58193 = x_58189 & x_58192;
assign x_58194 = x_26903 & x_26904;
assign x_58195 = x_26905 & x_26906;
assign x_58196 = x_58194 & x_58195;
assign x_58197 = x_26907 & x_26908;
assign x_58198 = x_26909 & x_26910;
assign x_58199 = x_58197 & x_58198;
assign x_58200 = x_58196 & x_58199;
assign x_58201 = x_58193 & x_58200;
assign x_58202 = x_26912 & x_26913;
assign x_58203 = x_26911 & x_58202;
assign x_58204 = x_26914 & x_26915;
assign x_58205 = x_26916 & x_26917;
assign x_58206 = x_58204 & x_58205;
assign x_58207 = x_58203 & x_58206;
assign x_58208 = x_26918 & x_26919;
assign x_58209 = x_26920 & x_26921;
assign x_58210 = x_58208 & x_58209;
assign x_58211 = x_26922 & x_26923;
assign x_58212 = x_26924 & x_26925;
assign x_58213 = x_58211 & x_58212;
assign x_58214 = x_58210 & x_58213;
assign x_58215 = x_58207 & x_58214;
assign x_58216 = x_58201 & x_58215;
assign x_58217 = x_26927 & x_26928;
assign x_58218 = x_26926 & x_58217;
assign x_58219 = x_26929 & x_26930;
assign x_58220 = x_26931 & x_26932;
assign x_58221 = x_58219 & x_58220;
assign x_58222 = x_58218 & x_58221;
assign x_58223 = x_26933 & x_26934;
assign x_58224 = x_26935 & x_26936;
assign x_58225 = x_58223 & x_58224;
assign x_58226 = x_26937 & x_26938;
assign x_58227 = x_26939 & x_26940;
assign x_58228 = x_58226 & x_58227;
assign x_58229 = x_58225 & x_58228;
assign x_58230 = x_58222 & x_58229;
assign x_58231 = x_26941 & x_26942;
assign x_58232 = x_26943 & x_26944;
assign x_58233 = x_58231 & x_58232;
assign x_58234 = x_26945 & x_26946;
assign x_58235 = x_26947 & x_26948;
assign x_58236 = x_58234 & x_58235;
assign x_58237 = x_58233 & x_58236;
assign x_58238 = x_26949 & x_26950;
assign x_58239 = x_26951 & x_26952;
assign x_58240 = x_58238 & x_58239;
assign x_58241 = x_26953 & x_26954;
assign x_58242 = x_26955 & x_26956;
assign x_58243 = x_58241 & x_58242;
assign x_58244 = x_58240 & x_58243;
assign x_58245 = x_58237 & x_58244;
assign x_58246 = x_58230 & x_58245;
assign x_58247 = x_58216 & x_58246;
assign x_58248 = x_26958 & x_26959;
assign x_58249 = x_26957 & x_58248;
assign x_58250 = x_26960 & x_26961;
assign x_58251 = x_26962 & x_26963;
assign x_58252 = x_58250 & x_58251;
assign x_58253 = x_58249 & x_58252;
assign x_58254 = x_26964 & x_26965;
assign x_58255 = x_26966 & x_26967;
assign x_58256 = x_58254 & x_58255;
assign x_58257 = x_26968 & x_26969;
assign x_58258 = x_26970 & x_26971;
assign x_58259 = x_58257 & x_58258;
assign x_58260 = x_58256 & x_58259;
assign x_58261 = x_58253 & x_58260;
assign x_58262 = x_26973 & x_26974;
assign x_58263 = x_26972 & x_58262;
assign x_58264 = x_26975 & x_26976;
assign x_58265 = x_26977 & x_26978;
assign x_58266 = x_58264 & x_58265;
assign x_58267 = x_58263 & x_58266;
assign x_58268 = x_26979 & x_26980;
assign x_58269 = x_26981 & x_26982;
assign x_58270 = x_58268 & x_58269;
assign x_58271 = x_26983 & x_26984;
assign x_58272 = x_26985 & x_26986;
assign x_58273 = x_58271 & x_58272;
assign x_58274 = x_58270 & x_58273;
assign x_58275 = x_58267 & x_58274;
assign x_58276 = x_58261 & x_58275;
assign x_58277 = x_26988 & x_26989;
assign x_58278 = x_26987 & x_58277;
assign x_58279 = x_26990 & x_26991;
assign x_58280 = x_26992 & x_26993;
assign x_58281 = x_58279 & x_58280;
assign x_58282 = x_58278 & x_58281;
assign x_58283 = x_26994 & x_26995;
assign x_58284 = x_26996 & x_26997;
assign x_58285 = x_58283 & x_58284;
assign x_58286 = x_26998 & x_26999;
assign x_58287 = x_27000 & x_27001;
assign x_58288 = x_58286 & x_58287;
assign x_58289 = x_58285 & x_58288;
assign x_58290 = x_58282 & x_58289;
assign x_58291 = x_27002 & x_27003;
assign x_58292 = x_27004 & x_27005;
assign x_58293 = x_58291 & x_58292;
assign x_58294 = x_27006 & x_27007;
assign x_58295 = x_27008 & x_27009;
assign x_58296 = x_58294 & x_58295;
assign x_58297 = x_58293 & x_58296;
assign x_58298 = x_27010 & x_27011;
assign x_58299 = x_27012 & x_27013;
assign x_58300 = x_58298 & x_58299;
assign x_58301 = x_27014 & x_27015;
assign x_58302 = x_27016 & x_27017;
assign x_58303 = x_58301 & x_58302;
assign x_58304 = x_58300 & x_58303;
assign x_58305 = x_58297 & x_58304;
assign x_58306 = x_58290 & x_58305;
assign x_58307 = x_58276 & x_58306;
assign x_58308 = x_58247 & x_58307;
assign x_58309 = x_27019 & x_27020;
assign x_58310 = x_27018 & x_58309;
assign x_58311 = x_27021 & x_27022;
assign x_58312 = x_27023 & x_27024;
assign x_58313 = x_58311 & x_58312;
assign x_58314 = x_58310 & x_58313;
assign x_58315 = x_27025 & x_27026;
assign x_58316 = x_27027 & x_27028;
assign x_58317 = x_58315 & x_58316;
assign x_58318 = x_27029 & x_27030;
assign x_58319 = x_27031 & x_27032;
assign x_58320 = x_58318 & x_58319;
assign x_58321 = x_58317 & x_58320;
assign x_58322 = x_58314 & x_58321;
assign x_58323 = x_27034 & x_27035;
assign x_58324 = x_27033 & x_58323;
assign x_58325 = x_27036 & x_27037;
assign x_58326 = x_27038 & x_27039;
assign x_58327 = x_58325 & x_58326;
assign x_58328 = x_58324 & x_58327;
assign x_58329 = x_27040 & x_27041;
assign x_58330 = x_27042 & x_27043;
assign x_58331 = x_58329 & x_58330;
assign x_58332 = x_27044 & x_27045;
assign x_58333 = x_27046 & x_27047;
assign x_58334 = x_58332 & x_58333;
assign x_58335 = x_58331 & x_58334;
assign x_58336 = x_58328 & x_58335;
assign x_58337 = x_58322 & x_58336;
assign x_58338 = x_27049 & x_27050;
assign x_58339 = x_27048 & x_58338;
assign x_58340 = x_27051 & x_27052;
assign x_58341 = x_27053 & x_27054;
assign x_58342 = x_58340 & x_58341;
assign x_58343 = x_58339 & x_58342;
assign x_58344 = x_27055 & x_27056;
assign x_58345 = x_27057 & x_27058;
assign x_58346 = x_58344 & x_58345;
assign x_58347 = x_27059 & x_27060;
assign x_58348 = x_27061 & x_27062;
assign x_58349 = x_58347 & x_58348;
assign x_58350 = x_58346 & x_58349;
assign x_58351 = x_58343 & x_58350;
assign x_58352 = x_27063 & x_27064;
assign x_58353 = x_27065 & x_27066;
assign x_58354 = x_58352 & x_58353;
assign x_58355 = x_27067 & x_27068;
assign x_58356 = x_27069 & x_27070;
assign x_58357 = x_58355 & x_58356;
assign x_58358 = x_58354 & x_58357;
assign x_58359 = x_27071 & x_27072;
assign x_58360 = x_27073 & x_27074;
assign x_58361 = x_58359 & x_58360;
assign x_58362 = x_27075 & x_27076;
assign x_58363 = x_27077 & x_27078;
assign x_58364 = x_58362 & x_58363;
assign x_58365 = x_58361 & x_58364;
assign x_58366 = x_58358 & x_58365;
assign x_58367 = x_58351 & x_58366;
assign x_58368 = x_58337 & x_58367;
assign x_58369 = x_27080 & x_27081;
assign x_58370 = x_27079 & x_58369;
assign x_58371 = x_27082 & x_27083;
assign x_58372 = x_27084 & x_27085;
assign x_58373 = x_58371 & x_58372;
assign x_58374 = x_58370 & x_58373;
assign x_58375 = x_27086 & x_27087;
assign x_58376 = x_27088 & x_27089;
assign x_58377 = x_58375 & x_58376;
assign x_58378 = x_27090 & x_27091;
assign x_58379 = x_27092 & x_27093;
assign x_58380 = x_58378 & x_58379;
assign x_58381 = x_58377 & x_58380;
assign x_58382 = x_58374 & x_58381;
assign x_58383 = x_27095 & x_27096;
assign x_58384 = x_27094 & x_58383;
assign x_58385 = x_27097 & x_27098;
assign x_58386 = x_27099 & x_27100;
assign x_58387 = x_58385 & x_58386;
assign x_58388 = x_58384 & x_58387;
assign x_58389 = x_27101 & x_27102;
assign x_58390 = x_27103 & x_27104;
assign x_58391 = x_58389 & x_58390;
assign x_58392 = x_27105 & x_27106;
assign x_58393 = x_27107 & x_27108;
assign x_58394 = x_58392 & x_58393;
assign x_58395 = x_58391 & x_58394;
assign x_58396 = x_58388 & x_58395;
assign x_58397 = x_58382 & x_58396;
assign x_58398 = x_27110 & x_27111;
assign x_58399 = x_27109 & x_58398;
assign x_58400 = x_27112 & x_27113;
assign x_58401 = x_27114 & x_27115;
assign x_58402 = x_58400 & x_58401;
assign x_58403 = x_58399 & x_58402;
assign x_58404 = x_27116 & x_27117;
assign x_58405 = x_27118 & x_27119;
assign x_58406 = x_58404 & x_58405;
assign x_58407 = x_27120 & x_27121;
assign x_58408 = x_27122 & x_27123;
assign x_58409 = x_58407 & x_58408;
assign x_58410 = x_58406 & x_58409;
assign x_58411 = x_58403 & x_58410;
assign x_58412 = x_27124 & x_27125;
assign x_58413 = x_27126 & x_27127;
assign x_58414 = x_58412 & x_58413;
assign x_58415 = x_27128 & x_27129;
assign x_58416 = x_27130 & x_27131;
assign x_58417 = x_58415 & x_58416;
assign x_58418 = x_58414 & x_58417;
assign x_58419 = x_27132 & x_27133;
assign x_58420 = x_27134 & x_27135;
assign x_58421 = x_58419 & x_58420;
assign x_58422 = x_27136 & x_27137;
assign x_58423 = x_27138 & x_27139;
assign x_58424 = x_58422 & x_58423;
assign x_58425 = x_58421 & x_58424;
assign x_58426 = x_58418 & x_58425;
assign x_58427 = x_58411 & x_58426;
assign x_58428 = x_58397 & x_58427;
assign x_58429 = x_58368 & x_58428;
assign x_58430 = x_58308 & x_58429;
assign x_58431 = x_27141 & x_27142;
assign x_58432 = x_27140 & x_58431;
assign x_58433 = x_27143 & x_27144;
assign x_58434 = x_27145 & x_27146;
assign x_58435 = x_58433 & x_58434;
assign x_58436 = x_58432 & x_58435;
assign x_58437 = x_27147 & x_27148;
assign x_58438 = x_27149 & x_27150;
assign x_58439 = x_58437 & x_58438;
assign x_58440 = x_27151 & x_27152;
assign x_58441 = x_27153 & x_27154;
assign x_58442 = x_58440 & x_58441;
assign x_58443 = x_58439 & x_58442;
assign x_58444 = x_58436 & x_58443;
assign x_58445 = x_27156 & x_27157;
assign x_58446 = x_27155 & x_58445;
assign x_58447 = x_27158 & x_27159;
assign x_58448 = x_27160 & x_27161;
assign x_58449 = x_58447 & x_58448;
assign x_58450 = x_58446 & x_58449;
assign x_58451 = x_27162 & x_27163;
assign x_58452 = x_27164 & x_27165;
assign x_58453 = x_58451 & x_58452;
assign x_58454 = x_27166 & x_27167;
assign x_58455 = x_27168 & x_27169;
assign x_58456 = x_58454 & x_58455;
assign x_58457 = x_58453 & x_58456;
assign x_58458 = x_58450 & x_58457;
assign x_58459 = x_58444 & x_58458;
assign x_58460 = x_27171 & x_27172;
assign x_58461 = x_27170 & x_58460;
assign x_58462 = x_27173 & x_27174;
assign x_58463 = x_27175 & x_27176;
assign x_58464 = x_58462 & x_58463;
assign x_58465 = x_58461 & x_58464;
assign x_58466 = x_27177 & x_27178;
assign x_58467 = x_27179 & x_27180;
assign x_58468 = x_58466 & x_58467;
assign x_58469 = x_27181 & x_27182;
assign x_58470 = x_27183 & x_27184;
assign x_58471 = x_58469 & x_58470;
assign x_58472 = x_58468 & x_58471;
assign x_58473 = x_58465 & x_58472;
assign x_58474 = x_27185 & x_27186;
assign x_58475 = x_27187 & x_27188;
assign x_58476 = x_58474 & x_58475;
assign x_58477 = x_27189 & x_27190;
assign x_58478 = x_27191 & x_27192;
assign x_58479 = x_58477 & x_58478;
assign x_58480 = x_58476 & x_58479;
assign x_58481 = x_27193 & x_27194;
assign x_58482 = x_27195 & x_27196;
assign x_58483 = x_58481 & x_58482;
assign x_58484 = x_27197 & x_27198;
assign x_58485 = x_27199 & x_27200;
assign x_58486 = x_58484 & x_58485;
assign x_58487 = x_58483 & x_58486;
assign x_58488 = x_58480 & x_58487;
assign x_58489 = x_58473 & x_58488;
assign x_58490 = x_58459 & x_58489;
assign x_58491 = x_27202 & x_27203;
assign x_58492 = x_27201 & x_58491;
assign x_58493 = x_27204 & x_27205;
assign x_58494 = x_27206 & x_27207;
assign x_58495 = x_58493 & x_58494;
assign x_58496 = x_58492 & x_58495;
assign x_58497 = x_27208 & x_27209;
assign x_58498 = x_27210 & x_27211;
assign x_58499 = x_58497 & x_58498;
assign x_58500 = x_27212 & x_27213;
assign x_58501 = x_27214 & x_27215;
assign x_58502 = x_58500 & x_58501;
assign x_58503 = x_58499 & x_58502;
assign x_58504 = x_58496 & x_58503;
assign x_58505 = x_27217 & x_27218;
assign x_58506 = x_27216 & x_58505;
assign x_58507 = x_27219 & x_27220;
assign x_58508 = x_27221 & x_27222;
assign x_58509 = x_58507 & x_58508;
assign x_58510 = x_58506 & x_58509;
assign x_58511 = x_27223 & x_27224;
assign x_58512 = x_27225 & x_27226;
assign x_58513 = x_58511 & x_58512;
assign x_58514 = x_27227 & x_27228;
assign x_58515 = x_27229 & x_27230;
assign x_58516 = x_58514 & x_58515;
assign x_58517 = x_58513 & x_58516;
assign x_58518 = x_58510 & x_58517;
assign x_58519 = x_58504 & x_58518;
assign x_58520 = x_27232 & x_27233;
assign x_58521 = x_27231 & x_58520;
assign x_58522 = x_27234 & x_27235;
assign x_58523 = x_27236 & x_27237;
assign x_58524 = x_58522 & x_58523;
assign x_58525 = x_58521 & x_58524;
assign x_58526 = x_27238 & x_27239;
assign x_58527 = x_27240 & x_27241;
assign x_58528 = x_58526 & x_58527;
assign x_58529 = x_27242 & x_27243;
assign x_58530 = x_27244 & x_27245;
assign x_58531 = x_58529 & x_58530;
assign x_58532 = x_58528 & x_58531;
assign x_58533 = x_58525 & x_58532;
assign x_58534 = x_27246 & x_27247;
assign x_58535 = x_27248 & x_27249;
assign x_58536 = x_58534 & x_58535;
assign x_58537 = x_27250 & x_27251;
assign x_58538 = x_27252 & x_27253;
assign x_58539 = x_58537 & x_58538;
assign x_58540 = x_58536 & x_58539;
assign x_58541 = x_27254 & x_27255;
assign x_58542 = x_27256 & x_27257;
assign x_58543 = x_58541 & x_58542;
assign x_58544 = x_27258 & x_27259;
assign x_58545 = x_27260 & x_27261;
assign x_58546 = x_58544 & x_58545;
assign x_58547 = x_58543 & x_58546;
assign x_58548 = x_58540 & x_58547;
assign x_58549 = x_58533 & x_58548;
assign x_58550 = x_58519 & x_58549;
assign x_58551 = x_58490 & x_58550;
assign x_58552 = x_27263 & x_27264;
assign x_58553 = x_27262 & x_58552;
assign x_58554 = x_27265 & x_27266;
assign x_58555 = x_27267 & x_27268;
assign x_58556 = x_58554 & x_58555;
assign x_58557 = x_58553 & x_58556;
assign x_58558 = x_27269 & x_27270;
assign x_58559 = x_27271 & x_27272;
assign x_58560 = x_58558 & x_58559;
assign x_58561 = x_27273 & x_27274;
assign x_58562 = x_27275 & x_27276;
assign x_58563 = x_58561 & x_58562;
assign x_58564 = x_58560 & x_58563;
assign x_58565 = x_58557 & x_58564;
assign x_58566 = x_27278 & x_27279;
assign x_58567 = x_27277 & x_58566;
assign x_58568 = x_27280 & x_27281;
assign x_58569 = x_27282 & x_27283;
assign x_58570 = x_58568 & x_58569;
assign x_58571 = x_58567 & x_58570;
assign x_58572 = x_27284 & x_27285;
assign x_58573 = x_27286 & x_27287;
assign x_58574 = x_58572 & x_58573;
assign x_58575 = x_27288 & x_27289;
assign x_58576 = x_27290 & x_27291;
assign x_58577 = x_58575 & x_58576;
assign x_58578 = x_58574 & x_58577;
assign x_58579 = x_58571 & x_58578;
assign x_58580 = x_58565 & x_58579;
assign x_58581 = x_27293 & x_27294;
assign x_58582 = x_27292 & x_58581;
assign x_58583 = x_27295 & x_27296;
assign x_58584 = x_27297 & x_27298;
assign x_58585 = x_58583 & x_58584;
assign x_58586 = x_58582 & x_58585;
assign x_58587 = x_27299 & x_27300;
assign x_58588 = x_27301 & x_27302;
assign x_58589 = x_58587 & x_58588;
assign x_58590 = x_27303 & x_27304;
assign x_58591 = x_27305 & x_27306;
assign x_58592 = x_58590 & x_58591;
assign x_58593 = x_58589 & x_58592;
assign x_58594 = x_58586 & x_58593;
assign x_58595 = x_27307 & x_27308;
assign x_58596 = x_27309 & x_27310;
assign x_58597 = x_58595 & x_58596;
assign x_58598 = x_27311 & x_27312;
assign x_58599 = x_27313 & x_27314;
assign x_58600 = x_58598 & x_58599;
assign x_58601 = x_58597 & x_58600;
assign x_58602 = x_27315 & x_27316;
assign x_58603 = x_27317 & x_27318;
assign x_58604 = x_58602 & x_58603;
assign x_58605 = x_27319 & x_27320;
assign x_58606 = x_27321 & x_27322;
assign x_58607 = x_58605 & x_58606;
assign x_58608 = x_58604 & x_58607;
assign x_58609 = x_58601 & x_58608;
assign x_58610 = x_58594 & x_58609;
assign x_58611 = x_58580 & x_58610;
assign x_58612 = x_27324 & x_27325;
assign x_58613 = x_27323 & x_58612;
assign x_58614 = x_27326 & x_27327;
assign x_58615 = x_27328 & x_27329;
assign x_58616 = x_58614 & x_58615;
assign x_58617 = x_58613 & x_58616;
assign x_58618 = x_27330 & x_27331;
assign x_58619 = x_27332 & x_27333;
assign x_58620 = x_58618 & x_58619;
assign x_58621 = x_27334 & x_27335;
assign x_58622 = x_27336 & x_27337;
assign x_58623 = x_58621 & x_58622;
assign x_58624 = x_58620 & x_58623;
assign x_58625 = x_58617 & x_58624;
assign x_58626 = x_27338 & x_27339;
assign x_58627 = x_27340 & x_27341;
assign x_58628 = x_58626 & x_58627;
assign x_58629 = x_27342 & x_27343;
assign x_58630 = x_27344 & x_27345;
assign x_58631 = x_58629 & x_58630;
assign x_58632 = x_58628 & x_58631;
assign x_58633 = x_27346 & x_27347;
assign x_58634 = x_27348 & x_27349;
assign x_58635 = x_58633 & x_58634;
assign x_58636 = x_27350 & x_27351;
assign x_58637 = x_27352 & x_27353;
assign x_58638 = x_58636 & x_58637;
assign x_58639 = x_58635 & x_58638;
assign x_58640 = x_58632 & x_58639;
assign x_58641 = x_58625 & x_58640;
assign x_58642 = x_27355 & x_27356;
assign x_58643 = x_27354 & x_58642;
assign x_58644 = x_27357 & x_27358;
assign x_58645 = x_27359 & x_27360;
assign x_58646 = x_58644 & x_58645;
assign x_58647 = x_58643 & x_58646;
assign x_58648 = x_27361 & x_27362;
assign x_58649 = x_27363 & x_27364;
assign x_58650 = x_58648 & x_58649;
assign x_58651 = x_27365 & x_27366;
assign x_58652 = x_27367 & x_27368;
assign x_58653 = x_58651 & x_58652;
assign x_58654 = x_58650 & x_58653;
assign x_58655 = x_58647 & x_58654;
assign x_58656 = x_27369 & x_27370;
assign x_58657 = x_27371 & x_27372;
assign x_58658 = x_58656 & x_58657;
assign x_58659 = x_27373 & x_27374;
assign x_58660 = x_27375 & x_27376;
assign x_58661 = x_58659 & x_58660;
assign x_58662 = x_58658 & x_58661;
assign x_58663 = x_27377 & x_27378;
assign x_58664 = x_27379 & x_27380;
assign x_58665 = x_58663 & x_58664;
assign x_58666 = x_27381 & x_27382;
assign x_58667 = x_27383 & x_27384;
assign x_58668 = x_58666 & x_58667;
assign x_58669 = x_58665 & x_58668;
assign x_58670 = x_58662 & x_58669;
assign x_58671 = x_58655 & x_58670;
assign x_58672 = x_58641 & x_58671;
assign x_58673 = x_58611 & x_58672;
assign x_58674 = x_58551 & x_58673;
assign x_58675 = x_58430 & x_58674;
assign x_58676 = x_58187 & x_58675;
assign x_58677 = x_57699 & x_58676;
assign x_58678 = x_56722 & x_58677;
assign x_58679 = x_27386 & x_27387;
assign x_58680 = x_27385 & x_58679;
assign x_58681 = x_27388 & x_27389;
assign x_58682 = x_27390 & x_27391;
assign x_58683 = x_58681 & x_58682;
assign x_58684 = x_58680 & x_58683;
assign x_58685 = x_27392 & x_27393;
assign x_58686 = x_27394 & x_27395;
assign x_58687 = x_58685 & x_58686;
assign x_58688 = x_27396 & x_27397;
assign x_58689 = x_27398 & x_27399;
assign x_58690 = x_58688 & x_58689;
assign x_58691 = x_58687 & x_58690;
assign x_58692 = x_58684 & x_58691;
assign x_58693 = x_27401 & x_27402;
assign x_58694 = x_27400 & x_58693;
assign x_58695 = x_27403 & x_27404;
assign x_58696 = x_27405 & x_27406;
assign x_58697 = x_58695 & x_58696;
assign x_58698 = x_58694 & x_58697;
assign x_58699 = x_27407 & x_27408;
assign x_58700 = x_27409 & x_27410;
assign x_58701 = x_58699 & x_58700;
assign x_58702 = x_27411 & x_27412;
assign x_58703 = x_27413 & x_27414;
assign x_58704 = x_58702 & x_58703;
assign x_58705 = x_58701 & x_58704;
assign x_58706 = x_58698 & x_58705;
assign x_58707 = x_58692 & x_58706;
assign x_58708 = x_27416 & x_27417;
assign x_58709 = x_27415 & x_58708;
assign x_58710 = x_27418 & x_27419;
assign x_58711 = x_27420 & x_27421;
assign x_58712 = x_58710 & x_58711;
assign x_58713 = x_58709 & x_58712;
assign x_58714 = x_27422 & x_27423;
assign x_58715 = x_27424 & x_27425;
assign x_58716 = x_58714 & x_58715;
assign x_58717 = x_27426 & x_27427;
assign x_58718 = x_27428 & x_27429;
assign x_58719 = x_58717 & x_58718;
assign x_58720 = x_58716 & x_58719;
assign x_58721 = x_58713 & x_58720;
assign x_58722 = x_27430 & x_27431;
assign x_58723 = x_27432 & x_27433;
assign x_58724 = x_58722 & x_58723;
assign x_58725 = x_27434 & x_27435;
assign x_58726 = x_27436 & x_27437;
assign x_58727 = x_58725 & x_58726;
assign x_58728 = x_58724 & x_58727;
assign x_58729 = x_27438 & x_27439;
assign x_58730 = x_27440 & x_27441;
assign x_58731 = x_58729 & x_58730;
assign x_58732 = x_27442 & x_27443;
assign x_58733 = x_27444 & x_27445;
assign x_58734 = x_58732 & x_58733;
assign x_58735 = x_58731 & x_58734;
assign x_58736 = x_58728 & x_58735;
assign x_58737 = x_58721 & x_58736;
assign x_58738 = x_58707 & x_58737;
assign x_58739 = x_27447 & x_27448;
assign x_58740 = x_27446 & x_58739;
assign x_58741 = x_27449 & x_27450;
assign x_58742 = x_27451 & x_27452;
assign x_58743 = x_58741 & x_58742;
assign x_58744 = x_58740 & x_58743;
assign x_58745 = x_27453 & x_27454;
assign x_58746 = x_27455 & x_27456;
assign x_58747 = x_58745 & x_58746;
assign x_58748 = x_27457 & x_27458;
assign x_58749 = x_27459 & x_27460;
assign x_58750 = x_58748 & x_58749;
assign x_58751 = x_58747 & x_58750;
assign x_58752 = x_58744 & x_58751;
assign x_58753 = x_27462 & x_27463;
assign x_58754 = x_27461 & x_58753;
assign x_58755 = x_27464 & x_27465;
assign x_58756 = x_27466 & x_27467;
assign x_58757 = x_58755 & x_58756;
assign x_58758 = x_58754 & x_58757;
assign x_58759 = x_27468 & x_27469;
assign x_58760 = x_27470 & x_27471;
assign x_58761 = x_58759 & x_58760;
assign x_58762 = x_27472 & x_27473;
assign x_58763 = x_27474 & x_27475;
assign x_58764 = x_58762 & x_58763;
assign x_58765 = x_58761 & x_58764;
assign x_58766 = x_58758 & x_58765;
assign x_58767 = x_58752 & x_58766;
assign x_58768 = x_27477 & x_27478;
assign x_58769 = x_27476 & x_58768;
assign x_58770 = x_27479 & x_27480;
assign x_58771 = x_27481 & x_27482;
assign x_58772 = x_58770 & x_58771;
assign x_58773 = x_58769 & x_58772;
assign x_58774 = x_27483 & x_27484;
assign x_58775 = x_27485 & x_27486;
assign x_58776 = x_58774 & x_58775;
assign x_58777 = x_27487 & x_27488;
assign x_58778 = x_27489 & x_27490;
assign x_58779 = x_58777 & x_58778;
assign x_58780 = x_58776 & x_58779;
assign x_58781 = x_58773 & x_58780;
assign x_58782 = x_27491 & x_27492;
assign x_58783 = x_27493 & x_27494;
assign x_58784 = x_58782 & x_58783;
assign x_58785 = x_27495 & x_27496;
assign x_58786 = x_27497 & x_27498;
assign x_58787 = x_58785 & x_58786;
assign x_58788 = x_58784 & x_58787;
assign x_58789 = x_27499 & x_27500;
assign x_58790 = x_27501 & x_27502;
assign x_58791 = x_58789 & x_58790;
assign x_58792 = x_27503 & x_27504;
assign x_58793 = x_27505 & x_27506;
assign x_58794 = x_58792 & x_58793;
assign x_58795 = x_58791 & x_58794;
assign x_58796 = x_58788 & x_58795;
assign x_58797 = x_58781 & x_58796;
assign x_58798 = x_58767 & x_58797;
assign x_58799 = x_58738 & x_58798;
assign x_58800 = x_27508 & x_27509;
assign x_58801 = x_27507 & x_58800;
assign x_58802 = x_27510 & x_27511;
assign x_58803 = x_27512 & x_27513;
assign x_58804 = x_58802 & x_58803;
assign x_58805 = x_58801 & x_58804;
assign x_58806 = x_27514 & x_27515;
assign x_58807 = x_27516 & x_27517;
assign x_58808 = x_58806 & x_58807;
assign x_58809 = x_27518 & x_27519;
assign x_58810 = x_27520 & x_27521;
assign x_58811 = x_58809 & x_58810;
assign x_58812 = x_58808 & x_58811;
assign x_58813 = x_58805 & x_58812;
assign x_58814 = x_27523 & x_27524;
assign x_58815 = x_27522 & x_58814;
assign x_58816 = x_27525 & x_27526;
assign x_58817 = x_27527 & x_27528;
assign x_58818 = x_58816 & x_58817;
assign x_58819 = x_58815 & x_58818;
assign x_58820 = x_27529 & x_27530;
assign x_58821 = x_27531 & x_27532;
assign x_58822 = x_58820 & x_58821;
assign x_58823 = x_27533 & x_27534;
assign x_58824 = x_27535 & x_27536;
assign x_58825 = x_58823 & x_58824;
assign x_58826 = x_58822 & x_58825;
assign x_58827 = x_58819 & x_58826;
assign x_58828 = x_58813 & x_58827;
assign x_58829 = x_27538 & x_27539;
assign x_58830 = x_27537 & x_58829;
assign x_58831 = x_27540 & x_27541;
assign x_58832 = x_27542 & x_27543;
assign x_58833 = x_58831 & x_58832;
assign x_58834 = x_58830 & x_58833;
assign x_58835 = x_27544 & x_27545;
assign x_58836 = x_27546 & x_27547;
assign x_58837 = x_58835 & x_58836;
assign x_58838 = x_27548 & x_27549;
assign x_58839 = x_27550 & x_27551;
assign x_58840 = x_58838 & x_58839;
assign x_58841 = x_58837 & x_58840;
assign x_58842 = x_58834 & x_58841;
assign x_58843 = x_27552 & x_27553;
assign x_58844 = x_27554 & x_27555;
assign x_58845 = x_58843 & x_58844;
assign x_58846 = x_27556 & x_27557;
assign x_58847 = x_27558 & x_27559;
assign x_58848 = x_58846 & x_58847;
assign x_58849 = x_58845 & x_58848;
assign x_58850 = x_27560 & x_27561;
assign x_58851 = x_27562 & x_27563;
assign x_58852 = x_58850 & x_58851;
assign x_58853 = x_27564 & x_27565;
assign x_58854 = x_27566 & x_27567;
assign x_58855 = x_58853 & x_58854;
assign x_58856 = x_58852 & x_58855;
assign x_58857 = x_58849 & x_58856;
assign x_58858 = x_58842 & x_58857;
assign x_58859 = x_58828 & x_58858;
assign x_58860 = x_27569 & x_27570;
assign x_58861 = x_27568 & x_58860;
assign x_58862 = x_27571 & x_27572;
assign x_58863 = x_27573 & x_27574;
assign x_58864 = x_58862 & x_58863;
assign x_58865 = x_58861 & x_58864;
assign x_58866 = x_27575 & x_27576;
assign x_58867 = x_27577 & x_27578;
assign x_58868 = x_58866 & x_58867;
assign x_58869 = x_27579 & x_27580;
assign x_58870 = x_27581 & x_27582;
assign x_58871 = x_58869 & x_58870;
assign x_58872 = x_58868 & x_58871;
assign x_58873 = x_58865 & x_58872;
assign x_58874 = x_27584 & x_27585;
assign x_58875 = x_27583 & x_58874;
assign x_58876 = x_27586 & x_27587;
assign x_58877 = x_27588 & x_27589;
assign x_58878 = x_58876 & x_58877;
assign x_58879 = x_58875 & x_58878;
assign x_58880 = x_27590 & x_27591;
assign x_58881 = x_27592 & x_27593;
assign x_58882 = x_58880 & x_58881;
assign x_58883 = x_27594 & x_27595;
assign x_58884 = x_27596 & x_27597;
assign x_58885 = x_58883 & x_58884;
assign x_58886 = x_58882 & x_58885;
assign x_58887 = x_58879 & x_58886;
assign x_58888 = x_58873 & x_58887;
assign x_58889 = x_27599 & x_27600;
assign x_58890 = x_27598 & x_58889;
assign x_58891 = x_27601 & x_27602;
assign x_58892 = x_27603 & x_27604;
assign x_58893 = x_58891 & x_58892;
assign x_58894 = x_58890 & x_58893;
assign x_58895 = x_27605 & x_27606;
assign x_58896 = x_27607 & x_27608;
assign x_58897 = x_58895 & x_58896;
assign x_58898 = x_27609 & x_27610;
assign x_58899 = x_27611 & x_27612;
assign x_58900 = x_58898 & x_58899;
assign x_58901 = x_58897 & x_58900;
assign x_58902 = x_58894 & x_58901;
assign x_58903 = x_27613 & x_27614;
assign x_58904 = x_27615 & x_27616;
assign x_58905 = x_58903 & x_58904;
assign x_58906 = x_27617 & x_27618;
assign x_58907 = x_27619 & x_27620;
assign x_58908 = x_58906 & x_58907;
assign x_58909 = x_58905 & x_58908;
assign x_58910 = x_27621 & x_27622;
assign x_58911 = x_27623 & x_27624;
assign x_58912 = x_58910 & x_58911;
assign x_58913 = x_27625 & x_27626;
assign x_58914 = x_27627 & x_27628;
assign x_58915 = x_58913 & x_58914;
assign x_58916 = x_58912 & x_58915;
assign x_58917 = x_58909 & x_58916;
assign x_58918 = x_58902 & x_58917;
assign x_58919 = x_58888 & x_58918;
assign x_58920 = x_58859 & x_58919;
assign x_58921 = x_58799 & x_58920;
assign x_58922 = x_27630 & x_27631;
assign x_58923 = x_27629 & x_58922;
assign x_58924 = x_27632 & x_27633;
assign x_58925 = x_27634 & x_27635;
assign x_58926 = x_58924 & x_58925;
assign x_58927 = x_58923 & x_58926;
assign x_58928 = x_27636 & x_27637;
assign x_58929 = x_27638 & x_27639;
assign x_58930 = x_58928 & x_58929;
assign x_58931 = x_27640 & x_27641;
assign x_58932 = x_27642 & x_27643;
assign x_58933 = x_58931 & x_58932;
assign x_58934 = x_58930 & x_58933;
assign x_58935 = x_58927 & x_58934;
assign x_58936 = x_27645 & x_27646;
assign x_58937 = x_27644 & x_58936;
assign x_58938 = x_27647 & x_27648;
assign x_58939 = x_27649 & x_27650;
assign x_58940 = x_58938 & x_58939;
assign x_58941 = x_58937 & x_58940;
assign x_58942 = x_27651 & x_27652;
assign x_58943 = x_27653 & x_27654;
assign x_58944 = x_58942 & x_58943;
assign x_58945 = x_27655 & x_27656;
assign x_58946 = x_27657 & x_27658;
assign x_58947 = x_58945 & x_58946;
assign x_58948 = x_58944 & x_58947;
assign x_58949 = x_58941 & x_58948;
assign x_58950 = x_58935 & x_58949;
assign x_58951 = x_27660 & x_27661;
assign x_58952 = x_27659 & x_58951;
assign x_58953 = x_27662 & x_27663;
assign x_58954 = x_27664 & x_27665;
assign x_58955 = x_58953 & x_58954;
assign x_58956 = x_58952 & x_58955;
assign x_58957 = x_27666 & x_27667;
assign x_58958 = x_27668 & x_27669;
assign x_58959 = x_58957 & x_58958;
assign x_58960 = x_27670 & x_27671;
assign x_58961 = x_27672 & x_27673;
assign x_58962 = x_58960 & x_58961;
assign x_58963 = x_58959 & x_58962;
assign x_58964 = x_58956 & x_58963;
assign x_58965 = x_27674 & x_27675;
assign x_58966 = x_27676 & x_27677;
assign x_58967 = x_58965 & x_58966;
assign x_58968 = x_27678 & x_27679;
assign x_58969 = x_27680 & x_27681;
assign x_58970 = x_58968 & x_58969;
assign x_58971 = x_58967 & x_58970;
assign x_58972 = x_27682 & x_27683;
assign x_58973 = x_27684 & x_27685;
assign x_58974 = x_58972 & x_58973;
assign x_58975 = x_27686 & x_27687;
assign x_58976 = x_27688 & x_27689;
assign x_58977 = x_58975 & x_58976;
assign x_58978 = x_58974 & x_58977;
assign x_58979 = x_58971 & x_58978;
assign x_58980 = x_58964 & x_58979;
assign x_58981 = x_58950 & x_58980;
assign x_58982 = x_27691 & x_27692;
assign x_58983 = x_27690 & x_58982;
assign x_58984 = x_27693 & x_27694;
assign x_58985 = x_27695 & x_27696;
assign x_58986 = x_58984 & x_58985;
assign x_58987 = x_58983 & x_58986;
assign x_58988 = x_27697 & x_27698;
assign x_58989 = x_27699 & x_27700;
assign x_58990 = x_58988 & x_58989;
assign x_58991 = x_27701 & x_27702;
assign x_58992 = x_27703 & x_27704;
assign x_58993 = x_58991 & x_58992;
assign x_58994 = x_58990 & x_58993;
assign x_58995 = x_58987 & x_58994;
assign x_58996 = x_27706 & x_27707;
assign x_58997 = x_27705 & x_58996;
assign x_58998 = x_27708 & x_27709;
assign x_58999 = x_27710 & x_27711;
assign x_59000 = x_58998 & x_58999;
assign x_59001 = x_58997 & x_59000;
assign x_59002 = x_27712 & x_27713;
assign x_59003 = x_27714 & x_27715;
assign x_59004 = x_59002 & x_59003;
assign x_59005 = x_27716 & x_27717;
assign x_59006 = x_27718 & x_27719;
assign x_59007 = x_59005 & x_59006;
assign x_59008 = x_59004 & x_59007;
assign x_59009 = x_59001 & x_59008;
assign x_59010 = x_58995 & x_59009;
assign x_59011 = x_27721 & x_27722;
assign x_59012 = x_27720 & x_59011;
assign x_59013 = x_27723 & x_27724;
assign x_59014 = x_27725 & x_27726;
assign x_59015 = x_59013 & x_59014;
assign x_59016 = x_59012 & x_59015;
assign x_59017 = x_27727 & x_27728;
assign x_59018 = x_27729 & x_27730;
assign x_59019 = x_59017 & x_59018;
assign x_59020 = x_27731 & x_27732;
assign x_59021 = x_27733 & x_27734;
assign x_59022 = x_59020 & x_59021;
assign x_59023 = x_59019 & x_59022;
assign x_59024 = x_59016 & x_59023;
assign x_59025 = x_27735 & x_27736;
assign x_59026 = x_27737 & x_27738;
assign x_59027 = x_59025 & x_59026;
assign x_59028 = x_27739 & x_27740;
assign x_59029 = x_27741 & x_27742;
assign x_59030 = x_59028 & x_59029;
assign x_59031 = x_59027 & x_59030;
assign x_59032 = x_27743 & x_27744;
assign x_59033 = x_27745 & x_27746;
assign x_59034 = x_59032 & x_59033;
assign x_59035 = x_27747 & x_27748;
assign x_59036 = x_27749 & x_27750;
assign x_59037 = x_59035 & x_59036;
assign x_59038 = x_59034 & x_59037;
assign x_59039 = x_59031 & x_59038;
assign x_59040 = x_59024 & x_59039;
assign x_59041 = x_59010 & x_59040;
assign x_59042 = x_58981 & x_59041;
assign x_59043 = x_27752 & x_27753;
assign x_59044 = x_27751 & x_59043;
assign x_59045 = x_27754 & x_27755;
assign x_59046 = x_27756 & x_27757;
assign x_59047 = x_59045 & x_59046;
assign x_59048 = x_59044 & x_59047;
assign x_59049 = x_27758 & x_27759;
assign x_59050 = x_27760 & x_27761;
assign x_59051 = x_59049 & x_59050;
assign x_59052 = x_27762 & x_27763;
assign x_59053 = x_27764 & x_27765;
assign x_59054 = x_59052 & x_59053;
assign x_59055 = x_59051 & x_59054;
assign x_59056 = x_59048 & x_59055;
assign x_59057 = x_27767 & x_27768;
assign x_59058 = x_27766 & x_59057;
assign x_59059 = x_27769 & x_27770;
assign x_59060 = x_27771 & x_27772;
assign x_59061 = x_59059 & x_59060;
assign x_59062 = x_59058 & x_59061;
assign x_59063 = x_27773 & x_27774;
assign x_59064 = x_27775 & x_27776;
assign x_59065 = x_59063 & x_59064;
assign x_59066 = x_27777 & x_27778;
assign x_59067 = x_27779 & x_27780;
assign x_59068 = x_59066 & x_59067;
assign x_59069 = x_59065 & x_59068;
assign x_59070 = x_59062 & x_59069;
assign x_59071 = x_59056 & x_59070;
assign x_59072 = x_27782 & x_27783;
assign x_59073 = x_27781 & x_59072;
assign x_59074 = x_27784 & x_27785;
assign x_59075 = x_27786 & x_27787;
assign x_59076 = x_59074 & x_59075;
assign x_59077 = x_59073 & x_59076;
assign x_59078 = x_27788 & x_27789;
assign x_59079 = x_27790 & x_27791;
assign x_59080 = x_59078 & x_59079;
assign x_59081 = x_27792 & x_27793;
assign x_59082 = x_27794 & x_27795;
assign x_59083 = x_59081 & x_59082;
assign x_59084 = x_59080 & x_59083;
assign x_59085 = x_59077 & x_59084;
assign x_59086 = x_27796 & x_27797;
assign x_59087 = x_27798 & x_27799;
assign x_59088 = x_59086 & x_59087;
assign x_59089 = x_27800 & x_27801;
assign x_59090 = x_27802 & x_27803;
assign x_59091 = x_59089 & x_59090;
assign x_59092 = x_59088 & x_59091;
assign x_59093 = x_27804 & x_27805;
assign x_59094 = x_27806 & x_27807;
assign x_59095 = x_59093 & x_59094;
assign x_59096 = x_27808 & x_27809;
assign x_59097 = x_27810 & x_27811;
assign x_59098 = x_59096 & x_59097;
assign x_59099 = x_59095 & x_59098;
assign x_59100 = x_59092 & x_59099;
assign x_59101 = x_59085 & x_59100;
assign x_59102 = x_59071 & x_59101;
assign x_59103 = x_27813 & x_27814;
assign x_59104 = x_27812 & x_59103;
assign x_59105 = x_27815 & x_27816;
assign x_59106 = x_27817 & x_27818;
assign x_59107 = x_59105 & x_59106;
assign x_59108 = x_59104 & x_59107;
assign x_59109 = x_27819 & x_27820;
assign x_59110 = x_27821 & x_27822;
assign x_59111 = x_59109 & x_59110;
assign x_59112 = x_27823 & x_27824;
assign x_59113 = x_27825 & x_27826;
assign x_59114 = x_59112 & x_59113;
assign x_59115 = x_59111 & x_59114;
assign x_59116 = x_59108 & x_59115;
assign x_59117 = x_27827 & x_27828;
assign x_59118 = x_27829 & x_27830;
assign x_59119 = x_59117 & x_59118;
assign x_59120 = x_27831 & x_27832;
assign x_59121 = x_27833 & x_27834;
assign x_59122 = x_59120 & x_59121;
assign x_59123 = x_59119 & x_59122;
assign x_59124 = x_27835 & x_27836;
assign x_59125 = x_27837 & x_27838;
assign x_59126 = x_59124 & x_59125;
assign x_59127 = x_27839 & x_27840;
assign x_59128 = x_27841 & x_27842;
assign x_59129 = x_59127 & x_59128;
assign x_59130 = x_59126 & x_59129;
assign x_59131 = x_59123 & x_59130;
assign x_59132 = x_59116 & x_59131;
assign x_59133 = x_27844 & x_27845;
assign x_59134 = x_27843 & x_59133;
assign x_59135 = x_27846 & x_27847;
assign x_59136 = x_27848 & x_27849;
assign x_59137 = x_59135 & x_59136;
assign x_59138 = x_59134 & x_59137;
assign x_59139 = x_27850 & x_27851;
assign x_59140 = x_27852 & x_27853;
assign x_59141 = x_59139 & x_59140;
assign x_59142 = x_27854 & x_27855;
assign x_59143 = x_27856 & x_27857;
assign x_59144 = x_59142 & x_59143;
assign x_59145 = x_59141 & x_59144;
assign x_59146 = x_59138 & x_59145;
assign x_59147 = x_27858 & x_27859;
assign x_59148 = x_27860 & x_27861;
assign x_59149 = x_59147 & x_59148;
assign x_59150 = x_27862 & x_27863;
assign x_59151 = x_27864 & x_27865;
assign x_59152 = x_59150 & x_59151;
assign x_59153 = x_59149 & x_59152;
assign x_59154 = x_27866 & x_27867;
assign x_59155 = x_27868 & x_27869;
assign x_59156 = x_59154 & x_59155;
assign x_59157 = x_27870 & x_27871;
assign x_59158 = x_27872 & x_27873;
assign x_59159 = x_59157 & x_59158;
assign x_59160 = x_59156 & x_59159;
assign x_59161 = x_59153 & x_59160;
assign x_59162 = x_59146 & x_59161;
assign x_59163 = x_59132 & x_59162;
assign x_59164 = x_59102 & x_59163;
assign x_59165 = x_59042 & x_59164;
assign x_59166 = x_58921 & x_59165;
assign x_59167 = x_27875 & x_27876;
assign x_59168 = x_27874 & x_59167;
assign x_59169 = x_27877 & x_27878;
assign x_59170 = x_27879 & x_27880;
assign x_59171 = x_59169 & x_59170;
assign x_59172 = x_59168 & x_59171;
assign x_59173 = x_27881 & x_27882;
assign x_59174 = x_27883 & x_27884;
assign x_59175 = x_59173 & x_59174;
assign x_59176 = x_27885 & x_27886;
assign x_59177 = x_27887 & x_27888;
assign x_59178 = x_59176 & x_59177;
assign x_59179 = x_59175 & x_59178;
assign x_59180 = x_59172 & x_59179;
assign x_59181 = x_27890 & x_27891;
assign x_59182 = x_27889 & x_59181;
assign x_59183 = x_27892 & x_27893;
assign x_59184 = x_27894 & x_27895;
assign x_59185 = x_59183 & x_59184;
assign x_59186 = x_59182 & x_59185;
assign x_59187 = x_27896 & x_27897;
assign x_59188 = x_27898 & x_27899;
assign x_59189 = x_59187 & x_59188;
assign x_59190 = x_27900 & x_27901;
assign x_59191 = x_27902 & x_27903;
assign x_59192 = x_59190 & x_59191;
assign x_59193 = x_59189 & x_59192;
assign x_59194 = x_59186 & x_59193;
assign x_59195 = x_59180 & x_59194;
assign x_59196 = x_27905 & x_27906;
assign x_59197 = x_27904 & x_59196;
assign x_59198 = x_27907 & x_27908;
assign x_59199 = x_27909 & x_27910;
assign x_59200 = x_59198 & x_59199;
assign x_59201 = x_59197 & x_59200;
assign x_59202 = x_27911 & x_27912;
assign x_59203 = x_27913 & x_27914;
assign x_59204 = x_59202 & x_59203;
assign x_59205 = x_27915 & x_27916;
assign x_59206 = x_27917 & x_27918;
assign x_59207 = x_59205 & x_59206;
assign x_59208 = x_59204 & x_59207;
assign x_59209 = x_59201 & x_59208;
assign x_59210 = x_27919 & x_27920;
assign x_59211 = x_27921 & x_27922;
assign x_59212 = x_59210 & x_59211;
assign x_59213 = x_27923 & x_27924;
assign x_59214 = x_27925 & x_27926;
assign x_59215 = x_59213 & x_59214;
assign x_59216 = x_59212 & x_59215;
assign x_59217 = x_27927 & x_27928;
assign x_59218 = x_27929 & x_27930;
assign x_59219 = x_59217 & x_59218;
assign x_59220 = x_27931 & x_27932;
assign x_59221 = x_27933 & x_27934;
assign x_59222 = x_59220 & x_59221;
assign x_59223 = x_59219 & x_59222;
assign x_59224 = x_59216 & x_59223;
assign x_59225 = x_59209 & x_59224;
assign x_59226 = x_59195 & x_59225;
assign x_59227 = x_27936 & x_27937;
assign x_59228 = x_27935 & x_59227;
assign x_59229 = x_27938 & x_27939;
assign x_59230 = x_27940 & x_27941;
assign x_59231 = x_59229 & x_59230;
assign x_59232 = x_59228 & x_59231;
assign x_59233 = x_27942 & x_27943;
assign x_59234 = x_27944 & x_27945;
assign x_59235 = x_59233 & x_59234;
assign x_59236 = x_27946 & x_27947;
assign x_59237 = x_27948 & x_27949;
assign x_59238 = x_59236 & x_59237;
assign x_59239 = x_59235 & x_59238;
assign x_59240 = x_59232 & x_59239;
assign x_59241 = x_27951 & x_27952;
assign x_59242 = x_27950 & x_59241;
assign x_59243 = x_27953 & x_27954;
assign x_59244 = x_27955 & x_27956;
assign x_59245 = x_59243 & x_59244;
assign x_59246 = x_59242 & x_59245;
assign x_59247 = x_27957 & x_27958;
assign x_59248 = x_27959 & x_27960;
assign x_59249 = x_59247 & x_59248;
assign x_59250 = x_27961 & x_27962;
assign x_59251 = x_27963 & x_27964;
assign x_59252 = x_59250 & x_59251;
assign x_59253 = x_59249 & x_59252;
assign x_59254 = x_59246 & x_59253;
assign x_59255 = x_59240 & x_59254;
assign x_59256 = x_27966 & x_27967;
assign x_59257 = x_27965 & x_59256;
assign x_59258 = x_27968 & x_27969;
assign x_59259 = x_27970 & x_27971;
assign x_59260 = x_59258 & x_59259;
assign x_59261 = x_59257 & x_59260;
assign x_59262 = x_27972 & x_27973;
assign x_59263 = x_27974 & x_27975;
assign x_59264 = x_59262 & x_59263;
assign x_59265 = x_27976 & x_27977;
assign x_59266 = x_27978 & x_27979;
assign x_59267 = x_59265 & x_59266;
assign x_59268 = x_59264 & x_59267;
assign x_59269 = x_59261 & x_59268;
assign x_59270 = x_27980 & x_27981;
assign x_59271 = x_27982 & x_27983;
assign x_59272 = x_59270 & x_59271;
assign x_59273 = x_27984 & x_27985;
assign x_59274 = x_27986 & x_27987;
assign x_59275 = x_59273 & x_59274;
assign x_59276 = x_59272 & x_59275;
assign x_59277 = x_27988 & x_27989;
assign x_59278 = x_27990 & x_27991;
assign x_59279 = x_59277 & x_59278;
assign x_59280 = x_27992 & x_27993;
assign x_59281 = x_27994 & x_27995;
assign x_59282 = x_59280 & x_59281;
assign x_59283 = x_59279 & x_59282;
assign x_59284 = x_59276 & x_59283;
assign x_59285 = x_59269 & x_59284;
assign x_59286 = x_59255 & x_59285;
assign x_59287 = x_59226 & x_59286;
assign x_59288 = x_27997 & x_27998;
assign x_59289 = x_27996 & x_59288;
assign x_59290 = x_27999 & x_28000;
assign x_59291 = x_28001 & x_28002;
assign x_59292 = x_59290 & x_59291;
assign x_59293 = x_59289 & x_59292;
assign x_59294 = x_28003 & x_28004;
assign x_59295 = x_28005 & x_28006;
assign x_59296 = x_59294 & x_59295;
assign x_59297 = x_28007 & x_28008;
assign x_59298 = x_28009 & x_28010;
assign x_59299 = x_59297 & x_59298;
assign x_59300 = x_59296 & x_59299;
assign x_59301 = x_59293 & x_59300;
assign x_59302 = x_28012 & x_28013;
assign x_59303 = x_28011 & x_59302;
assign x_59304 = x_28014 & x_28015;
assign x_59305 = x_28016 & x_28017;
assign x_59306 = x_59304 & x_59305;
assign x_59307 = x_59303 & x_59306;
assign x_59308 = x_28018 & x_28019;
assign x_59309 = x_28020 & x_28021;
assign x_59310 = x_59308 & x_59309;
assign x_59311 = x_28022 & x_28023;
assign x_59312 = x_28024 & x_28025;
assign x_59313 = x_59311 & x_59312;
assign x_59314 = x_59310 & x_59313;
assign x_59315 = x_59307 & x_59314;
assign x_59316 = x_59301 & x_59315;
assign x_59317 = x_28027 & x_28028;
assign x_59318 = x_28026 & x_59317;
assign x_59319 = x_28029 & x_28030;
assign x_59320 = x_28031 & x_28032;
assign x_59321 = x_59319 & x_59320;
assign x_59322 = x_59318 & x_59321;
assign x_59323 = x_28033 & x_28034;
assign x_59324 = x_28035 & x_28036;
assign x_59325 = x_59323 & x_59324;
assign x_59326 = x_28037 & x_28038;
assign x_59327 = x_28039 & x_28040;
assign x_59328 = x_59326 & x_59327;
assign x_59329 = x_59325 & x_59328;
assign x_59330 = x_59322 & x_59329;
assign x_59331 = x_28041 & x_28042;
assign x_59332 = x_28043 & x_28044;
assign x_59333 = x_59331 & x_59332;
assign x_59334 = x_28045 & x_28046;
assign x_59335 = x_28047 & x_28048;
assign x_59336 = x_59334 & x_59335;
assign x_59337 = x_59333 & x_59336;
assign x_59338 = x_28049 & x_28050;
assign x_59339 = x_28051 & x_28052;
assign x_59340 = x_59338 & x_59339;
assign x_59341 = x_28053 & x_28054;
assign x_59342 = x_28055 & x_28056;
assign x_59343 = x_59341 & x_59342;
assign x_59344 = x_59340 & x_59343;
assign x_59345 = x_59337 & x_59344;
assign x_59346 = x_59330 & x_59345;
assign x_59347 = x_59316 & x_59346;
assign x_59348 = x_28058 & x_28059;
assign x_59349 = x_28057 & x_59348;
assign x_59350 = x_28060 & x_28061;
assign x_59351 = x_28062 & x_28063;
assign x_59352 = x_59350 & x_59351;
assign x_59353 = x_59349 & x_59352;
assign x_59354 = x_28064 & x_28065;
assign x_59355 = x_28066 & x_28067;
assign x_59356 = x_59354 & x_59355;
assign x_59357 = x_28068 & x_28069;
assign x_59358 = x_28070 & x_28071;
assign x_59359 = x_59357 & x_59358;
assign x_59360 = x_59356 & x_59359;
assign x_59361 = x_59353 & x_59360;
assign x_59362 = x_28073 & x_28074;
assign x_59363 = x_28072 & x_59362;
assign x_59364 = x_28075 & x_28076;
assign x_59365 = x_28077 & x_28078;
assign x_59366 = x_59364 & x_59365;
assign x_59367 = x_59363 & x_59366;
assign x_59368 = x_28079 & x_28080;
assign x_59369 = x_28081 & x_28082;
assign x_59370 = x_59368 & x_59369;
assign x_59371 = x_28083 & x_28084;
assign x_59372 = x_28085 & x_28086;
assign x_59373 = x_59371 & x_59372;
assign x_59374 = x_59370 & x_59373;
assign x_59375 = x_59367 & x_59374;
assign x_59376 = x_59361 & x_59375;
assign x_59377 = x_28088 & x_28089;
assign x_59378 = x_28087 & x_59377;
assign x_59379 = x_28090 & x_28091;
assign x_59380 = x_28092 & x_28093;
assign x_59381 = x_59379 & x_59380;
assign x_59382 = x_59378 & x_59381;
assign x_59383 = x_28094 & x_28095;
assign x_59384 = x_28096 & x_28097;
assign x_59385 = x_59383 & x_59384;
assign x_59386 = x_28098 & x_28099;
assign x_59387 = x_28100 & x_28101;
assign x_59388 = x_59386 & x_59387;
assign x_59389 = x_59385 & x_59388;
assign x_59390 = x_59382 & x_59389;
assign x_59391 = x_28102 & x_28103;
assign x_59392 = x_28104 & x_28105;
assign x_59393 = x_59391 & x_59392;
assign x_59394 = x_28106 & x_28107;
assign x_59395 = x_28108 & x_28109;
assign x_59396 = x_59394 & x_59395;
assign x_59397 = x_59393 & x_59396;
assign x_59398 = x_28110 & x_28111;
assign x_59399 = x_28112 & x_28113;
assign x_59400 = x_59398 & x_59399;
assign x_59401 = x_28114 & x_28115;
assign x_59402 = x_28116 & x_28117;
assign x_59403 = x_59401 & x_59402;
assign x_59404 = x_59400 & x_59403;
assign x_59405 = x_59397 & x_59404;
assign x_59406 = x_59390 & x_59405;
assign x_59407 = x_59376 & x_59406;
assign x_59408 = x_59347 & x_59407;
assign x_59409 = x_59287 & x_59408;
assign x_59410 = x_28119 & x_28120;
assign x_59411 = x_28118 & x_59410;
assign x_59412 = x_28121 & x_28122;
assign x_59413 = x_28123 & x_28124;
assign x_59414 = x_59412 & x_59413;
assign x_59415 = x_59411 & x_59414;
assign x_59416 = x_28125 & x_28126;
assign x_59417 = x_28127 & x_28128;
assign x_59418 = x_59416 & x_59417;
assign x_59419 = x_28129 & x_28130;
assign x_59420 = x_28131 & x_28132;
assign x_59421 = x_59419 & x_59420;
assign x_59422 = x_59418 & x_59421;
assign x_59423 = x_59415 & x_59422;
assign x_59424 = x_28134 & x_28135;
assign x_59425 = x_28133 & x_59424;
assign x_59426 = x_28136 & x_28137;
assign x_59427 = x_28138 & x_28139;
assign x_59428 = x_59426 & x_59427;
assign x_59429 = x_59425 & x_59428;
assign x_59430 = x_28140 & x_28141;
assign x_59431 = x_28142 & x_28143;
assign x_59432 = x_59430 & x_59431;
assign x_59433 = x_28144 & x_28145;
assign x_59434 = x_28146 & x_28147;
assign x_59435 = x_59433 & x_59434;
assign x_59436 = x_59432 & x_59435;
assign x_59437 = x_59429 & x_59436;
assign x_59438 = x_59423 & x_59437;
assign x_59439 = x_28149 & x_28150;
assign x_59440 = x_28148 & x_59439;
assign x_59441 = x_28151 & x_28152;
assign x_59442 = x_28153 & x_28154;
assign x_59443 = x_59441 & x_59442;
assign x_59444 = x_59440 & x_59443;
assign x_59445 = x_28155 & x_28156;
assign x_59446 = x_28157 & x_28158;
assign x_59447 = x_59445 & x_59446;
assign x_59448 = x_28159 & x_28160;
assign x_59449 = x_28161 & x_28162;
assign x_59450 = x_59448 & x_59449;
assign x_59451 = x_59447 & x_59450;
assign x_59452 = x_59444 & x_59451;
assign x_59453 = x_28163 & x_28164;
assign x_59454 = x_28165 & x_28166;
assign x_59455 = x_59453 & x_59454;
assign x_59456 = x_28167 & x_28168;
assign x_59457 = x_28169 & x_28170;
assign x_59458 = x_59456 & x_59457;
assign x_59459 = x_59455 & x_59458;
assign x_59460 = x_28171 & x_28172;
assign x_59461 = x_28173 & x_28174;
assign x_59462 = x_59460 & x_59461;
assign x_59463 = x_28175 & x_28176;
assign x_59464 = x_28177 & x_28178;
assign x_59465 = x_59463 & x_59464;
assign x_59466 = x_59462 & x_59465;
assign x_59467 = x_59459 & x_59466;
assign x_59468 = x_59452 & x_59467;
assign x_59469 = x_59438 & x_59468;
assign x_59470 = x_28180 & x_28181;
assign x_59471 = x_28179 & x_59470;
assign x_59472 = x_28182 & x_28183;
assign x_59473 = x_28184 & x_28185;
assign x_59474 = x_59472 & x_59473;
assign x_59475 = x_59471 & x_59474;
assign x_59476 = x_28186 & x_28187;
assign x_59477 = x_28188 & x_28189;
assign x_59478 = x_59476 & x_59477;
assign x_59479 = x_28190 & x_28191;
assign x_59480 = x_28192 & x_28193;
assign x_59481 = x_59479 & x_59480;
assign x_59482 = x_59478 & x_59481;
assign x_59483 = x_59475 & x_59482;
assign x_59484 = x_28195 & x_28196;
assign x_59485 = x_28194 & x_59484;
assign x_59486 = x_28197 & x_28198;
assign x_59487 = x_28199 & x_28200;
assign x_59488 = x_59486 & x_59487;
assign x_59489 = x_59485 & x_59488;
assign x_59490 = x_28201 & x_28202;
assign x_59491 = x_28203 & x_28204;
assign x_59492 = x_59490 & x_59491;
assign x_59493 = x_28205 & x_28206;
assign x_59494 = x_28207 & x_28208;
assign x_59495 = x_59493 & x_59494;
assign x_59496 = x_59492 & x_59495;
assign x_59497 = x_59489 & x_59496;
assign x_59498 = x_59483 & x_59497;
assign x_59499 = x_28210 & x_28211;
assign x_59500 = x_28209 & x_59499;
assign x_59501 = x_28212 & x_28213;
assign x_59502 = x_28214 & x_28215;
assign x_59503 = x_59501 & x_59502;
assign x_59504 = x_59500 & x_59503;
assign x_59505 = x_28216 & x_28217;
assign x_59506 = x_28218 & x_28219;
assign x_59507 = x_59505 & x_59506;
assign x_59508 = x_28220 & x_28221;
assign x_59509 = x_28222 & x_28223;
assign x_59510 = x_59508 & x_59509;
assign x_59511 = x_59507 & x_59510;
assign x_59512 = x_59504 & x_59511;
assign x_59513 = x_28224 & x_28225;
assign x_59514 = x_28226 & x_28227;
assign x_59515 = x_59513 & x_59514;
assign x_59516 = x_28228 & x_28229;
assign x_59517 = x_28230 & x_28231;
assign x_59518 = x_59516 & x_59517;
assign x_59519 = x_59515 & x_59518;
assign x_59520 = x_28232 & x_28233;
assign x_59521 = x_28234 & x_28235;
assign x_59522 = x_59520 & x_59521;
assign x_59523 = x_28236 & x_28237;
assign x_59524 = x_28238 & x_28239;
assign x_59525 = x_59523 & x_59524;
assign x_59526 = x_59522 & x_59525;
assign x_59527 = x_59519 & x_59526;
assign x_59528 = x_59512 & x_59527;
assign x_59529 = x_59498 & x_59528;
assign x_59530 = x_59469 & x_59529;
assign x_59531 = x_28241 & x_28242;
assign x_59532 = x_28240 & x_59531;
assign x_59533 = x_28243 & x_28244;
assign x_59534 = x_28245 & x_28246;
assign x_59535 = x_59533 & x_59534;
assign x_59536 = x_59532 & x_59535;
assign x_59537 = x_28247 & x_28248;
assign x_59538 = x_28249 & x_28250;
assign x_59539 = x_59537 & x_59538;
assign x_59540 = x_28251 & x_28252;
assign x_59541 = x_28253 & x_28254;
assign x_59542 = x_59540 & x_59541;
assign x_59543 = x_59539 & x_59542;
assign x_59544 = x_59536 & x_59543;
assign x_59545 = x_28256 & x_28257;
assign x_59546 = x_28255 & x_59545;
assign x_59547 = x_28258 & x_28259;
assign x_59548 = x_28260 & x_28261;
assign x_59549 = x_59547 & x_59548;
assign x_59550 = x_59546 & x_59549;
assign x_59551 = x_28262 & x_28263;
assign x_59552 = x_28264 & x_28265;
assign x_59553 = x_59551 & x_59552;
assign x_59554 = x_28266 & x_28267;
assign x_59555 = x_28268 & x_28269;
assign x_59556 = x_59554 & x_59555;
assign x_59557 = x_59553 & x_59556;
assign x_59558 = x_59550 & x_59557;
assign x_59559 = x_59544 & x_59558;
assign x_59560 = x_28271 & x_28272;
assign x_59561 = x_28270 & x_59560;
assign x_59562 = x_28273 & x_28274;
assign x_59563 = x_28275 & x_28276;
assign x_59564 = x_59562 & x_59563;
assign x_59565 = x_59561 & x_59564;
assign x_59566 = x_28277 & x_28278;
assign x_59567 = x_28279 & x_28280;
assign x_59568 = x_59566 & x_59567;
assign x_59569 = x_28281 & x_28282;
assign x_59570 = x_28283 & x_28284;
assign x_59571 = x_59569 & x_59570;
assign x_59572 = x_59568 & x_59571;
assign x_59573 = x_59565 & x_59572;
assign x_59574 = x_28285 & x_28286;
assign x_59575 = x_28287 & x_28288;
assign x_59576 = x_59574 & x_59575;
assign x_59577 = x_28289 & x_28290;
assign x_59578 = x_28291 & x_28292;
assign x_59579 = x_59577 & x_59578;
assign x_59580 = x_59576 & x_59579;
assign x_59581 = x_28293 & x_28294;
assign x_59582 = x_28295 & x_28296;
assign x_59583 = x_59581 & x_59582;
assign x_59584 = x_28297 & x_28298;
assign x_59585 = x_28299 & x_28300;
assign x_59586 = x_59584 & x_59585;
assign x_59587 = x_59583 & x_59586;
assign x_59588 = x_59580 & x_59587;
assign x_59589 = x_59573 & x_59588;
assign x_59590 = x_59559 & x_59589;
assign x_59591 = x_28302 & x_28303;
assign x_59592 = x_28301 & x_59591;
assign x_59593 = x_28304 & x_28305;
assign x_59594 = x_28306 & x_28307;
assign x_59595 = x_59593 & x_59594;
assign x_59596 = x_59592 & x_59595;
assign x_59597 = x_28308 & x_28309;
assign x_59598 = x_28310 & x_28311;
assign x_59599 = x_59597 & x_59598;
assign x_59600 = x_28312 & x_28313;
assign x_59601 = x_28314 & x_28315;
assign x_59602 = x_59600 & x_59601;
assign x_59603 = x_59599 & x_59602;
assign x_59604 = x_59596 & x_59603;
assign x_59605 = x_28316 & x_28317;
assign x_59606 = x_28318 & x_28319;
assign x_59607 = x_59605 & x_59606;
assign x_59608 = x_28320 & x_28321;
assign x_59609 = x_28322 & x_28323;
assign x_59610 = x_59608 & x_59609;
assign x_59611 = x_59607 & x_59610;
assign x_59612 = x_28324 & x_28325;
assign x_59613 = x_28326 & x_28327;
assign x_59614 = x_59612 & x_59613;
assign x_59615 = x_28328 & x_28329;
assign x_59616 = x_28330 & x_28331;
assign x_59617 = x_59615 & x_59616;
assign x_59618 = x_59614 & x_59617;
assign x_59619 = x_59611 & x_59618;
assign x_59620 = x_59604 & x_59619;
assign x_59621 = x_28333 & x_28334;
assign x_59622 = x_28332 & x_59621;
assign x_59623 = x_28335 & x_28336;
assign x_59624 = x_28337 & x_28338;
assign x_59625 = x_59623 & x_59624;
assign x_59626 = x_59622 & x_59625;
assign x_59627 = x_28339 & x_28340;
assign x_59628 = x_28341 & x_28342;
assign x_59629 = x_59627 & x_59628;
assign x_59630 = x_28343 & x_28344;
assign x_59631 = x_28345 & x_28346;
assign x_59632 = x_59630 & x_59631;
assign x_59633 = x_59629 & x_59632;
assign x_59634 = x_59626 & x_59633;
assign x_59635 = x_28347 & x_28348;
assign x_59636 = x_28349 & x_28350;
assign x_59637 = x_59635 & x_59636;
assign x_59638 = x_28351 & x_28352;
assign x_59639 = x_28353 & x_28354;
assign x_59640 = x_59638 & x_59639;
assign x_59641 = x_59637 & x_59640;
assign x_59642 = x_28355 & x_28356;
assign x_59643 = x_28357 & x_28358;
assign x_59644 = x_59642 & x_59643;
assign x_59645 = x_28359 & x_28360;
assign x_59646 = x_28361 & x_28362;
assign x_59647 = x_59645 & x_59646;
assign x_59648 = x_59644 & x_59647;
assign x_59649 = x_59641 & x_59648;
assign x_59650 = x_59634 & x_59649;
assign x_59651 = x_59620 & x_59650;
assign x_59652 = x_59590 & x_59651;
assign x_59653 = x_59530 & x_59652;
assign x_59654 = x_59409 & x_59653;
assign x_59655 = x_59166 & x_59654;
assign x_59656 = x_28364 & x_28365;
assign x_59657 = x_28363 & x_59656;
assign x_59658 = x_28366 & x_28367;
assign x_59659 = x_28368 & x_28369;
assign x_59660 = x_59658 & x_59659;
assign x_59661 = x_59657 & x_59660;
assign x_59662 = x_28370 & x_28371;
assign x_59663 = x_28372 & x_28373;
assign x_59664 = x_59662 & x_59663;
assign x_59665 = x_28374 & x_28375;
assign x_59666 = x_28376 & x_28377;
assign x_59667 = x_59665 & x_59666;
assign x_59668 = x_59664 & x_59667;
assign x_59669 = x_59661 & x_59668;
assign x_59670 = x_28379 & x_28380;
assign x_59671 = x_28378 & x_59670;
assign x_59672 = x_28381 & x_28382;
assign x_59673 = x_28383 & x_28384;
assign x_59674 = x_59672 & x_59673;
assign x_59675 = x_59671 & x_59674;
assign x_59676 = x_28385 & x_28386;
assign x_59677 = x_28387 & x_28388;
assign x_59678 = x_59676 & x_59677;
assign x_59679 = x_28389 & x_28390;
assign x_59680 = x_28391 & x_28392;
assign x_59681 = x_59679 & x_59680;
assign x_59682 = x_59678 & x_59681;
assign x_59683 = x_59675 & x_59682;
assign x_59684 = x_59669 & x_59683;
assign x_59685 = x_28394 & x_28395;
assign x_59686 = x_28393 & x_59685;
assign x_59687 = x_28396 & x_28397;
assign x_59688 = x_28398 & x_28399;
assign x_59689 = x_59687 & x_59688;
assign x_59690 = x_59686 & x_59689;
assign x_59691 = x_28400 & x_28401;
assign x_59692 = x_28402 & x_28403;
assign x_59693 = x_59691 & x_59692;
assign x_59694 = x_28404 & x_28405;
assign x_59695 = x_28406 & x_28407;
assign x_59696 = x_59694 & x_59695;
assign x_59697 = x_59693 & x_59696;
assign x_59698 = x_59690 & x_59697;
assign x_59699 = x_28408 & x_28409;
assign x_59700 = x_28410 & x_28411;
assign x_59701 = x_59699 & x_59700;
assign x_59702 = x_28412 & x_28413;
assign x_59703 = x_28414 & x_28415;
assign x_59704 = x_59702 & x_59703;
assign x_59705 = x_59701 & x_59704;
assign x_59706 = x_28416 & x_28417;
assign x_59707 = x_28418 & x_28419;
assign x_59708 = x_59706 & x_59707;
assign x_59709 = x_28420 & x_28421;
assign x_59710 = x_28422 & x_28423;
assign x_59711 = x_59709 & x_59710;
assign x_59712 = x_59708 & x_59711;
assign x_59713 = x_59705 & x_59712;
assign x_59714 = x_59698 & x_59713;
assign x_59715 = x_59684 & x_59714;
assign x_59716 = x_28425 & x_28426;
assign x_59717 = x_28424 & x_59716;
assign x_59718 = x_28427 & x_28428;
assign x_59719 = x_28429 & x_28430;
assign x_59720 = x_59718 & x_59719;
assign x_59721 = x_59717 & x_59720;
assign x_59722 = x_28431 & x_28432;
assign x_59723 = x_28433 & x_28434;
assign x_59724 = x_59722 & x_59723;
assign x_59725 = x_28435 & x_28436;
assign x_59726 = x_28437 & x_28438;
assign x_59727 = x_59725 & x_59726;
assign x_59728 = x_59724 & x_59727;
assign x_59729 = x_59721 & x_59728;
assign x_59730 = x_28440 & x_28441;
assign x_59731 = x_28439 & x_59730;
assign x_59732 = x_28442 & x_28443;
assign x_59733 = x_28444 & x_28445;
assign x_59734 = x_59732 & x_59733;
assign x_59735 = x_59731 & x_59734;
assign x_59736 = x_28446 & x_28447;
assign x_59737 = x_28448 & x_28449;
assign x_59738 = x_59736 & x_59737;
assign x_59739 = x_28450 & x_28451;
assign x_59740 = x_28452 & x_28453;
assign x_59741 = x_59739 & x_59740;
assign x_59742 = x_59738 & x_59741;
assign x_59743 = x_59735 & x_59742;
assign x_59744 = x_59729 & x_59743;
assign x_59745 = x_28455 & x_28456;
assign x_59746 = x_28454 & x_59745;
assign x_59747 = x_28457 & x_28458;
assign x_59748 = x_28459 & x_28460;
assign x_59749 = x_59747 & x_59748;
assign x_59750 = x_59746 & x_59749;
assign x_59751 = x_28461 & x_28462;
assign x_59752 = x_28463 & x_28464;
assign x_59753 = x_59751 & x_59752;
assign x_59754 = x_28465 & x_28466;
assign x_59755 = x_28467 & x_28468;
assign x_59756 = x_59754 & x_59755;
assign x_59757 = x_59753 & x_59756;
assign x_59758 = x_59750 & x_59757;
assign x_59759 = x_28469 & x_28470;
assign x_59760 = x_28471 & x_28472;
assign x_59761 = x_59759 & x_59760;
assign x_59762 = x_28473 & x_28474;
assign x_59763 = x_28475 & x_28476;
assign x_59764 = x_59762 & x_59763;
assign x_59765 = x_59761 & x_59764;
assign x_59766 = x_28477 & x_28478;
assign x_59767 = x_28479 & x_28480;
assign x_59768 = x_59766 & x_59767;
assign x_59769 = x_28481 & x_28482;
assign x_59770 = x_28483 & x_28484;
assign x_59771 = x_59769 & x_59770;
assign x_59772 = x_59768 & x_59771;
assign x_59773 = x_59765 & x_59772;
assign x_59774 = x_59758 & x_59773;
assign x_59775 = x_59744 & x_59774;
assign x_59776 = x_59715 & x_59775;
assign x_59777 = x_28486 & x_28487;
assign x_59778 = x_28485 & x_59777;
assign x_59779 = x_28488 & x_28489;
assign x_59780 = x_28490 & x_28491;
assign x_59781 = x_59779 & x_59780;
assign x_59782 = x_59778 & x_59781;
assign x_59783 = x_28492 & x_28493;
assign x_59784 = x_28494 & x_28495;
assign x_59785 = x_59783 & x_59784;
assign x_59786 = x_28496 & x_28497;
assign x_59787 = x_28498 & x_28499;
assign x_59788 = x_59786 & x_59787;
assign x_59789 = x_59785 & x_59788;
assign x_59790 = x_59782 & x_59789;
assign x_59791 = x_28501 & x_28502;
assign x_59792 = x_28500 & x_59791;
assign x_59793 = x_28503 & x_28504;
assign x_59794 = x_28505 & x_28506;
assign x_59795 = x_59793 & x_59794;
assign x_59796 = x_59792 & x_59795;
assign x_59797 = x_28507 & x_28508;
assign x_59798 = x_28509 & x_28510;
assign x_59799 = x_59797 & x_59798;
assign x_59800 = x_28511 & x_28512;
assign x_59801 = x_28513 & x_28514;
assign x_59802 = x_59800 & x_59801;
assign x_59803 = x_59799 & x_59802;
assign x_59804 = x_59796 & x_59803;
assign x_59805 = x_59790 & x_59804;
assign x_59806 = x_28516 & x_28517;
assign x_59807 = x_28515 & x_59806;
assign x_59808 = x_28518 & x_28519;
assign x_59809 = x_28520 & x_28521;
assign x_59810 = x_59808 & x_59809;
assign x_59811 = x_59807 & x_59810;
assign x_59812 = x_28522 & x_28523;
assign x_59813 = x_28524 & x_28525;
assign x_59814 = x_59812 & x_59813;
assign x_59815 = x_28526 & x_28527;
assign x_59816 = x_28528 & x_28529;
assign x_59817 = x_59815 & x_59816;
assign x_59818 = x_59814 & x_59817;
assign x_59819 = x_59811 & x_59818;
assign x_59820 = x_28530 & x_28531;
assign x_59821 = x_28532 & x_28533;
assign x_59822 = x_59820 & x_59821;
assign x_59823 = x_28534 & x_28535;
assign x_59824 = x_28536 & x_28537;
assign x_59825 = x_59823 & x_59824;
assign x_59826 = x_59822 & x_59825;
assign x_59827 = x_28538 & x_28539;
assign x_59828 = x_28540 & x_28541;
assign x_59829 = x_59827 & x_59828;
assign x_59830 = x_28542 & x_28543;
assign x_59831 = x_28544 & x_28545;
assign x_59832 = x_59830 & x_59831;
assign x_59833 = x_59829 & x_59832;
assign x_59834 = x_59826 & x_59833;
assign x_59835 = x_59819 & x_59834;
assign x_59836 = x_59805 & x_59835;
assign x_59837 = x_28547 & x_28548;
assign x_59838 = x_28546 & x_59837;
assign x_59839 = x_28549 & x_28550;
assign x_59840 = x_28551 & x_28552;
assign x_59841 = x_59839 & x_59840;
assign x_59842 = x_59838 & x_59841;
assign x_59843 = x_28553 & x_28554;
assign x_59844 = x_28555 & x_28556;
assign x_59845 = x_59843 & x_59844;
assign x_59846 = x_28557 & x_28558;
assign x_59847 = x_28559 & x_28560;
assign x_59848 = x_59846 & x_59847;
assign x_59849 = x_59845 & x_59848;
assign x_59850 = x_59842 & x_59849;
assign x_59851 = x_28562 & x_28563;
assign x_59852 = x_28561 & x_59851;
assign x_59853 = x_28564 & x_28565;
assign x_59854 = x_28566 & x_28567;
assign x_59855 = x_59853 & x_59854;
assign x_59856 = x_59852 & x_59855;
assign x_59857 = x_28568 & x_28569;
assign x_59858 = x_28570 & x_28571;
assign x_59859 = x_59857 & x_59858;
assign x_59860 = x_28572 & x_28573;
assign x_59861 = x_28574 & x_28575;
assign x_59862 = x_59860 & x_59861;
assign x_59863 = x_59859 & x_59862;
assign x_59864 = x_59856 & x_59863;
assign x_59865 = x_59850 & x_59864;
assign x_59866 = x_28577 & x_28578;
assign x_59867 = x_28576 & x_59866;
assign x_59868 = x_28579 & x_28580;
assign x_59869 = x_28581 & x_28582;
assign x_59870 = x_59868 & x_59869;
assign x_59871 = x_59867 & x_59870;
assign x_59872 = x_28583 & x_28584;
assign x_59873 = x_28585 & x_28586;
assign x_59874 = x_59872 & x_59873;
assign x_59875 = x_28587 & x_28588;
assign x_59876 = x_28589 & x_28590;
assign x_59877 = x_59875 & x_59876;
assign x_59878 = x_59874 & x_59877;
assign x_59879 = x_59871 & x_59878;
assign x_59880 = x_28591 & x_28592;
assign x_59881 = x_28593 & x_28594;
assign x_59882 = x_59880 & x_59881;
assign x_59883 = x_28595 & x_28596;
assign x_59884 = x_28597 & x_28598;
assign x_59885 = x_59883 & x_59884;
assign x_59886 = x_59882 & x_59885;
assign x_59887 = x_28599 & x_28600;
assign x_59888 = x_28601 & x_28602;
assign x_59889 = x_59887 & x_59888;
assign x_59890 = x_28603 & x_28604;
assign x_59891 = x_28605 & x_28606;
assign x_59892 = x_59890 & x_59891;
assign x_59893 = x_59889 & x_59892;
assign x_59894 = x_59886 & x_59893;
assign x_59895 = x_59879 & x_59894;
assign x_59896 = x_59865 & x_59895;
assign x_59897 = x_59836 & x_59896;
assign x_59898 = x_59776 & x_59897;
assign x_59899 = x_28608 & x_28609;
assign x_59900 = x_28607 & x_59899;
assign x_59901 = x_28610 & x_28611;
assign x_59902 = x_28612 & x_28613;
assign x_59903 = x_59901 & x_59902;
assign x_59904 = x_59900 & x_59903;
assign x_59905 = x_28614 & x_28615;
assign x_59906 = x_28616 & x_28617;
assign x_59907 = x_59905 & x_59906;
assign x_59908 = x_28618 & x_28619;
assign x_59909 = x_28620 & x_28621;
assign x_59910 = x_59908 & x_59909;
assign x_59911 = x_59907 & x_59910;
assign x_59912 = x_59904 & x_59911;
assign x_59913 = x_28623 & x_28624;
assign x_59914 = x_28622 & x_59913;
assign x_59915 = x_28625 & x_28626;
assign x_59916 = x_28627 & x_28628;
assign x_59917 = x_59915 & x_59916;
assign x_59918 = x_59914 & x_59917;
assign x_59919 = x_28629 & x_28630;
assign x_59920 = x_28631 & x_28632;
assign x_59921 = x_59919 & x_59920;
assign x_59922 = x_28633 & x_28634;
assign x_59923 = x_28635 & x_28636;
assign x_59924 = x_59922 & x_59923;
assign x_59925 = x_59921 & x_59924;
assign x_59926 = x_59918 & x_59925;
assign x_59927 = x_59912 & x_59926;
assign x_59928 = x_28638 & x_28639;
assign x_59929 = x_28637 & x_59928;
assign x_59930 = x_28640 & x_28641;
assign x_59931 = x_28642 & x_28643;
assign x_59932 = x_59930 & x_59931;
assign x_59933 = x_59929 & x_59932;
assign x_59934 = x_28644 & x_28645;
assign x_59935 = x_28646 & x_28647;
assign x_59936 = x_59934 & x_59935;
assign x_59937 = x_28648 & x_28649;
assign x_59938 = x_28650 & x_28651;
assign x_59939 = x_59937 & x_59938;
assign x_59940 = x_59936 & x_59939;
assign x_59941 = x_59933 & x_59940;
assign x_59942 = x_28652 & x_28653;
assign x_59943 = x_28654 & x_28655;
assign x_59944 = x_59942 & x_59943;
assign x_59945 = x_28656 & x_28657;
assign x_59946 = x_28658 & x_28659;
assign x_59947 = x_59945 & x_59946;
assign x_59948 = x_59944 & x_59947;
assign x_59949 = x_28660 & x_28661;
assign x_59950 = x_28662 & x_28663;
assign x_59951 = x_59949 & x_59950;
assign x_59952 = x_28664 & x_28665;
assign x_59953 = x_28666 & x_28667;
assign x_59954 = x_59952 & x_59953;
assign x_59955 = x_59951 & x_59954;
assign x_59956 = x_59948 & x_59955;
assign x_59957 = x_59941 & x_59956;
assign x_59958 = x_59927 & x_59957;
assign x_59959 = x_28669 & x_28670;
assign x_59960 = x_28668 & x_59959;
assign x_59961 = x_28671 & x_28672;
assign x_59962 = x_28673 & x_28674;
assign x_59963 = x_59961 & x_59962;
assign x_59964 = x_59960 & x_59963;
assign x_59965 = x_28675 & x_28676;
assign x_59966 = x_28677 & x_28678;
assign x_59967 = x_59965 & x_59966;
assign x_59968 = x_28679 & x_28680;
assign x_59969 = x_28681 & x_28682;
assign x_59970 = x_59968 & x_59969;
assign x_59971 = x_59967 & x_59970;
assign x_59972 = x_59964 & x_59971;
assign x_59973 = x_28684 & x_28685;
assign x_59974 = x_28683 & x_59973;
assign x_59975 = x_28686 & x_28687;
assign x_59976 = x_28688 & x_28689;
assign x_59977 = x_59975 & x_59976;
assign x_59978 = x_59974 & x_59977;
assign x_59979 = x_28690 & x_28691;
assign x_59980 = x_28692 & x_28693;
assign x_59981 = x_59979 & x_59980;
assign x_59982 = x_28694 & x_28695;
assign x_59983 = x_28696 & x_28697;
assign x_59984 = x_59982 & x_59983;
assign x_59985 = x_59981 & x_59984;
assign x_59986 = x_59978 & x_59985;
assign x_59987 = x_59972 & x_59986;
assign x_59988 = x_28699 & x_28700;
assign x_59989 = x_28698 & x_59988;
assign x_59990 = x_28701 & x_28702;
assign x_59991 = x_28703 & x_28704;
assign x_59992 = x_59990 & x_59991;
assign x_59993 = x_59989 & x_59992;
assign x_59994 = x_28705 & x_28706;
assign x_59995 = x_28707 & x_28708;
assign x_59996 = x_59994 & x_59995;
assign x_59997 = x_28709 & x_28710;
assign x_59998 = x_28711 & x_28712;
assign x_59999 = x_59997 & x_59998;
assign x_60000 = x_59996 & x_59999;
assign x_60001 = x_59993 & x_60000;
assign x_60002 = x_28713 & x_28714;
assign x_60003 = x_28715 & x_28716;
assign x_60004 = x_60002 & x_60003;
assign x_60005 = x_28717 & x_28718;
assign x_60006 = x_28719 & x_28720;
assign x_60007 = x_60005 & x_60006;
assign x_60008 = x_60004 & x_60007;
assign x_60009 = x_28721 & x_28722;
assign x_60010 = x_28723 & x_28724;
assign x_60011 = x_60009 & x_60010;
assign x_60012 = x_28725 & x_28726;
assign x_60013 = x_28727 & x_28728;
assign x_60014 = x_60012 & x_60013;
assign x_60015 = x_60011 & x_60014;
assign x_60016 = x_60008 & x_60015;
assign x_60017 = x_60001 & x_60016;
assign x_60018 = x_59987 & x_60017;
assign x_60019 = x_59958 & x_60018;
assign x_60020 = x_28730 & x_28731;
assign x_60021 = x_28729 & x_60020;
assign x_60022 = x_28732 & x_28733;
assign x_60023 = x_28734 & x_28735;
assign x_60024 = x_60022 & x_60023;
assign x_60025 = x_60021 & x_60024;
assign x_60026 = x_28736 & x_28737;
assign x_60027 = x_28738 & x_28739;
assign x_60028 = x_60026 & x_60027;
assign x_60029 = x_28740 & x_28741;
assign x_60030 = x_28742 & x_28743;
assign x_60031 = x_60029 & x_60030;
assign x_60032 = x_60028 & x_60031;
assign x_60033 = x_60025 & x_60032;
assign x_60034 = x_28745 & x_28746;
assign x_60035 = x_28744 & x_60034;
assign x_60036 = x_28747 & x_28748;
assign x_60037 = x_28749 & x_28750;
assign x_60038 = x_60036 & x_60037;
assign x_60039 = x_60035 & x_60038;
assign x_60040 = x_28751 & x_28752;
assign x_60041 = x_28753 & x_28754;
assign x_60042 = x_60040 & x_60041;
assign x_60043 = x_28755 & x_28756;
assign x_60044 = x_28757 & x_28758;
assign x_60045 = x_60043 & x_60044;
assign x_60046 = x_60042 & x_60045;
assign x_60047 = x_60039 & x_60046;
assign x_60048 = x_60033 & x_60047;
assign x_60049 = x_28760 & x_28761;
assign x_60050 = x_28759 & x_60049;
assign x_60051 = x_28762 & x_28763;
assign x_60052 = x_28764 & x_28765;
assign x_60053 = x_60051 & x_60052;
assign x_60054 = x_60050 & x_60053;
assign x_60055 = x_28766 & x_28767;
assign x_60056 = x_28768 & x_28769;
assign x_60057 = x_60055 & x_60056;
assign x_60058 = x_28770 & x_28771;
assign x_60059 = x_28772 & x_28773;
assign x_60060 = x_60058 & x_60059;
assign x_60061 = x_60057 & x_60060;
assign x_60062 = x_60054 & x_60061;
assign x_60063 = x_28774 & x_28775;
assign x_60064 = x_28776 & x_28777;
assign x_60065 = x_60063 & x_60064;
assign x_60066 = x_28778 & x_28779;
assign x_60067 = x_28780 & x_28781;
assign x_60068 = x_60066 & x_60067;
assign x_60069 = x_60065 & x_60068;
assign x_60070 = x_28782 & x_28783;
assign x_60071 = x_28784 & x_28785;
assign x_60072 = x_60070 & x_60071;
assign x_60073 = x_28786 & x_28787;
assign x_60074 = x_28788 & x_28789;
assign x_60075 = x_60073 & x_60074;
assign x_60076 = x_60072 & x_60075;
assign x_60077 = x_60069 & x_60076;
assign x_60078 = x_60062 & x_60077;
assign x_60079 = x_60048 & x_60078;
assign x_60080 = x_28791 & x_28792;
assign x_60081 = x_28790 & x_60080;
assign x_60082 = x_28793 & x_28794;
assign x_60083 = x_28795 & x_28796;
assign x_60084 = x_60082 & x_60083;
assign x_60085 = x_60081 & x_60084;
assign x_60086 = x_28797 & x_28798;
assign x_60087 = x_28799 & x_28800;
assign x_60088 = x_60086 & x_60087;
assign x_60089 = x_28801 & x_28802;
assign x_60090 = x_28803 & x_28804;
assign x_60091 = x_60089 & x_60090;
assign x_60092 = x_60088 & x_60091;
assign x_60093 = x_60085 & x_60092;
assign x_60094 = x_28805 & x_28806;
assign x_60095 = x_28807 & x_28808;
assign x_60096 = x_60094 & x_60095;
assign x_60097 = x_28809 & x_28810;
assign x_60098 = x_28811 & x_28812;
assign x_60099 = x_60097 & x_60098;
assign x_60100 = x_60096 & x_60099;
assign x_60101 = x_28813 & x_28814;
assign x_60102 = x_28815 & x_28816;
assign x_60103 = x_60101 & x_60102;
assign x_60104 = x_28817 & x_28818;
assign x_60105 = x_28819 & x_28820;
assign x_60106 = x_60104 & x_60105;
assign x_60107 = x_60103 & x_60106;
assign x_60108 = x_60100 & x_60107;
assign x_60109 = x_60093 & x_60108;
assign x_60110 = x_28822 & x_28823;
assign x_60111 = x_28821 & x_60110;
assign x_60112 = x_28824 & x_28825;
assign x_60113 = x_28826 & x_28827;
assign x_60114 = x_60112 & x_60113;
assign x_60115 = x_60111 & x_60114;
assign x_60116 = x_28828 & x_28829;
assign x_60117 = x_28830 & x_28831;
assign x_60118 = x_60116 & x_60117;
assign x_60119 = x_28832 & x_28833;
assign x_60120 = x_28834 & x_28835;
assign x_60121 = x_60119 & x_60120;
assign x_60122 = x_60118 & x_60121;
assign x_60123 = x_60115 & x_60122;
assign x_60124 = x_28836 & x_28837;
assign x_60125 = x_28838 & x_28839;
assign x_60126 = x_60124 & x_60125;
assign x_60127 = x_28840 & x_28841;
assign x_60128 = x_28842 & x_28843;
assign x_60129 = x_60127 & x_60128;
assign x_60130 = x_60126 & x_60129;
assign x_60131 = x_28844 & x_28845;
assign x_60132 = x_28846 & x_28847;
assign x_60133 = x_60131 & x_60132;
assign x_60134 = x_28848 & x_28849;
assign x_60135 = x_28850 & x_28851;
assign x_60136 = x_60134 & x_60135;
assign x_60137 = x_60133 & x_60136;
assign x_60138 = x_60130 & x_60137;
assign x_60139 = x_60123 & x_60138;
assign x_60140 = x_60109 & x_60139;
assign x_60141 = x_60079 & x_60140;
assign x_60142 = x_60019 & x_60141;
assign x_60143 = x_59898 & x_60142;
assign x_60144 = x_28853 & x_28854;
assign x_60145 = x_28852 & x_60144;
assign x_60146 = x_28855 & x_28856;
assign x_60147 = x_28857 & x_28858;
assign x_60148 = x_60146 & x_60147;
assign x_60149 = x_60145 & x_60148;
assign x_60150 = x_28859 & x_28860;
assign x_60151 = x_28861 & x_28862;
assign x_60152 = x_60150 & x_60151;
assign x_60153 = x_28863 & x_28864;
assign x_60154 = x_28865 & x_28866;
assign x_60155 = x_60153 & x_60154;
assign x_60156 = x_60152 & x_60155;
assign x_60157 = x_60149 & x_60156;
assign x_60158 = x_28868 & x_28869;
assign x_60159 = x_28867 & x_60158;
assign x_60160 = x_28870 & x_28871;
assign x_60161 = x_28872 & x_28873;
assign x_60162 = x_60160 & x_60161;
assign x_60163 = x_60159 & x_60162;
assign x_60164 = x_28874 & x_28875;
assign x_60165 = x_28876 & x_28877;
assign x_60166 = x_60164 & x_60165;
assign x_60167 = x_28878 & x_28879;
assign x_60168 = x_28880 & x_28881;
assign x_60169 = x_60167 & x_60168;
assign x_60170 = x_60166 & x_60169;
assign x_60171 = x_60163 & x_60170;
assign x_60172 = x_60157 & x_60171;
assign x_60173 = x_28883 & x_28884;
assign x_60174 = x_28882 & x_60173;
assign x_60175 = x_28885 & x_28886;
assign x_60176 = x_28887 & x_28888;
assign x_60177 = x_60175 & x_60176;
assign x_60178 = x_60174 & x_60177;
assign x_60179 = x_28889 & x_28890;
assign x_60180 = x_28891 & x_28892;
assign x_60181 = x_60179 & x_60180;
assign x_60182 = x_28893 & x_28894;
assign x_60183 = x_28895 & x_28896;
assign x_60184 = x_60182 & x_60183;
assign x_60185 = x_60181 & x_60184;
assign x_60186 = x_60178 & x_60185;
assign x_60187 = x_28897 & x_28898;
assign x_60188 = x_28899 & x_28900;
assign x_60189 = x_60187 & x_60188;
assign x_60190 = x_28901 & x_28902;
assign x_60191 = x_28903 & x_28904;
assign x_60192 = x_60190 & x_60191;
assign x_60193 = x_60189 & x_60192;
assign x_60194 = x_28905 & x_28906;
assign x_60195 = x_28907 & x_28908;
assign x_60196 = x_60194 & x_60195;
assign x_60197 = x_28909 & x_28910;
assign x_60198 = x_28911 & x_28912;
assign x_60199 = x_60197 & x_60198;
assign x_60200 = x_60196 & x_60199;
assign x_60201 = x_60193 & x_60200;
assign x_60202 = x_60186 & x_60201;
assign x_60203 = x_60172 & x_60202;
assign x_60204 = x_28914 & x_28915;
assign x_60205 = x_28913 & x_60204;
assign x_60206 = x_28916 & x_28917;
assign x_60207 = x_28918 & x_28919;
assign x_60208 = x_60206 & x_60207;
assign x_60209 = x_60205 & x_60208;
assign x_60210 = x_28920 & x_28921;
assign x_60211 = x_28922 & x_28923;
assign x_60212 = x_60210 & x_60211;
assign x_60213 = x_28924 & x_28925;
assign x_60214 = x_28926 & x_28927;
assign x_60215 = x_60213 & x_60214;
assign x_60216 = x_60212 & x_60215;
assign x_60217 = x_60209 & x_60216;
assign x_60218 = x_28929 & x_28930;
assign x_60219 = x_28928 & x_60218;
assign x_60220 = x_28931 & x_28932;
assign x_60221 = x_28933 & x_28934;
assign x_60222 = x_60220 & x_60221;
assign x_60223 = x_60219 & x_60222;
assign x_60224 = x_28935 & x_28936;
assign x_60225 = x_28937 & x_28938;
assign x_60226 = x_60224 & x_60225;
assign x_60227 = x_28939 & x_28940;
assign x_60228 = x_28941 & x_28942;
assign x_60229 = x_60227 & x_60228;
assign x_60230 = x_60226 & x_60229;
assign x_60231 = x_60223 & x_60230;
assign x_60232 = x_60217 & x_60231;
assign x_60233 = x_28944 & x_28945;
assign x_60234 = x_28943 & x_60233;
assign x_60235 = x_28946 & x_28947;
assign x_60236 = x_28948 & x_28949;
assign x_60237 = x_60235 & x_60236;
assign x_60238 = x_60234 & x_60237;
assign x_60239 = x_28950 & x_28951;
assign x_60240 = x_28952 & x_28953;
assign x_60241 = x_60239 & x_60240;
assign x_60242 = x_28954 & x_28955;
assign x_60243 = x_28956 & x_28957;
assign x_60244 = x_60242 & x_60243;
assign x_60245 = x_60241 & x_60244;
assign x_60246 = x_60238 & x_60245;
assign x_60247 = x_28958 & x_28959;
assign x_60248 = x_28960 & x_28961;
assign x_60249 = x_60247 & x_60248;
assign x_60250 = x_28962 & x_28963;
assign x_60251 = x_28964 & x_28965;
assign x_60252 = x_60250 & x_60251;
assign x_60253 = x_60249 & x_60252;
assign x_60254 = x_28966 & x_28967;
assign x_60255 = x_28968 & x_28969;
assign x_60256 = x_60254 & x_60255;
assign x_60257 = x_28970 & x_28971;
assign x_60258 = x_28972 & x_28973;
assign x_60259 = x_60257 & x_60258;
assign x_60260 = x_60256 & x_60259;
assign x_60261 = x_60253 & x_60260;
assign x_60262 = x_60246 & x_60261;
assign x_60263 = x_60232 & x_60262;
assign x_60264 = x_60203 & x_60263;
assign x_60265 = x_28975 & x_28976;
assign x_60266 = x_28974 & x_60265;
assign x_60267 = x_28977 & x_28978;
assign x_60268 = x_28979 & x_28980;
assign x_60269 = x_60267 & x_60268;
assign x_60270 = x_60266 & x_60269;
assign x_60271 = x_28981 & x_28982;
assign x_60272 = x_28983 & x_28984;
assign x_60273 = x_60271 & x_60272;
assign x_60274 = x_28985 & x_28986;
assign x_60275 = x_28987 & x_28988;
assign x_60276 = x_60274 & x_60275;
assign x_60277 = x_60273 & x_60276;
assign x_60278 = x_60270 & x_60277;
assign x_60279 = x_28990 & x_28991;
assign x_60280 = x_28989 & x_60279;
assign x_60281 = x_28992 & x_28993;
assign x_60282 = x_28994 & x_28995;
assign x_60283 = x_60281 & x_60282;
assign x_60284 = x_60280 & x_60283;
assign x_60285 = x_28996 & x_28997;
assign x_60286 = x_28998 & x_28999;
assign x_60287 = x_60285 & x_60286;
assign x_60288 = x_29000 & x_29001;
assign x_60289 = x_29002 & x_29003;
assign x_60290 = x_60288 & x_60289;
assign x_60291 = x_60287 & x_60290;
assign x_60292 = x_60284 & x_60291;
assign x_60293 = x_60278 & x_60292;
assign x_60294 = x_29005 & x_29006;
assign x_60295 = x_29004 & x_60294;
assign x_60296 = x_29007 & x_29008;
assign x_60297 = x_29009 & x_29010;
assign x_60298 = x_60296 & x_60297;
assign x_60299 = x_60295 & x_60298;
assign x_60300 = x_29011 & x_29012;
assign x_60301 = x_29013 & x_29014;
assign x_60302 = x_60300 & x_60301;
assign x_60303 = x_29015 & x_29016;
assign x_60304 = x_29017 & x_29018;
assign x_60305 = x_60303 & x_60304;
assign x_60306 = x_60302 & x_60305;
assign x_60307 = x_60299 & x_60306;
assign x_60308 = x_29019 & x_29020;
assign x_60309 = x_29021 & x_29022;
assign x_60310 = x_60308 & x_60309;
assign x_60311 = x_29023 & x_29024;
assign x_60312 = x_29025 & x_29026;
assign x_60313 = x_60311 & x_60312;
assign x_60314 = x_60310 & x_60313;
assign x_60315 = x_29027 & x_29028;
assign x_60316 = x_29029 & x_29030;
assign x_60317 = x_60315 & x_60316;
assign x_60318 = x_29031 & x_29032;
assign x_60319 = x_29033 & x_29034;
assign x_60320 = x_60318 & x_60319;
assign x_60321 = x_60317 & x_60320;
assign x_60322 = x_60314 & x_60321;
assign x_60323 = x_60307 & x_60322;
assign x_60324 = x_60293 & x_60323;
assign x_60325 = x_29036 & x_29037;
assign x_60326 = x_29035 & x_60325;
assign x_60327 = x_29038 & x_29039;
assign x_60328 = x_29040 & x_29041;
assign x_60329 = x_60327 & x_60328;
assign x_60330 = x_60326 & x_60329;
assign x_60331 = x_29042 & x_29043;
assign x_60332 = x_29044 & x_29045;
assign x_60333 = x_60331 & x_60332;
assign x_60334 = x_29046 & x_29047;
assign x_60335 = x_29048 & x_29049;
assign x_60336 = x_60334 & x_60335;
assign x_60337 = x_60333 & x_60336;
assign x_60338 = x_60330 & x_60337;
assign x_60339 = x_29051 & x_29052;
assign x_60340 = x_29050 & x_60339;
assign x_60341 = x_29053 & x_29054;
assign x_60342 = x_29055 & x_29056;
assign x_60343 = x_60341 & x_60342;
assign x_60344 = x_60340 & x_60343;
assign x_60345 = x_29057 & x_29058;
assign x_60346 = x_29059 & x_29060;
assign x_60347 = x_60345 & x_60346;
assign x_60348 = x_29061 & x_29062;
assign x_60349 = x_29063 & x_29064;
assign x_60350 = x_60348 & x_60349;
assign x_60351 = x_60347 & x_60350;
assign x_60352 = x_60344 & x_60351;
assign x_60353 = x_60338 & x_60352;
assign x_60354 = x_29066 & x_29067;
assign x_60355 = x_29065 & x_60354;
assign x_60356 = x_29068 & x_29069;
assign x_60357 = x_29070 & x_29071;
assign x_60358 = x_60356 & x_60357;
assign x_60359 = x_60355 & x_60358;
assign x_60360 = x_29072 & x_29073;
assign x_60361 = x_29074 & x_29075;
assign x_60362 = x_60360 & x_60361;
assign x_60363 = x_29076 & x_29077;
assign x_60364 = x_29078 & x_29079;
assign x_60365 = x_60363 & x_60364;
assign x_60366 = x_60362 & x_60365;
assign x_60367 = x_60359 & x_60366;
assign x_60368 = x_29080 & x_29081;
assign x_60369 = x_29082 & x_29083;
assign x_60370 = x_60368 & x_60369;
assign x_60371 = x_29084 & x_29085;
assign x_60372 = x_29086 & x_29087;
assign x_60373 = x_60371 & x_60372;
assign x_60374 = x_60370 & x_60373;
assign x_60375 = x_29088 & x_29089;
assign x_60376 = x_29090 & x_29091;
assign x_60377 = x_60375 & x_60376;
assign x_60378 = x_29092 & x_29093;
assign x_60379 = x_29094 & x_29095;
assign x_60380 = x_60378 & x_60379;
assign x_60381 = x_60377 & x_60380;
assign x_60382 = x_60374 & x_60381;
assign x_60383 = x_60367 & x_60382;
assign x_60384 = x_60353 & x_60383;
assign x_60385 = x_60324 & x_60384;
assign x_60386 = x_60264 & x_60385;
assign x_60387 = x_29097 & x_29098;
assign x_60388 = x_29096 & x_60387;
assign x_60389 = x_29099 & x_29100;
assign x_60390 = x_29101 & x_29102;
assign x_60391 = x_60389 & x_60390;
assign x_60392 = x_60388 & x_60391;
assign x_60393 = x_29103 & x_29104;
assign x_60394 = x_29105 & x_29106;
assign x_60395 = x_60393 & x_60394;
assign x_60396 = x_29107 & x_29108;
assign x_60397 = x_29109 & x_29110;
assign x_60398 = x_60396 & x_60397;
assign x_60399 = x_60395 & x_60398;
assign x_60400 = x_60392 & x_60399;
assign x_60401 = x_29112 & x_29113;
assign x_60402 = x_29111 & x_60401;
assign x_60403 = x_29114 & x_29115;
assign x_60404 = x_29116 & x_29117;
assign x_60405 = x_60403 & x_60404;
assign x_60406 = x_60402 & x_60405;
assign x_60407 = x_29118 & x_29119;
assign x_60408 = x_29120 & x_29121;
assign x_60409 = x_60407 & x_60408;
assign x_60410 = x_29122 & x_29123;
assign x_60411 = x_29124 & x_29125;
assign x_60412 = x_60410 & x_60411;
assign x_60413 = x_60409 & x_60412;
assign x_60414 = x_60406 & x_60413;
assign x_60415 = x_60400 & x_60414;
assign x_60416 = x_29127 & x_29128;
assign x_60417 = x_29126 & x_60416;
assign x_60418 = x_29129 & x_29130;
assign x_60419 = x_29131 & x_29132;
assign x_60420 = x_60418 & x_60419;
assign x_60421 = x_60417 & x_60420;
assign x_60422 = x_29133 & x_29134;
assign x_60423 = x_29135 & x_29136;
assign x_60424 = x_60422 & x_60423;
assign x_60425 = x_29137 & x_29138;
assign x_60426 = x_29139 & x_29140;
assign x_60427 = x_60425 & x_60426;
assign x_60428 = x_60424 & x_60427;
assign x_60429 = x_60421 & x_60428;
assign x_60430 = x_29141 & x_29142;
assign x_60431 = x_29143 & x_29144;
assign x_60432 = x_60430 & x_60431;
assign x_60433 = x_29145 & x_29146;
assign x_60434 = x_29147 & x_29148;
assign x_60435 = x_60433 & x_60434;
assign x_60436 = x_60432 & x_60435;
assign x_60437 = x_29149 & x_29150;
assign x_60438 = x_29151 & x_29152;
assign x_60439 = x_60437 & x_60438;
assign x_60440 = x_29153 & x_29154;
assign x_60441 = x_29155 & x_29156;
assign x_60442 = x_60440 & x_60441;
assign x_60443 = x_60439 & x_60442;
assign x_60444 = x_60436 & x_60443;
assign x_60445 = x_60429 & x_60444;
assign x_60446 = x_60415 & x_60445;
assign x_60447 = x_29158 & x_29159;
assign x_60448 = x_29157 & x_60447;
assign x_60449 = x_29160 & x_29161;
assign x_60450 = x_29162 & x_29163;
assign x_60451 = x_60449 & x_60450;
assign x_60452 = x_60448 & x_60451;
assign x_60453 = x_29164 & x_29165;
assign x_60454 = x_29166 & x_29167;
assign x_60455 = x_60453 & x_60454;
assign x_60456 = x_29168 & x_29169;
assign x_60457 = x_29170 & x_29171;
assign x_60458 = x_60456 & x_60457;
assign x_60459 = x_60455 & x_60458;
assign x_60460 = x_60452 & x_60459;
assign x_60461 = x_29173 & x_29174;
assign x_60462 = x_29172 & x_60461;
assign x_60463 = x_29175 & x_29176;
assign x_60464 = x_29177 & x_29178;
assign x_60465 = x_60463 & x_60464;
assign x_60466 = x_60462 & x_60465;
assign x_60467 = x_29179 & x_29180;
assign x_60468 = x_29181 & x_29182;
assign x_60469 = x_60467 & x_60468;
assign x_60470 = x_29183 & x_29184;
assign x_60471 = x_29185 & x_29186;
assign x_60472 = x_60470 & x_60471;
assign x_60473 = x_60469 & x_60472;
assign x_60474 = x_60466 & x_60473;
assign x_60475 = x_60460 & x_60474;
assign x_60476 = x_29188 & x_29189;
assign x_60477 = x_29187 & x_60476;
assign x_60478 = x_29190 & x_29191;
assign x_60479 = x_29192 & x_29193;
assign x_60480 = x_60478 & x_60479;
assign x_60481 = x_60477 & x_60480;
assign x_60482 = x_29194 & x_29195;
assign x_60483 = x_29196 & x_29197;
assign x_60484 = x_60482 & x_60483;
assign x_60485 = x_29198 & x_29199;
assign x_60486 = x_29200 & x_29201;
assign x_60487 = x_60485 & x_60486;
assign x_60488 = x_60484 & x_60487;
assign x_60489 = x_60481 & x_60488;
assign x_60490 = x_29202 & x_29203;
assign x_60491 = x_29204 & x_29205;
assign x_60492 = x_60490 & x_60491;
assign x_60493 = x_29206 & x_29207;
assign x_60494 = x_29208 & x_29209;
assign x_60495 = x_60493 & x_60494;
assign x_60496 = x_60492 & x_60495;
assign x_60497 = x_29210 & x_29211;
assign x_60498 = x_29212 & x_29213;
assign x_60499 = x_60497 & x_60498;
assign x_60500 = x_29214 & x_29215;
assign x_60501 = x_29216 & x_29217;
assign x_60502 = x_60500 & x_60501;
assign x_60503 = x_60499 & x_60502;
assign x_60504 = x_60496 & x_60503;
assign x_60505 = x_60489 & x_60504;
assign x_60506 = x_60475 & x_60505;
assign x_60507 = x_60446 & x_60506;
assign x_60508 = x_29219 & x_29220;
assign x_60509 = x_29218 & x_60508;
assign x_60510 = x_29221 & x_29222;
assign x_60511 = x_29223 & x_29224;
assign x_60512 = x_60510 & x_60511;
assign x_60513 = x_60509 & x_60512;
assign x_60514 = x_29225 & x_29226;
assign x_60515 = x_29227 & x_29228;
assign x_60516 = x_60514 & x_60515;
assign x_60517 = x_29229 & x_29230;
assign x_60518 = x_29231 & x_29232;
assign x_60519 = x_60517 & x_60518;
assign x_60520 = x_60516 & x_60519;
assign x_60521 = x_60513 & x_60520;
assign x_60522 = x_29234 & x_29235;
assign x_60523 = x_29233 & x_60522;
assign x_60524 = x_29236 & x_29237;
assign x_60525 = x_29238 & x_29239;
assign x_60526 = x_60524 & x_60525;
assign x_60527 = x_60523 & x_60526;
assign x_60528 = x_29240 & x_29241;
assign x_60529 = x_29242 & x_29243;
assign x_60530 = x_60528 & x_60529;
assign x_60531 = x_29244 & x_29245;
assign x_60532 = x_29246 & x_29247;
assign x_60533 = x_60531 & x_60532;
assign x_60534 = x_60530 & x_60533;
assign x_60535 = x_60527 & x_60534;
assign x_60536 = x_60521 & x_60535;
assign x_60537 = x_29249 & x_29250;
assign x_60538 = x_29248 & x_60537;
assign x_60539 = x_29251 & x_29252;
assign x_60540 = x_29253 & x_29254;
assign x_60541 = x_60539 & x_60540;
assign x_60542 = x_60538 & x_60541;
assign x_60543 = x_29255 & x_29256;
assign x_60544 = x_29257 & x_29258;
assign x_60545 = x_60543 & x_60544;
assign x_60546 = x_29259 & x_29260;
assign x_60547 = x_29261 & x_29262;
assign x_60548 = x_60546 & x_60547;
assign x_60549 = x_60545 & x_60548;
assign x_60550 = x_60542 & x_60549;
assign x_60551 = x_29263 & x_29264;
assign x_60552 = x_29265 & x_29266;
assign x_60553 = x_60551 & x_60552;
assign x_60554 = x_29267 & x_29268;
assign x_60555 = x_29269 & x_29270;
assign x_60556 = x_60554 & x_60555;
assign x_60557 = x_60553 & x_60556;
assign x_60558 = x_29271 & x_29272;
assign x_60559 = x_29273 & x_29274;
assign x_60560 = x_60558 & x_60559;
assign x_60561 = x_29275 & x_29276;
assign x_60562 = x_29277 & x_29278;
assign x_60563 = x_60561 & x_60562;
assign x_60564 = x_60560 & x_60563;
assign x_60565 = x_60557 & x_60564;
assign x_60566 = x_60550 & x_60565;
assign x_60567 = x_60536 & x_60566;
assign x_60568 = x_29280 & x_29281;
assign x_60569 = x_29279 & x_60568;
assign x_60570 = x_29282 & x_29283;
assign x_60571 = x_29284 & x_29285;
assign x_60572 = x_60570 & x_60571;
assign x_60573 = x_60569 & x_60572;
assign x_60574 = x_29286 & x_29287;
assign x_60575 = x_29288 & x_29289;
assign x_60576 = x_60574 & x_60575;
assign x_60577 = x_29290 & x_29291;
assign x_60578 = x_29292 & x_29293;
assign x_60579 = x_60577 & x_60578;
assign x_60580 = x_60576 & x_60579;
assign x_60581 = x_60573 & x_60580;
assign x_60582 = x_29294 & x_29295;
assign x_60583 = x_29296 & x_29297;
assign x_60584 = x_60582 & x_60583;
assign x_60585 = x_29298 & x_29299;
assign x_60586 = x_29300 & x_29301;
assign x_60587 = x_60585 & x_60586;
assign x_60588 = x_60584 & x_60587;
assign x_60589 = x_29302 & x_29303;
assign x_60590 = x_29304 & x_29305;
assign x_60591 = x_60589 & x_60590;
assign x_60592 = x_29306 & x_29307;
assign x_60593 = x_29308 & x_29309;
assign x_60594 = x_60592 & x_60593;
assign x_60595 = x_60591 & x_60594;
assign x_60596 = x_60588 & x_60595;
assign x_60597 = x_60581 & x_60596;
assign x_60598 = x_29311 & x_29312;
assign x_60599 = x_29310 & x_60598;
assign x_60600 = x_29313 & x_29314;
assign x_60601 = x_29315 & x_29316;
assign x_60602 = x_60600 & x_60601;
assign x_60603 = x_60599 & x_60602;
assign x_60604 = x_29317 & x_29318;
assign x_60605 = x_29319 & x_29320;
assign x_60606 = x_60604 & x_60605;
assign x_60607 = x_29321 & x_29322;
assign x_60608 = x_29323 & x_29324;
assign x_60609 = x_60607 & x_60608;
assign x_60610 = x_60606 & x_60609;
assign x_60611 = x_60603 & x_60610;
assign x_60612 = x_29325 & x_29326;
assign x_60613 = x_29327 & x_29328;
assign x_60614 = x_60612 & x_60613;
assign x_60615 = x_29329 & x_29330;
assign x_60616 = x_29331 & x_29332;
assign x_60617 = x_60615 & x_60616;
assign x_60618 = x_60614 & x_60617;
assign x_60619 = x_29333 & x_29334;
assign x_60620 = x_29335 & x_29336;
assign x_60621 = x_60619 & x_60620;
assign x_60622 = x_29337 & x_29338;
assign x_60623 = x_29339 & x_29340;
assign x_60624 = x_60622 & x_60623;
assign x_60625 = x_60621 & x_60624;
assign x_60626 = x_60618 & x_60625;
assign x_60627 = x_60611 & x_60626;
assign x_60628 = x_60597 & x_60627;
assign x_60629 = x_60567 & x_60628;
assign x_60630 = x_60507 & x_60629;
assign x_60631 = x_60386 & x_60630;
assign x_60632 = x_60143 & x_60631;
assign x_60633 = x_59655 & x_60632;
assign x_60634 = x_29342 & x_29343;
assign x_60635 = x_29341 & x_60634;
assign x_60636 = x_29344 & x_29345;
assign x_60637 = x_29346 & x_29347;
assign x_60638 = x_60636 & x_60637;
assign x_60639 = x_60635 & x_60638;
assign x_60640 = x_29348 & x_29349;
assign x_60641 = x_29350 & x_29351;
assign x_60642 = x_60640 & x_60641;
assign x_60643 = x_29352 & x_29353;
assign x_60644 = x_29354 & x_29355;
assign x_60645 = x_60643 & x_60644;
assign x_60646 = x_60642 & x_60645;
assign x_60647 = x_60639 & x_60646;
assign x_60648 = x_29357 & x_29358;
assign x_60649 = x_29356 & x_60648;
assign x_60650 = x_29359 & x_29360;
assign x_60651 = x_29361 & x_29362;
assign x_60652 = x_60650 & x_60651;
assign x_60653 = x_60649 & x_60652;
assign x_60654 = x_29363 & x_29364;
assign x_60655 = x_29365 & x_29366;
assign x_60656 = x_60654 & x_60655;
assign x_60657 = x_29367 & x_29368;
assign x_60658 = x_29369 & x_29370;
assign x_60659 = x_60657 & x_60658;
assign x_60660 = x_60656 & x_60659;
assign x_60661 = x_60653 & x_60660;
assign x_60662 = x_60647 & x_60661;
assign x_60663 = x_29372 & x_29373;
assign x_60664 = x_29371 & x_60663;
assign x_60665 = x_29374 & x_29375;
assign x_60666 = x_29376 & x_29377;
assign x_60667 = x_60665 & x_60666;
assign x_60668 = x_60664 & x_60667;
assign x_60669 = x_29378 & x_29379;
assign x_60670 = x_29380 & x_29381;
assign x_60671 = x_60669 & x_60670;
assign x_60672 = x_29382 & x_29383;
assign x_60673 = x_29384 & x_29385;
assign x_60674 = x_60672 & x_60673;
assign x_60675 = x_60671 & x_60674;
assign x_60676 = x_60668 & x_60675;
assign x_60677 = x_29386 & x_29387;
assign x_60678 = x_29388 & x_29389;
assign x_60679 = x_60677 & x_60678;
assign x_60680 = x_29390 & x_29391;
assign x_60681 = x_29392 & x_29393;
assign x_60682 = x_60680 & x_60681;
assign x_60683 = x_60679 & x_60682;
assign x_60684 = x_29394 & x_29395;
assign x_60685 = x_29396 & x_29397;
assign x_60686 = x_60684 & x_60685;
assign x_60687 = x_29398 & x_29399;
assign x_60688 = x_29400 & x_29401;
assign x_60689 = x_60687 & x_60688;
assign x_60690 = x_60686 & x_60689;
assign x_60691 = x_60683 & x_60690;
assign x_60692 = x_60676 & x_60691;
assign x_60693 = x_60662 & x_60692;
assign x_60694 = x_29403 & x_29404;
assign x_60695 = x_29402 & x_60694;
assign x_60696 = x_29405 & x_29406;
assign x_60697 = x_29407 & x_29408;
assign x_60698 = x_60696 & x_60697;
assign x_60699 = x_60695 & x_60698;
assign x_60700 = x_29409 & x_29410;
assign x_60701 = x_29411 & x_29412;
assign x_60702 = x_60700 & x_60701;
assign x_60703 = x_29413 & x_29414;
assign x_60704 = x_29415 & x_29416;
assign x_60705 = x_60703 & x_60704;
assign x_60706 = x_60702 & x_60705;
assign x_60707 = x_60699 & x_60706;
assign x_60708 = x_29418 & x_29419;
assign x_60709 = x_29417 & x_60708;
assign x_60710 = x_29420 & x_29421;
assign x_60711 = x_29422 & x_29423;
assign x_60712 = x_60710 & x_60711;
assign x_60713 = x_60709 & x_60712;
assign x_60714 = x_29424 & x_29425;
assign x_60715 = x_29426 & x_29427;
assign x_60716 = x_60714 & x_60715;
assign x_60717 = x_29428 & x_29429;
assign x_60718 = x_29430 & x_29431;
assign x_60719 = x_60717 & x_60718;
assign x_60720 = x_60716 & x_60719;
assign x_60721 = x_60713 & x_60720;
assign x_60722 = x_60707 & x_60721;
assign x_60723 = x_29433 & x_29434;
assign x_60724 = x_29432 & x_60723;
assign x_60725 = x_29435 & x_29436;
assign x_60726 = x_29437 & x_29438;
assign x_60727 = x_60725 & x_60726;
assign x_60728 = x_60724 & x_60727;
assign x_60729 = x_29439 & x_29440;
assign x_60730 = x_29441 & x_29442;
assign x_60731 = x_60729 & x_60730;
assign x_60732 = x_29443 & x_29444;
assign x_60733 = x_29445 & x_29446;
assign x_60734 = x_60732 & x_60733;
assign x_60735 = x_60731 & x_60734;
assign x_60736 = x_60728 & x_60735;
assign x_60737 = x_29447 & x_29448;
assign x_60738 = x_29449 & x_29450;
assign x_60739 = x_60737 & x_60738;
assign x_60740 = x_29451 & x_29452;
assign x_60741 = x_29453 & x_29454;
assign x_60742 = x_60740 & x_60741;
assign x_60743 = x_60739 & x_60742;
assign x_60744 = x_29455 & x_29456;
assign x_60745 = x_29457 & x_29458;
assign x_60746 = x_60744 & x_60745;
assign x_60747 = x_29459 & x_29460;
assign x_60748 = x_29461 & x_29462;
assign x_60749 = x_60747 & x_60748;
assign x_60750 = x_60746 & x_60749;
assign x_60751 = x_60743 & x_60750;
assign x_60752 = x_60736 & x_60751;
assign x_60753 = x_60722 & x_60752;
assign x_60754 = x_60693 & x_60753;
assign x_60755 = x_29464 & x_29465;
assign x_60756 = x_29463 & x_60755;
assign x_60757 = x_29466 & x_29467;
assign x_60758 = x_29468 & x_29469;
assign x_60759 = x_60757 & x_60758;
assign x_60760 = x_60756 & x_60759;
assign x_60761 = x_29470 & x_29471;
assign x_60762 = x_29472 & x_29473;
assign x_60763 = x_60761 & x_60762;
assign x_60764 = x_29474 & x_29475;
assign x_60765 = x_29476 & x_29477;
assign x_60766 = x_60764 & x_60765;
assign x_60767 = x_60763 & x_60766;
assign x_60768 = x_60760 & x_60767;
assign x_60769 = x_29479 & x_29480;
assign x_60770 = x_29478 & x_60769;
assign x_60771 = x_29481 & x_29482;
assign x_60772 = x_29483 & x_29484;
assign x_60773 = x_60771 & x_60772;
assign x_60774 = x_60770 & x_60773;
assign x_60775 = x_29485 & x_29486;
assign x_60776 = x_29487 & x_29488;
assign x_60777 = x_60775 & x_60776;
assign x_60778 = x_29489 & x_29490;
assign x_60779 = x_29491 & x_29492;
assign x_60780 = x_60778 & x_60779;
assign x_60781 = x_60777 & x_60780;
assign x_60782 = x_60774 & x_60781;
assign x_60783 = x_60768 & x_60782;
assign x_60784 = x_29494 & x_29495;
assign x_60785 = x_29493 & x_60784;
assign x_60786 = x_29496 & x_29497;
assign x_60787 = x_29498 & x_29499;
assign x_60788 = x_60786 & x_60787;
assign x_60789 = x_60785 & x_60788;
assign x_60790 = x_29500 & x_29501;
assign x_60791 = x_29502 & x_29503;
assign x_60792 = x_60790 & x_60791;
assign x_60793 = x_29504 & x_29505;
assign x_60794 = x_29506 & x_29507;
assign x_60795 = x_60793 & x_60794;
assign x_60796 = x_60792 & x_60795;
assign x_60797 = x_60789 & x_60796;
assign x_60798 = x_29508 & x_29509;
assign x_60799 = x_29510 & x_29511;
assign x_60800 = x_60798 & x_60799;
assign x_60801 = x_29512 & x_29513;
assign x_60802 = x_29514 & x_29515;
assign x_60803 = x_60801 & x_60802;
assign x_60804 = x_60800 & x_60803;
assign x_60805 = x_29516 & x_29517;
assign x_60806 = x_29518 & x_29519;
assign x_60807 = x_60805 & x_60806;
assign x_60808 = x_29520 & x_29521;
assign x_60809 = x_29522 & x_29523;
assign x_60810 = x_60808 & x_60809;
assign x_60811 = x_60807 & x_60810;
assign x_60812 = x_60804 & x_60811;
assign x_60813 = x_60797 & x_60812;
assign x_60814 = x_60783 & x_60813;
assign x_60815 = x_29525 & x_29526;
assign x_60816 = x_29524 & x_60815;
assign x_60817 = x_29527 & x_29528;
assign x_60818 = x_29529 & x_29530;
assign x_60819 = x_60817 & x_60818;
assign x_60820 = x_60816 & x_60819;
assign x_60821 = x_29531 & x_29532;
assign x_60822 = x_29533 & x_29534;
assign x_60823 = x_60821 & x_60822;
assign x_60824 = x_29535 & x_29536;
assign x_60825 = x_29537 & x_29538;
assign x_60826 = x_60824 & x_60825;
assign x_60827 = x_60823 & x_60826;
assign x_60828 = x_60820 & x_60827;
assign x_60829 = x_29540 & x_29541;
assign x_60830 = x_29539 & x_60829;
assign x_60831 = x_29542 & x_29543;
assign x_60832 = x_29544 & x_29545;
assign x_60833 = x_60831 & x_60832;
assign x_60834 = x_60830 & x_60833;
assign x_60835 = x_29546 & x_29547;
assign x_60836 = x_29548 & x_29549;
assign x_60837 = x_60835 & x_60836;
assign x_60838 = x_29550 & x_29551;
assign x_60839 = x_29552 & x_29553;
assign x_60840 = x_60838 & x_60839;
assign x_60841 = x_60837 & x_60840;
assign x_60842 = x_60834 & x_60841;
assign x_60843 = x_60828 & x_60842;
assign x_60844 = x_29555 & x_29556;
assign x_60845 = x_29554 & x_60844;
assign x_60846 = x_29557 & x_29558;
assign x_60847 = x_29559 & x_29560;
assign x_60848 = x_60846 & x_60847;
assign x_60849 = x_60845 & x_60848;
assign x_60850 = x_29561 & x_29562;
assign x_60851 = x_29563 & x_29564;
assign x_60852 = x_60850 & x_60851;
assign x_60853 = x_29565 & x_29566;
assign x_60854 = x_29567 & x_29568;
assign x_60855 = x_60853 & x_60854;
assign x_60856 = x_60852 & x_60855;
assign x_60857 = x_60849 & x_60856;
assign x_60858 = x_29569 & x_29570;
assign x_60859 = x_29571 & x_29572;
assign x_60860 = x_60858 & x_60859;
assign x_60861 = x_29573 & x_29574;
assign x_60862 = x_29575 & x_29576;
assign x_60863 = x_60861 & x_60862;
assign x_60864 = x_60860 & x_60863;
assign x_60865 = x_29577 & x_29578;
assign x_60866 = x_29579 & x_29580;
assign x_60867 = x_60865 & x_60866;
assign x_60868 = x_29581 & x_29582;
assign x_60869 = x_29583 & x_29584;
assign x_60870 = x_60868 & x_60869;
assign x_60871 = x_60867 & x_60870;
assign x_60872 = x_60864 & x_60871;
assign x_60873 = x_60857 & x_60872;
assign x_60874 = x_60843 & x_60873;
assign x_60875 = x_60814 & x_60874;
assign x_60876 = x_60754 & x_60875;
assign x_60877 = x_29586 & x_29587;
assign x_60878 = x_29585 & x_60877;
assign x_60879 = x_29588 & x_29589;
assign x_60880 = x_29590 & x_29591;
assign x_60881 = x_60879 & x_60880;
assign x_60882 = x_60878 & x_60881;
assign x_60883 = x_29592 & x_29593;
assign x_60884 = x_29594 & x_29595;
assign x_60885 = x_60883 & x_60884;
assign x_60886 = x_29596 & x_29597;
assign x_60887 = x_29598 & x_29599;
assign x_60888 = x_60886 & x_60887;
assign x_60889 = x_60885 & x_60888;
assign x_60890 = x_60882 & x_60889;
assign x_60891 = x_29601 & x_29602;
assign x_60892 = x_29600 & x_60891;
assign x_60893 = x_29603 & x_29604;
assign x_60894 = x_29605 & x_29606;
assign x_60895 = x_60893 & x_60894;
assign x_60896 = x_60892 & x_60895;
assign x_60897 = x_29607 & x_29608;
assign x_60898 = x_29609 & x_29610;
assign x_60899 = x_60897 & x_60898;
assign x_60900 = x_29611 & x_29612;
assign x_60901 = x_29613 & x_29614;
assign x_60902 = x_60900 & x_60901;
assign x_60903 = x_60899 & x_60902;
assign x_60904 = x_60896 & x_60903;
assign x_60905 = x_60890 & x_60904;
assign x_60906 = x_29616 & x_29617;
assign x_60907 = x_29615 & x_60906;
assign x_60908 = x_29618 & x_29619;
assign x_60909 = x_29620 & x_29621;
assign x_60910 = x_60908 & x_60909;
assign x_60911 = x_60907 & x_60910;
assign x_60912 = x_29622 & x_29623;
assign x_60913 = x_29624 & x_29625;
assign x_60914 = x_60912 & x_60913;
assign x_60915 = x_29626 & x_29627;
assign x_60916 = x_29628 & x_29629;
assign x_60917 = x_60915 & x_60916;
assign x_60918 = x_60914 & x_60917;
assign x_60919 = x_60911 & x_60918;
assign x_60920 = x_29630 & x_29631;
assign x_60921 = x_29632 & x_29633;
assign x_60922 = x_60920 & x_60921;
assign x_60923 = x_29634 & x_29635;
assign x_60924 = x_29636 & x_29637;
assign x_60925 = x_60923 & x_60924;
assign x_60926 = x_60922 & x_60925;
assign x_60927 = x_29638 & x_29639;
assign x_60928 = x_29640 & x_29641;
assign x_60929 = x_60927 & x_60928;
assign x_60930 = x_29642 & x_29643;
assign x_60931 = x_29644 & x_29645;
assign x_60932 = x_60930 & x_60931;
assign x_60933 = x_60929 & x_60932;
assign x_60934 = x_60926 & x_60933;
assign x_60935 = x_60919 & x_60934;
assign x_60936 = x_60905 & x_60935;
assign x_60937 = x_29647 & x_29648;
assign x_60938 = x_29646 & x_60937;
assign x_60939 = x_29649 & x_29650;
assign x_60940 = x_29651 & x_29652;
assign x_60941 = x_60939 & x_60940;
assign x_60942 = x_60938 & x_60941;
assign x_60943 = x_29653 & x_29654;
assign x_60944 = x_29655 & x_29656;
assign x_60945 = x_60943 & x_60944;
assign x_60946 = x_29657 & x_29658;
assign x_60947 = x_29659 & x_29660;
assign x_60948 = x_60946 & x_60947;
assign x_60949 = x_60945 & x_60948;
assign x_60950 = x_60942 & x_60949;
assign x_60951 = x_29662 & x_29663;
assign x_60952 = x_29661 & x_60951;
assign x_60953 = x_29664 & x_29665;
assign x_60954 = x_29666 & x_29667;
assign x_60955 = x_60953 & x_60954;
assign x_60956 = x_60952 & x_60955;
assign x_60957 = x_29668 & x_29669;
assign x_60958 = x_29670 & x_29671;
assign x_60959 = x_60957 & x_60958;
assign x_60960 = x_29672 & x_29673;
assign x_60961 = x_29674 & x_29675;
assign x_60962 = x_60960 & x_60961;
assign x_60963 = x_60959 & x_60962;
assign x_60964 = x_60956 & x_60963;
assign x_60965 = x_60950 & x_60964;
assign x_60966 = x_29677 & x_29678;
assign x_60967 = x_29676 & x_60966;
assign x_60968 = x_29679 & x_29680;
assign x_60969 = x_29681 & x_29682;
assign x_60970 = x_60968 & x_60969;
assign x_60971 = x_60967 & x_60970;
assign x_60972 = x_29683 & x_29684;
assign x_60973 = x_29685 & x_29686;
assign x_60974 = x_60972 & x_60973;
assign x_60975 = x_29687 & x_29688;
assign x_60976 = x_29689 & x_29690;
assign x_60977 = x_60975 & x_60976;
assign x_60978 = x_60974 & x_60977;
assign x_60979 = x_60971 & x_60978;
assign x_60980 = x_29691 & x_29692;
assign x_60981 = x_29693 & x_29694;
assign x_60982 = x_60980 & x_60981;
assign x_60983 = x_29695 & x_29696;
assign x_60984 = x_29697 & x_29698;
assign x_60985 = x_60983 & x_60984;
assign x_60986 = x_60982 & x_60985;
assign x_60987 = x_29699 & x_29700;
assign x_60988 = x_29701 & x_29702;
assign x_60989 = x_60987 & x_60988;
assign x_60990 = x_29703 & x_29704;
assign x_60991 = x_29705 & x_29706;
assign x_60992 = x_60990 & x_60991;
assign x_60993 = x_60989 & x_60992;
assign x_60994 = x_60986 & x_60993;
assign x_60995 = x_60979 & x_60994;
assign x_60996 = x_60965 & x_60995;
assign x_60997 = x_60936 & x_60996;
assign x_60998 = x_29708 & x_29709;
assign x_60999 = x_29707 & x_60998;
assign x_61000 = x_29710 & x_29711;
assign x_61001 = x_29712 & x_29713;
assign x_61002 = x_61000 & x_61001;
assign x_61003 = x_60999 & x_61002;
assign x_61004 = x_29714 & x_29715;
assign x_61005 = x_29716 & x_29717;
assign x_61006 = x_61004 & x_61005;
assign x_61007 = x_29718 & x_29719;
assign x_61008 = x_29720 & x_29721;
assign x_61009 = x_61007 & x_61008;
assign x_61010 = x_61006 & x_61009;
assign x_61011 = x_61003 & x_61010;
assign x_61012 = x_29723 & x_29724;
assign x_61013 = x_29722 & x_61012;
assign x_61014 = x_29725 & x_29726;
assign x_61015 = x_29727 & x_29728;
assign x_61016 = x_61014 & x_61015;
assign x_61017 = x_61013 & x_61016;
assign x_61018 = x_29729 & x_29730;
assign x_61019 = x_29731 & x_29732;
assign x_61020 = x_61018 & x_61019;
assign x_61021 = x_29733 & x_29734;
assign x_61022 = x_29735 & x_29736;
assign x_61023 = x_61021 & x_61022;
assign x_61024 = x_61020 & x_61023;
assign x_61025 = x_61017 & x_61024;
assign x_61026 = x_61011 & x_61025;
assign x_61027 = x_29738 & x_29739;
assign x_61028 = x_29737 & x_61027;
assign x_61029 = x_29740 & x_29741;
assign x_61030 = x_29742 & x_29743;
assign x_61031 = x_61029 & x_61030;
assign x_61032 = x_61028 & x_61031;
assign x_61033 = x_29744 & x_29745;
assign x_61034 = x_29746 & x_29747;
assign x_61035 = x_61033 & x_61034;
assign x_61036 = x_29748 & x_29749;
assign x_61037 = x_29750 & x_29751;
assign x_61038 = x_61036 & x_61037;
assign x_61039 = x_61035 & x_61038;
assign x_61040 = x_61032 & x_61039;
assign x_61041 = x_29752 & x_29753;
assign x_61042 = x_29754 & x_29755;
assign x_61043 = x_61041 & x_61042;
assign x_61044 = x_29756 & x_29757;
assign x_61045 = x_29758 & x_29759;
assign x_61046 = x_61044 & x_61045;
assign x_61047 = x_61043 & x_61046;
assign x_61048 = x_29760 & x_29761;
assign x_61049 = x_29762 & x_29763;
assign x_61050 = x_61048 & x_61049;
assign x_61051 = x_29764 & x_29765;
assign x_61052 = x_29766 & x_29767;
assign x_61053 = x_61051 & x_61052;
assign x_61054 = x_61050 & x_61053;
assign x_61055 = x_61047 & x_61054;
assign x_61056 = x_61040 & x_61055;
assign x_61057 = x_61026 & x_61056;
assign x_61058 = x_29769 & x_29770;
assign x_61059 = x_29768 & x_61058;
assign x_61060 = x_29771 & x_29772;
assign x_61061 = x_29773 & x_29774;
assign x_61062 = x_61060 & x_61061;
assign x_61063 = x_61059 & x_61062;
assign x_61064 = x_29775 & x_29776;
assign x_61065 = x_29777 & x_29778;
assign x_61066 = x_61064 & x_61065;
assign x_61067 = x_29779 & x_29780;
assign x_61068 = x_29781 & x_29782;
assign x_61069 = x_61067 & x_61068;
assign x_61070 = x_61066 & x_61069;
assign x_61071 = x_61063 & x_61070;
assign x_61072 = x_29783 & x_29784;
assign x_61073 = x_29785 & x_29786;
assign x_61074 = x_61072 & x_61073;
assign x_61075 = x_29787 & x_29788;
assign x_61076 = x_29789 & x_29790;
assign x_61077 = x_61075 & x_61076;
assign x_61078 = x_61074 & x_61077;
assign x_61079 = x_29791 & x_29792;
assign x_61080 = x_29793 & x_29794;
assign x_61081 = x_61079 & x_61080;
assign x_61082 = x_29795 & x_29796;
assign x_61083 = x_29797 & x_29798;
assign x_61084 = x_61082 & x_61083;
assign x_61085 = x_61081 & x_61084;
assign x_61086 = x_61078 & x_61085;
assign x_61087 = x_61071 & x_61086;
assign x_61088 = x_29800 & x_29801;
assign x_61089 = x_29799 & x_61088;
assign x_61090 = x_29802 & x_29803;
assign x_61091 = x_29804 & x_29805;
assign x_61092 = x_61090 & x_61091;
assign x_61093 = x_61089 & x_61092;
assign x_61094 = x_29806 & x_29807;
assign x_61095 = x_29808 & x_29809;
assign x_61096 = x_61094 & x_61095;
assign x_61097 = x_29810 & x_29811;
assign x_61098 = x_29812 & x_29813;
assign x_61099 = x_61097 & x_61098;
assign x_61100 = x_61096 & x_61099;
assign x_61101 = x_61093 & x_61100;
assign x_61102 = x_29814 & x_29815;
assign x_61103 = x_29816 & x_29817;
assign x_61104 = x_61102 & x_61103;
assign x_61105 = x_29818 & x_29819;
assign x_61106 = x_29820 & x_29821;
assign x_61107 = x_61105 & x_61106;
assign x_61108 = x_61104 & x_61107;
assign x_61109 = x_29822 & x_29823;
assign x_61110 = x_29824 & x_29825;
assign x_61111 = x_61109 & x_61110;
assign x_61112 = x_29826 & x_29827;
assign x_61113 = x_29828 & x_29829;
assign x_61114 = x_61112 & x_61113;
assign x_61115 = x_61111 & x_61114;
assign x_61116 = x_61108 & x_61115;
assign x_61117 = x_61101 & x_61116;
assign x_61118 = x_61087 & x_61117;
assign x_61119 = x_61057 & x_61118;
assign x_61120 = x_60997 & x_61119;
assign x_61121 = x_60876 & x_61120;
assign x_61122 = x_29831 & x_29832;
assign x_61123 = x_29830 & x_61122;
assign x_61124 = x_29833 & x_29834;
assign x_61125 = x_29835 & x_29836;
assign x_61126 = x_61124 & x_61125;
assign x_61127 = x_61123 & x_61126;
assign x_61128 = x_29837 & x_29838;
assign x_61129 = x_29839 & x_29840;
assign x_61130 = x_61128 & x_61129;
assign x_61131 = x_29841 & x_29842;
assign x_61132 = x_29843 & x_29844;
assign x_61133 = x_61131 & x_61132;
assign x_61134 = x_61130 & x_61133;
assign x_61135 = x_61127 & x_61134;
assign x_61136 = x_29846 & x_29847;
assign x_61137 = x_29845 & x_61136;
assign x_61138 = x_29848 & x_29849;
assign x_61139 = x_29850 & x_29851;
assign x_61140 = x_61138 & x_61139;
assign x_61141 = x_61137 & x_61140;
assign x_61142 = x_29852 & x_29853;
assign x_61143 = x_29854 & x_29855;
assign x_61144 = x_61142 & x_61143;
assign x_61145 = x_29856 & x_29857;
assign x_61146 = x_29858 & x_29859;
assign x_61147 = x_61145 & x_61146;
assign x_61148 = x_61144 & x_61147;
assign x_61149 = x_61141 & x_61148;
assign x_61150 = x_61135 & x_61149;
assign x_61151 = x_29861 & x_29862;
assign x_61152 = x_29860 & x_61151;
assign x_61153 = x_29863 & x_29864;
assign x_61154 = x_29865 & x_29866;
assign x_61155 = x_61153 & x_61154;
assign x_61156 = x_61152 & x_61155;
assign x_61157 = x_29867 & x_29868;
assign x_61158 = x_29869 & x_29870;
assign x_61159 = x_61157 & x_61158;
assign x_61160 = x_29871 & x_29872;
assign x_61161 = x_29873 & x_29874;
assign x_61162 = x_61160 & x_61161;
assign x_61163 = x_61159 & x_61162;
assign x_61164 = x_61156 & x_61163;
assign x_61165 = x_29875 & x_29876;
assign x_61166 = x_29877 & x_29878;
assign x_61167 = x_61165 & x_61166;
assign x_61168 = x_29879 & x_29880;
assign x_61169 = x_29881 & x_29882;
assign x_61170 = x_61168 & x_61169;
assign x_61171 = x_61167 & x_61170;
assign x_61172 = x_29883 & x_29884;
assign x_61173 = x_29885 & x_29886;
assign x_61174 = x_61172 & x_61173;
assign x_61175 = x_29887 & x_29888;
assign x_61176 = x_29889 & x_29890;
assign x_61177 = x_61175 & x_61176;
assign x_61178 = x_61174 & x_61177;
assign x_61179 = x_61171 & x_61178;
assign x_61180 = x_61164 & x_61179;
assign x_61181 = x_61150 & x_61180;
assign x_61182 = x_29892 & x_29893;
assign x_61183 = x_29891 & x_61182;
assign x_61184 = x_29894 & x_29895;
assign x_61185 = x_29896 & x_29897;
assign x_61186 = x_61184 & x_61185;
assign x_61187 = x_61183 & x_61186;
assign x_61188 = x_29898 & x_29899;
assign x_61189 = x_29900 & x_29901;
assign x_61190 = x_61188 & x_61189;
assign x_61191 = x_29902 & x_29903;
assign x_61192 = x_29904 & x_29905;
assign x_61193 = x_61191 & x_61192;
assign x_61194 = x_61190 & x_61193;
assign x_61195 = x_61187 & x_61194;
assign x_61196 = x_29907 & x_29908;
assign x_61197 = x_29906 & x_61196;
assign x_61198 = x_29909 & x_29910;
assign x_61199 = x_29911 & x_29912;
assign x_61200 = x_61198 & x_61199;
assign x_61201 = x_61197 & x_61200;
assign x_61202 = x_29913 & x_29914;
assign x_61203 = x_29915 & x_29916;
assign x_61204 = x_61202 & x_61203;
assign x_61205 = x_29917 & x_29918;
assign x_61206 = x_29919 & x_29920;
assign x_61207 = x_61205 & x_61206;
assign x_61208 = x_61204 & x_61207;
assign x_61209 = x_61201 & x_61208;
assign x_61210 = x_61195 & x_61209;
assign x_61211 = x_29922 & x_29923;
assign x_61212 = x_29921 & x_61211;
assign x_61213 = x_29924 & x_29925;
assign x_61214 = x_29926 & x_29927;
assign x_61215 = x_61213 & x_61214;
assign x_61216 = x_61212 & x_61215;
assign x_61217 = x_29928 & x_29929;
assign x_61218 = x_29930 & x_29931;
assign x_61219 = x_61217 & x_61218;
assign x_61220 = x_29932 & x_29933;
assign x_61221 = x_29934 & x_29935;
assign x_61222 = x_61220 & x_61221;
assign x_61223 = x_61219 & x_61222;
assign x_61224 = x_61216 & x_61223;
assign x_61225 = x_29936 & x_29937;
assign x_61226 = x_29938 & x_29939;
assign x_61227 = x_61225 & x_61226;
assign x_61228 = x_29940 & x_29941;
assign x_61229 = x_29942 & x_29943;
assign x_61230 = x_61228 & x_61229;
assign x_61231 = x_61227 & x_61230;
assign x_61232 = x_29944 & x_29945;
assign x_61233 = x_29946 & x_29947;
assign x_61234 = x_61232 & x_61233;
assign x_61235 = x_29948 & x_29949;
assign x_61236 = x_29950 & x_29951;
assign x_61237 = x_61235 & x_61236;
assign x_61238 = x_61234 & x_61237;
assign x_61239 = x_61231 & x_61238;
assign x_61240 = x_61224 & x_61239;
assign x_61241 = x_61210 & x_61240;
assign x_61242 = x_61181 & x_61241;
assign x_61243 = x_29953 & x_29954;
assign x_61244 = x_29952 & x_61243;
assign x_61245 = x_29955 & x_29956;
assign x_61246 = x_29957 & x_29958;
assign x_61247 = x_61245 & x_61246;
assign x_61248 = x_61244 & x_61247;
assign x_61249 = x_29959 & x_29960;
assign x_61250 = x_29961 & x_29962;
assign x_61251 = x_61249 & x_61250;
assign x_61252 = x_29963 & x_29964;
assign x_61253 = x_29965 & x_29966;
assign x_61254 = x_61252 & x_61253;
assign x_61255 = x_61251 & x_61254;
assign x_61256 = x_61248 & x_61255;
assign x_61257 = x_29968 & x_29969;
assign x_61258 = x_29967 & x_61257;
assign x_61259 = x_29970 & x_29971;
assign x_61260 = x_29972 & x_29973;
assign x_61261 = x_61259 & x_61260;
assign x_61262 = x_61258 & x_61261;
assign x_61263 = x_29974 & x_29975;
assign x_61264 = x_29976 & x_29977;
assign x_61265 = x_61263 & x_61264;
assign x_61266 = x_29978 & x_29979;
assign x_61267 = x_29980 & x_29981;
assign x_61268 = x_61266 & x_61267;
assign x_61269 = x_61265 & x_61268;
assign x_61270 = x_61262 & x_61269;
assign x_61271 = x_61256 & x_61270;
assign x_61272 = x_29983 & x_29984;
assign x_61273 = x_29982 & x_61272;
assign x_61274 = x_29985 & x_29986;
assign x_61275 = x_29987 & x_29988;
assign x_61276 = x_61274 & x_61275;
assign x_61277 = x_61273 & x_61276;
assign x_61278 = x_29989 & x_29990;
assign x_61279 = x_29991 & x_29992;
assign x_61280 = x_61278 & x_61279;
assign x_61281 = x_29993 & x_29994;
assign x_61282 = x_29995 & x_29996;
assign x_61283 = x_61281 & x_61282;
assign x_61284 = x_61280 & x_61283;
assign x_61285 = x_61277 & x_61284;
assign x_61286 = x_29997 & x_29998;
assign x_61287 = x_29999 & x_30000;
assign x_61288 = x_61286 & x_61287;
assign x_61289 = x_30001 & x_30002;
assign x_61290 = x_30003 & x_30004;
assign x_61291 = x_61289 & x_61290;
assign x_61292 = x_61288 & x_61291;
assign x_61293 = x_30005 & x_30006;
assign x_61294 = x_30007 & x_30008;
assign x_61295 = x_61293 & x_61294;
assign x_61296 = x_30009 & x_30010;
assign x_61297 = x_30011 & x_30012;
assign x_61298 = x_61296 & x_61297;
assign x_61299 = x_61295 & x_61298;
assign x_61300 = x_61292 & x_61299;
assign x_61301 = x_61285 & x_61300;
assign x_61302 = x_61271 & x_61301;
assign x_61303 = x_30014 & x_30015;
assign x_61304 = x_30013 & x_61303;
assign x_61305 = x_30016 & x_30017;
assign x_61306 = x_30018 & x_30019;
assign x_61307 = x_61305 & x_61306;
assign x_61308 = x_61304 & x_61307;
assign x_61309 = x_30020 & x_30021;
assign x_61310 = x_30022 & x_30023;
assign x_61311 = x_61309 & x_61310;
assign x_61312 = x_30024 & x_30025;
assign x_61313 = x_30026 & x_30027;
assign x_61314 = x_61312 & x_61313;
assign x_61315 = x_61311 & x_61314;
assign x_61316 = x_61308 & x_61315;
assign x_61317 = x_30029 & x_30030;
assign x_61318 = x_30028 & x_61317;
assign x_61319 = x_30031 & x_30032;
assign x_61320 = x_30033 & x_30034;
assign x_61321 = x_61319 & x_61320;
assign x_61322 = x_61318 & x_61321;
assign x_61323 = x_30035 & x_30036;
assign x_61324 = x_30037 & x_30038;
assign x_61325 = x_61323 & x_61324;
assign x_61326 = x_30039 & x_30040;
assign x_61327 = x_30041 & x_30042;
assign x_61328 = x_61326 & x_61327;
assign x_61329 = x_61325 & x_61328;
assign x_61330 = x_61322 & x_61329;
assign x_61331 = x_61316 & x_61330;
assign x_61332 = x_30044 & x_30045;
assign x_61333 = x_30043 & x_61332;
assign x_61334 = x_30046 & x_30047;
assign x_61335 = x_30048 & x_30049;
assign x_61336 = x_61334 & x_61335;
assign x_61337 = x_61333 & x_61336;
assign x_61338 = x_30050 & x_30051;
assign x_61339 = x_30052 & x_30053;
assign x_61340 = x_61338 & x_61339;
assign x_61341 = x_30054 & x_30055;
assign x_61342 = x_30056 & x_30057;
assign x_61343 = x_61341 & x_61342;
assign x_61344 = x_61340 & x_61343;
assign x_61345 = x_61337 & x_61344;
assign x_61346 = x_30058 & x_30059;
assign x_61347 = x_30060 & x_30061;
assign x_61348 = x_61346 & x_61347;
assign x_61349 = x_30062 & x_30063;
assign x_61350 = x_30064 & x_30065;
assign x_61351 = x_61349 & x_61350;
assign x_61352 = x_61348 & x_61351;
assign x_61353 = x_30066 & x_30067;
assign x_61354 = x_30068 & x_30069;
assign x_61355 = x_61353 & x_61354;
assign x_61356 = x_30070 & x_30071;
assign x_61357 = x_30072 & x_30073;
assign x_61358 = x_61356 & x_61357;
assign x_61359 = x_61355 & x_61358;
assign x_61360 = x_61352 & x_61359;
assign x_61361 = x_61345 & x_61360;
assign x_61362 = x_61331 & x_61361;
assign x_61363 = x_61302 & x_61362;
assign x_61364 = x_61242 & x_61363;
assign x_61365 = x_30075 & x_30076;
assign x_61366 = x_30074 & x_61365;
assign x_61367 = x_30077 & x_30078;
assign x_61368 = x_30079 & x_30080;
assign x_61369 = x_61367 & x_61368;
assign x_61370 = x_61366 & x_61369;
assign x_61371 = x_30081 & x_30082;
assign x_61372 = x_30083 & x_30084;
assign x_61373 = x_61371 & x_61372;
assign x_61374 = x_30085 & x_30086;
assign x_61375 = x_30087 & x_30088;
assign x_61376 = x_61374 & x_61375;
assign x_61377 = x_61373 & x_61376;
assign x_61378 = x_61370 & x_61377;
assign x_61379 = x_30090 & x_30091;
assign x_61380 = x_30089 & x_61379;
assign x_61381 = x_30092 & x_30093;
assign x_61382 = x_30094 & x_30095;
assign x_61383 = x_61381 & x_61382;
assign x_61384 = x_61380 & x_61383;
assign x_61385 = x_30096 & x_30097;
assign x_61386 = x_30098 & x_30099;
assign x_61387 = x_61385 & x_61386;
assign x_61388 = x_30100 & x_30101;
assign x_61389 = x_30102 & x_30103;
assign x_61390 = x_61388 & x_61389;
assign x_61391 = x_61387 & x_61390;
assign x_61392 = x_61384 & x_61391;
assign x_61393 = x_61378 & x_61392;
assign x_61394 = x_30105 & x_30106;
assign x_61395 = x_30104 & x_61394;
assign x_61396 = x_30107 & x_30108;
assign x_61397 = x_30109 & x_30110;
assign x_61398 = x_61396 & x_61397;
assign x_61399 = x_61395 & x_61398;
assign x_61400 = x_30111 & x_30112;
assign x_61401 = x_30113 & x_30114;
assign x_61402 = x_61400 & x_61401;
assign x_61403 = x_30115 & x_30116;
assign x_61404 = x_30117 & x_30118;
assign x_61405 = x_61403 & x_61404;
assign x_61406 = x_61402 & x_61405;
assign x_61407 = x_61399 & x_61406;
assign x_61408 = x_30119 & x_30120;
assign x_61409 = x_30121 & x_30122;
assign x_61410 = x_61408 & x_61409;
assign x_61411 = x_30123 & x_30124;
assign x_61412 = x_30125 & x_30126;
assign x_61413 = x_61411 & x_61412;
assign x_61414 = x_61410 & x_61413;
assign x_61415 = x_30127 & x_30128;
assign x_61416 = x_30129 & x_30130;
assign x_61417 = x_61415 & x_61416;
assign x_61418 = x_30131 & x_30132;
assign x_61419 = x_30133 & x_30134;
assign x_61420 = x_61418 & x_61419;
assign x_61421 = x_61417 & x_61420;
assign x_61422 = x_61414 & x_61421;
assign x_61423 = x_61407 & x_61422;
assign x_61424 = x_61393 & x_61423;
assign x_61425 = x_30136 & x_30137;
assign x_61426 = x_30135 & x_61425;
assign x_61427 = x_30138 & x_30139;
assign x_61428 = x_30140 & x_30141;
assign x_61429 = x_61427 & x_61428;
assign x_61430 = x_61426 & x_61429;
assign x_61431 = x_30142 & x_30143;
assign x_61432 = x_30144 & x_30145;
assign x_61433 = x_61431 & x_61432;
assign x_61434 = x_30146 & x_30147;
assign x_61435 = x_30148 & x_30149;
assign x_61436 = x_61434 & x_61435;
assign x_61437 = x_61433 & x_61436;
assign x_61438 = x_61430 & x_61437;
assign x_61439 = x_30151 & x_30152;
assign x_61440 = x_30150 & x_61439;
assign x_61441 = x_30153 & x_30154;
assign x_61442 = x_30155 & x_30156;
assign x_61443 = x_61441 & x_61442;
assign x_61444 = x_61440 & x_61443;
assign x_61445 = x_30157 & x_30158;
assign x_61446 = x_30159 & x_30160;
assign x_61447 = x_61445 & x_61446;
assign x_61448 = x_30161 & x_30162;
assign x_61449 = x_30163 & x_30164;
assign x_61450 = x_61448 & x_61449;
assign x_61451 = x_61447 & x_61450;
assign x_61452 = x_61444 & x_61451;
assign x_61453 = x_61438 & x_61452;
assign x_61454 = x_30166 & x_30167;
assign x_61455 = x_30165 & x_61454;
assign x_61456 = x_30168 & x_30169;
assign x_61457 = x_30170 & x_30171;
assign x_61458 = x_61456 & x_61457;
assign x_61459 = x_61455 & x_61458;
assign x_61460 = x_30172 & x_30173;
assign x_61461 = x_30174 & x_30175;
assign x_61462 = x_61460 & x_61461;
assign x_61463 = x_30176 & x_30177;
assign x_61464 = x_30178 & x_30179;
assign x_61465 = x_61463 & x_61464;
assign x_61466 = x_61462 & x_61465;
assign x_61467 = x_61459 & x_61466;
assign x_61468 = x_30180 & x_30181;
assign x_61469 = x_30182 & x_30183;
assign x_61470 = x_61468 & x_61469;
assign x_61471 = x_30184 & x_30185;
assign x_61472 = x_30186 & x_30187;
assign x_61473 = x_61471 & x_61472;
assign x_61474 = x_61470 & x_61473;
assign x_61475 = x_30188 & x_30189;
assign x_61476 = x_30190 & x_30191;
assign x_61477 = x_61475 & x_61476;
assign x_61478 = x_30192 & x_30193;
assign x_61479 = x_30194 & x_30195;
assign x_61480 = x_61478 & x_61479;
assign x_61481 = x_61477 & x_61480;
assign x_61482 = x_61474 & x_61481;
assign x_61483 = x_61467 & x_61482;
assign x_61484 = x_61453 & x_61483;
assign x_61485 = x_61424 & x_61484;
assign x_61486 = x_30197 & x_30198;
assign x_61487 = x_30196 & x_61486;
assign x_61488 = x_30199 & x_30200;
assign x_61489 = x_30201 & x_30202;
assign x_61490 = x_61488 & x_61489;
assign x_61491 = x_61487 & x_61490;
assign x_61492 = x_30203 & x_30204;
assign x_61493 = x_30205 & x_30206;
assign x_61494 = x_61492 & x_61493;
assign x_61495 = x_30207 & x_30208;
assign x_61496 = x_30209 & x_30210;
assign x_61497 = x_61495 & x_61496;
assign x_61498 = x_61494 & x_61497;
assign x_61499 = x_61491 & x_61498;
assign x_61500 = x_30212 & x_30213;
assign x_61501 = x_30211 & x_61500;
assign x_61502 = x_30214 & x_30215;
assign x_61503 = x_30216 & x_30217;
assign x_61504 = x_61502 & x_61503;
assign x_61505 = x_61501 & x_61504;
assign x_61506 = x_30218 & x_30219;
assign x_61507 = x_30220 & x_30221;
assign x_61508 = x_61506 & x_61507;
assign x_61509 = x_30222 & x_30223;
assign x_61510 = x_30224 & x_30225;
assign x_61511 = x_61509 & x_61510;
assign x_61512 = x_61508 & x_61511;
assign x_61513 = x_61505 & x_61512;
assign x_61514 = x_61499 & x_61513;
assign x_61515 = x_30227 & x_30228;
assign x_61516 = x_30226 & x_61515;
assign x_61517 = x_30229 & x_30230;
assign x_61518 = x_30231 & x_30232;
assign x_61519 = x_61517 & x_61518;
assign x_61520 = x_61516 & x_61519;
assign x_61521 = x_30233 & x_30234;
assign x_61522 = x_30235 & x_30236;
assign x_61523 = x_61521 & x_61522;
assign x_61524 = x_30237 & x_30238;
assign x_61525 = x_30239 & x_30240;
assign x_61526 = x_61524 & x_61525;
assign x_61527 = x_61523 & x_61526;
assign x_61528 = x_61520 & x_61527;
assign x_61529 = x_30241 & x_30242;
assign x_61530 = x_30243 & x_30244;
assign x_61531 = x_61529 & x_61530;
assign x_61532 = x_30245 & x_30246;
assign x_61533 = x_30247 & x_30248;
assign x_61534 = x_61532 & x_61533;
assign x_61535 = x_61531 & x_61534;
assign x_61536 = x_30249 & x_30250;
assign x_61537 = x_30251 & x_30252;
assign x_61538 = x_61536 & x_61537;
assign x_61539 = x_30253 & x_30254;
assign x_61540 = x_30255 & x_30256;
assign x_61541 = x_61539 & x_61540;
assign x_61542 = x_61538 & x_61541;
assign x_61543 = x_61535 & x_61542;
assign x_61544 = x_61528 & x_61543;
assign x_61545 = x_61514 & x_61544;
assign x_61546 = x_30258 & x_30259;
assign x_61547 = x_30257 & x_61546;
assign x_61548 = x_30260 & x_30261;
assign x_61549 = x_30262 & x_30263;
assign x_61550 = x_61548 & x_61549;
assign x_61551 = x_61547 & x_61550;
assign x_61552 = x_30264 & x_30265;
assign x_61553 = x_30266 & x_30267;
assign x_61554 = x_61552 & x_61553;
assign x_61555 = x_30268 & x_30269;
assign x_61556 = x_30270 & x_30271;
assign x_61557 = x_61555 & x_61556;
assign x_61558 = x_61554 & x_61557;
assign x_61559 = x_61551 & x_61558;
assign x_61560 = x_30272 & x_30273;
assign x_61561 = x_30274 & x_30275;
assign x_61562 = x_61560 & x_61561;
assign x_61563 = x_30276 & x_30277;
assign x_61564 = x_30278 & x_30279;
assign x_61565 = x_61563 & x_61564;
assign x_61566 = x_61562 & x_61565;
assign x_61567 = x_30280 & x_30281;
assign x_61568 = x_30282 & x_30283;
assign x_61569 = x_61567 & x_61568;
assign x_61570 = x_30284 & x_30285;
assign x_61571 = x_30286 & x_30287;
assign x_61572 = x_61570 & x_61571;
assign x_61573 = x_61569 & x_61572;
assign x_61574 = x_61566 & x_61573;
assign x_61575 = x_61559 & x_61574;
assign x_61576 = x_30289 & x_30290;
assign x_61577 = x_30288 & x_61576;
assign x_61578 = x_30291 & x_30292;
assign x_61579 = x_30293 & x_30294;
assign x_61580 = x_61578 & x_61579;
assign x_61581 = x_61577 & x_61580;
assign x_61582 = x_30295 & x_30296;
assign x_61583 = x_30297 & x_30298;
assign x_61584 = x_61582 & x_61583;
assign x_61585 = x_30299 & x_30300;
assign x_61586 = x_30301 & x_30302;
assign x_61587 = x_61585 & x_61586;
assign x_61588 = x_61584 & x_61587;
assign x_61589 = x_61581 & x_61588;
assign x_61590 = x_30303 & x_30304;
assign x_61591 = x_30305 & x_30306;
assign x_61592 = x_61590 & x_61591;
assign x_61593 = x_30307 & x_30308;
assign x_61594 = x_30309 & x_30310;
assign x_61595 = x_61593 & x_61594;
assign x_61596 = x_61592 & x_61595;
assign x_61597 = x_30311 & x_30312;
assign x_61598 = x_30313 & x_30314;
assign x_61599 = x_61597 & x_61598;
assign x_61600 = x_30315 & x_30316;
assign x_61601 = x_30317 & x_30318;
assign x_61602 = x_61600 & x_61601;
assign x_61603 = x_61599 & x_61602;
assign x_61604 = x_61596 & x_61603;
assign x_61605 = x_61589 & x_61604;
assign x_61606 = x_61575 & x_61605;
assign x_61607 = x_61545 & x_61606;
assign x_61608 = x_61485 & x_61607;
assign x_61609 = x_61364 & x_61608;
assign x_61610 = x_61121 & x_61609;
assign x_61611 = x_30320 & x_30321;
assign x_61612 = x_30319 & x_61611;
assign x_61613 = x_30322 & x_30323;
assign x_61614 = x_30324 & x_30325;
assign x_61615 = x_61613 & x_61614;
assign x_61616 = x_61612 & x_61615;
assign x_61617 = x_30326 & x_30327;
assign x_61618 = x_30328 & x_30329;
assign x_61619 = x_61617 & x_61618;
assign x_61620 = x_30330 & x_30331;
assign x_61621 = x_30332 & x_30333;
assign x_61622 = x_61620 & x_61621;
assign x_61623 = x_61619 & x_61622;
assign x_61624 = x_61616 & x_61623;
assign x_61625 = x_30335 & x_30336;
assign x_61626 = x_30334 & x_61625;
assign x_61627 = x_30337 & x_30338;
assign x_61628 = x_30339 & x_30340;
assign x_61629 = x_61627 & x_61628;
assign x_61630 = x_61626 & x_61629;
assign x_61631 = x_30341 & x_30342;
assign x_61632 = x_30343 & x_30344;
assign x_61633 = x_61631 & x_61632;
assign x_61634 = x_30345 & x_30346;
assign x_61635 = x_30347 & x_30348;
assign x_61636 = x_61634 & x_61635;
assign x_61637 = x_61633 & x_61636;
assign x_61638 = x_61630 & x_61637;
assign x_61639 = x_61624 & x_61638;
assign x_61640 = x_30350 & x_30351;
assign x_61641 = x_30349 & x_61640;
assign x_61642 = x_30352 & x_30353;
assign x_61643 = x_30354 & x_30355;
assign x_61644 = x_61642 & x_61643;
assign x_61645 = x_61641 & x_61644;
assign x_61646 = x_30356 & x_30357;
assign x_61647 = x_30358 & x_30359;
assign x_61648 = x_61646 & x_61647;
assign x_61649 = x_30360 & x_30361;
assign x_61650 = x_30362 & x_30363;
assign x_61651 = x_61649 & x_61650;
assign x_61652 = x_61648 & x_61651;
assign x_61653 = x_61645 & x_61652;
assign x_61654 = x_30364 & x_30365;
assign x_61655 = x_30366 & x_30367;
assign x_61656 = x_61654 & x_61655;
assign x_61657 = x_30368 & x_30369;
assign x_61658 = x_30370 & x_30371;
assign x_61659 = x_61657 & x_61658;
assign x_61660 = x_61656 & x_61659;
assign x_61661 = x_30372 & x_30373;
assign x_61662 = x_30374 & x_30375;
assign x_61663 = x_61661 & x_61662;
assign x_61664 = x_30376 & x_30377;
assign x_61665 = x_30378 & x_30379;
assign x_61666 = x_61664 & x_61665;
assign x_61667 = x_61663 & x_61666;
assign x_61668 = x_61660 & x_61667;
assign x_61669 = x_61653 & x_61668;
assign x_61670 = x_61639 & x_61669;
assign x_61671 = x_30381 & x_30382;
assign x_61672 = x_30380 & x_61671;
assign x_61673 = x_30383 & x_30384;
assign x_61674 = x_30385 & x_30386;
assign x_61675 = x_61673 & x_61674;
assign x_61676 = x_61672 & x_61675;
assign x_61677 = x_30387 & x_30388;
assign x_61678 = x_30389 & x_30390;
assign x_61679 = x_61677 & x_61678;
assign x_61680 = x_30391 & x_30392;
assign x_61681 = x_30393 & x_30394;
assign x_61682 = x_61680 & x_61681;
assign x_61683 = x_61679 & x_61682;
assign x_61684 = x_61676 & x_61683;
assign x_61685 = x_30396 & x_30397;
assign x_61686 = x_30395 & x_61685;
assign x_61687 = x_30398 & x_30399;
assign x_61688 = x_30400 & x_30401;
assign x_61689 = x_61687 & x_61688;
assign x_61690 = x_61686 & x_61689;
assign x_61691 = x_30402 & x_30403;
assign x_61692 = x_30404 & x_30405;
assign x_61693 = x_61691 & x_61692;
assign x_61694 = x_30406 & x_30407;
assign x_61695 = x_30408 & x_30409;
assign x_61696 = x_61694 & x_61695;
assign x_61697 = x_61693 & x_61696;
assign x_61698 = x_61690 & x_61697;
assign x_61699 = x_61684 & x_61698;
assign x_61700 = x_30411 & x_30412;
assign x_61701 = x_30410 & x_61700;
assign x_61702 = x_30413 & x_30414;
assign x_61703 = x_30415 & x_30416;
assign x_61704 = x_61702 & x_61703;
assign x_61705 = x_61701 & x_61704;
assign x_61706 = x_30417 & x_30418;
assign x_61707 = x_30419 & x_30420;
assign x_61708 = x_61706 & x_61707;
assign x_61709 = x_30421 & x_30422;
assign x_61710 = x_30423 & x_30424;
assign x_61711 = x_61709 & x_61710;
assign x_61712 = x_61708 & x_61711;
assign x_61713 = x_61705 & x_61712;
assign x_61714 = x_30425 & x_30426;
assign x_61715 = x_30427 & x_30428;
assign x_61716 = x_61714 & x_61715;
assign x_61717 = x_30429 & x_30430;
assign x_61718 = x_30431 & x_30432;
assign x_61719 = x_61717 & x_61718;
assign x_61720 = x_61716 & x_61719;
assign x_61721 = x_30433 & x_30434;
assign x_61722 = x_30435 & x_30436;
assign x_61723 = x_61721 & x_61722;
assign x_61724 = x_30437 & x_30438;
assign x_61725 = x_30439 & x_30440;
assign x_61726 = x_61724 & x_61725;
assign x_61727 = x_61723 & x_61726;
assign x_61728 = x_61720 & x_61727;
assign x_61729 = x_61713 & x_61728;
assign x_61730 = x_61699 & x_61729;
assign x_61731 = x_61670 & x_61730;
assign x_61732 = x_30442 & x_30443;
assign x_61733 = x_30441 & x_61732;
assign x_61734 = x_30444 & x_30445;
assign x_61735 = x_30446 & x_30447;
assign x_61736 = x_61734 & x_61735;
assign x_61737 = x_61733 & x_61736;
assign x_61738 = x_30448 & x_30449;
assign x_61739 = x_30450 & x_30451;
assign x_61740 = x_61738 & x_61739;
assign x_61741 = x_30452 & x_30453;
assign x_61742 = x_30454 & x_30455;
assign x_61743 = x_61741 & x_61742;
assign x_61744 = x_61740 & x_61743;
assign x_61745 = x_61737 & x_61744;
assign x_61746 = x_30457 & x_30458;
assign x_61747 = x_30456 & x_61746;
assign x_61748 = x_30459 & x_30460;
assign x_61749 = x_30461 & x_30462;
assign x_61750 = x_61748 & x_61749;
assign x_61751 = x_61747 & x_61750;
assign x_61752 = x_30463 & x_30464;
assign x_61753 = x_30465 & x_30466;
assign x_61754 = x_61752 & x_61753;
assign x_61755 = x_30467 & x_30468;
assign x_61756 = x_30469 & x_30470;
assign x_61757 = x_61755 & x_61756;
assign x_61758 = x_61754 & x_61757;
assign x_61759 = x_61751 & x_61758;
assign x_61760 = x_61745 & x_61759;
assign x_61761 = x_30472 & x_30473;
assign x_61762 = x_30471 & x_61761;
assign x_61763 = x_30474 & x_30475;
assign x_61764 = x_30476 & x_30477;
assign x_61765 = x_61763 & x_61764;
assign x_61766 = x_61762 & x_61765;
assign x_61767 = x_30478 & x_30479;
assign x_61768 = x_30480 & x_30481;
assign x_61769 = x_61767 & x_61768;
assign x_61770 = x_30482 & x_30483;
assign x_61771 = x_30484 & x_30485;
assign x_61772 = x_61770 & x_61771;
assign x_61773 = x_61769 & x_61772;
assign x_61774 = x_61766 & x_61773;
assign x_61775 = x_30486 & x_30487;
assign x_61776 = x_30488 & x_30489;
assign x_61777 = x_61775 & x_61776;
assign x_61778 = x_30490 & x_30491;
assign x_61779 = x_30492 & x_30493;
assign x_61780 = x_61778 & x_61779;
assign x_61781 = x_61777 & x_61780;
assign x_61782 = x_30494 & x_30495;
assign x_61783 = x_30496 & x_30497;
assign x_61784 = x_61782 & x_61783;
assign x_61785 = x_30498 & x_30499;
assign x_61786 = x_30500 & x_30501;
assign x_61787 = x_61785 & x_61786;
assign x_61788 = x_61784 & x_61787;
assign x_61789 = x_61781 & x_61788;
assign x_61790 = x_61774 & x_61789;
assign x_61791 = x_61760 & x_61790;
assign x_61792 = x_30503 & x_30504;
assign x_61793 = x_30502 & x_61792;
assign x_61794 = x_30505 & x_30506;
assign x_61795 = x_30507 & x_30508;
assign x_61796 = x_61794 & x_61795;
assign x_61797 = x_61793 & x_61796;
assign x_61798 = x_30509 & x_30510;
assign x_61799 = x_30511 & x_30512;
assign x_61800 = x_61798 & x_61799;
assign x_61801 = x_30513 & x_30514;
assign x_61802 = x_30515 & x_30516;
assign x_61803 = x_61801 & x_61802;
assign x_61804 = x_61800 & x_61803;
assign x_61805 = x_61797 & x_61804;
assign x_61806 = x_30518 & x_30519;
assign x_61807 = x_30517 & x_61806;
assign x_61808 = x_30520 & x_30521;
assign x_61809 = x_30522 & x_30523;
assign x_61810 = x_61808 & x_61809;
assign x_61811 = x_61807 & x_61810;
assign x_61812 = x_30524 & x_30525;
assign x_61813 = x_30526 & x_30527;
assign x_61814 = x_61812 & x_61813;
assign x_61815 = x_30528 & x_30529;
assign x_61816 = x_30530 & x_30531;
assign x_61817 = x_61815 & x_61816;
assign x_61818 = x_61814 & x_61817;
assign x_61819 = x_61811 & x_61818;
assign x_61820 = x_61805 & x_61819;
assign x_61821 = x_30533 & x_30534;
assign x_61822 = x_30532 & x_61821;
assign x_61823 = x_30535 & x_30536;
assign x_61824 = x_30537 & x_30538;
assign x_61825 = x_61823 & x_61824;
assign x_61826 = x_61822 & x_61825;
assign x_61827 = x_30539 & x_30540;
assign x_61828 = x_30541 & x_30542;
assign x_61829 = x_61827 & x_61828;
assign x_61830 = x_30543 & x_30544;
assign x_61831 = x_30545 & x_30546;
assign x_61832 = x_61830 & x_61831;
assign x_61833 = x_61829 & x_61832;
assign x_61834 = x_61826 & x_61833;
assign x_61835 = x_30547 & x_30548;
assign x_61836 = x_30549 & x_30550;
assign x_61837 = x_61835 & x_61836;
assign x_61838 = x_30551 & x_30552;
assign x_61839 = x_30553 & x_30554;
assign x_61840 = x_61838 & x_61839;
assign x_61841 = x_61837 & x_61840;
assign x_61842 = x_30555 & x_30556;
assign x_61843 = x_30557 & x_30558;
assign x_61844 = x_61842 & x_61843;
assign x_61845 = x_30559 & x_30560;
assign x_61846 = x_30561 & x_30562;
assign x_61847 = x_61845 & x_61846;
assign x_61848 = x_61844 & x_61847;
assign x_61849 = x_61841 & x_61848;
assign x_61850 = x_61834 & x_61849;
assign x_61851 = x_61820 & x_61850;
assign x_61852 = x_61791 & x_61851;
assign x_61853 = x_61731 & x_61852;
assign x_61854 = x_30564 & x_30565;
assign x_61855 = x_30563 & x_61854;
assign x_61856 = x_30566 & x_30567;
assign x_61857 = x_30568 & x_30569;
assign x_61858 = x_61856 & x_61857;
assign x_61859 = x_61855 & x_61858;
assign x_61860 = x_30570 & x_30571;
assign x_61861 = x_30572 & x_30573;
assign x_61862 = x_61860 & x_61861;
assign x_61863 = x_30574 & x_30575;
assign x_61864 = x_30576 & x_30577;
assign x_61865 = x_61863 & x_61864;
assign x_61866 = x_61862 & x_61865;
assign x_61867 = x_61859 & x_61866;
assign x_61868 = x_30579 & x_30580;
assign x_61869 = x_30578 & x_61868;
assign x_61870 = x_30581 & x_30582;
assign x_61871 = x_30583 & x_30584;
assign x_61872 = x_61870 & x_61871;
assign x_61873 = x_61869 & x_61872;
assign x_61874 = x_30585 & x_30586;
assign x_61875 = x_30587 & x_30588;
assign x_61876 = x_61874 & x_61875;
assign x_61877 = x_30589 & x_30590;
assign x_61878 = x_30591 & x_30592;
assign x_61879 = x_61877 & x_61878;
assign x_61880 = x_61876 & x_61879;
assign x_61881 = x_61873 & x_61880;
assign x_61882 = x_61867 & x_61881;
assign x_61883 = x_30594 & x_30595;
assign x_61884 = x_30593 & x_61883;
assign x_61885 = x_30596 & x_30597;
assign x_61886 = x_30598 & x_30599;
assign x_61887 = x_61885 & x_61886;
assign x_61888 = x_61884 & x_61887;
assign x_61889 = x_30600 & x_30601;
assign x_61890 = x_30602 & x_30603;
assign x_61891 = x_61889 & x_61890;
assign x_61892 = x_30604 & x_30605;
assign x_61893 = x_30606 & x_30607;
assign x_61894 = x_61892 & x_61893;
assign x_61895 = x_61891 & x_61894;
assign x_61896 = x_61888 & x_61895;
assign x_61897 = x_30608 & x_30609;
assign x_61898 = x_30610 & x_30611;
assign x_61899 = x_61897 & x_61898;
assign x_61900 = x_30612 & x_30613;
assign x_61901 = x_30614 & x_30615;
assign x_61902 = x_61900 & x_61901;
assign x_61903 = x_61899 & x_61902;
assign x_61904 = x_30616 & x_30617;
assign x_61905 = x_30618 & x_30619;
assign x_61906 = x_61904 & x_61905;
assign x_61907 = x_30620 & x_30621;
assign x_61908 = x_30622 & x_30623;
assign x_61909 = x_61907 & x_61908;
assign x_61910 = x_61906 & x_61909;
assign x_61911 = x_61903 & x_61910;
assign x_61912 = x_61896 & x_61911;
assign x_61913 = x_61882 & x_61912;
assign x_61914 = x_30625 & x_30626;
assign x_61915 = x_30624 & x_61914;
assign x_61916 = x_30627 & x_30628;
assign x_61917 = x_30629 & x_30630;
assign x_61918 = x_61916 & x_61917;
assign x_61919 = x_61915 & x_61918;
assign x_61920 = x_30631 & x_30632;
assign x_61921 = x_30633 & x_30634;
assign x_61922 = x_61920 & x_61921;
assign x_61923 = x_30635 & x_30636;
assign x_61924 = x_30637 & x_30638;
assign x_61925 = x_61923 & x_61924;
assign x_61926 = x_61922 & x_61925;
assign x_61927 = x_61919 & x_61926;
assign x_61928 = x_30640 & x_30641;
assign x_61929 = x_30639 & x_61928;
assign x_61930 = x_30642 & x_30643;
assign x_61931 = x_30644 & x_30645;
assign x_61932 = x_61930 & x_61931;
assign x_61933 = x_61929 & x_61932;
assign x_61934 = x_30646 & x_30647;
assign x_61935 = x_30648 & x_30649;
assign x_61936 = x_61934 & x_61935;
assign x_61937 = x_30650 & x_30651;
assign x_61938 = x_30652 & x_30653;
assign x_61939 = x_61937 & x_61938;
assign x_61940 = x_61936 & x_61939;
assign x_61941 = x_61933 & x_61940;
assign x_61942 = x_61927 & x_61941;
assign x_61943 = x_30655 & x_30656;
assign x_61944 = x_30654 & x_61943;
assign x_61945 = x_30657 & x_30658;
assign x_61946 = x_30659 & x_30660;
assign x_61947 = x_61945 & x_61946;
assign x_61948 = x_61944 & x_61947;
assign x_61949 = x_30661 & x_30662;
assign x_61950 = x_30663 & x_30664;
assign x_61951 = x_61949 & x_61950;
assign x_61952 = x_30665 & x_30666;
assign x_61953 = x_30667 & x_30668;
assign x_61954 = x_61952 & x_61953;
assign x_61955 = x_61951 & x_61954;
assign x_61956 = x_61948 & x_61955;
assign x_61957 = x_30669 & x_30670;
assign x_61958 = x_30671 & x_30672;
assign x_61959 = x_61957 & x_61958;
assign x_61960 = x_30673 & x_30674;
assign x_61961 = x_30675 & x_30676;
assign x_61962 = x_61960 & x_61961;
assign x_61963 = x_61959 & x_61962;
assign x_61964 = x_30677 & x_30678;
assign x_61965 = x_30679 & x_30680;
assign x_61966 = x_61964 & x_61965;
assign x_61967 = x_30681 & x_30682;
assign x_61968 = x_30683 & x_30684;
assign x_61969 = x_61967 & x_61968;
assign x_61970 = x_61966 & x_61969;
assign x_61971 = x_61963 & x_61970;
assign x_61972 = x_61956 & x_61971;
assign x_61973 = x_61942 & x_61972;
assign x_61974 = x_61913 & x_61973;
assign x_61975 = x_30686 & x_30687;
assign x_61976 = x_30685 & x_61975;
assign x_61977 = x_30688 & x_30689;
assign x_61978 = x_30690 & x_30691;
assign x_61979 = x_61977 & x_61978;
assign x_61980 = x_61976 & x_61979;
assign x_61981 = x_30692 & x_30693;
assign x_61982 = x_30694 & x_30695;
assign x_61983 = x_61981 & x_61982;
assign x_61984 = x_30696 & x_30697;
assign x_61985 = x_30698 & x_30699;
assign x_61986 = x_61984 & x_61985;
assign x_61987 = x_61983 & x_61986;
assign x_61988 = x_61980 & x_61987;
assign x_61989 = x_30701 & x_30702;
assign x_61990 = x_30700 & x_61989;
assign x_61991 = x_30703 & x_30704;
assign x_61992 = x_30705 & x_30706;
assign x_61993 = x_61991 & x_61992;
assign x_61994 = x_61990 & x_61993;
assign x_61995 = x_30707 & x_30708;
assign x_61996 = x_30709 & x_30710;
assign x_61997 = x_61995 & x_61996;
assign x_61998 = x_30711 & x_30712;
assign x_61999 = x_30713 & x_30714;
assign x_62000 = x_61998 & x_61999;
assign x_62001 = x_61997 & x_62000;
assign x_62002 = x_61994 & x_62001;
assign x_62003 = x_61988 & x_62002;
assign x_62004 = x_30716 & x_30717;
assign x_62005 = x_30715 & x_62004;
assign x_62006 = x_30718 & x_30719;
assign x_62007 = x_30720 & x_30721;
assign x_62008 = x_62006 & x_62007;
assign x_62009 = x_62005 & x_62008;
assign x_62010 = x_30722 & x_30723;
assign x_62011 = x_30724 & x_30725;
assign x_62012 = x_62010 & x_62011;
assign x_62013 = x_30726 & x_30727;
assign x_62014 = x_30728 & x_30729;
assign x_62015 = x_62013 & x_62014;
assign x_62016 = x_62012 & x_62015;
assign x_62017 = x_62009 & x_62016;
assign x_62018 = x_30730 & x_30731;
assign x_62019 = x_30732 & x_30733;
assign x_62020 = x_62018 & x_62019;
assign x_62021 = x_30734 & x_30735;
assign x_62022 = x_30736 & x_30737;
assign x_62023 = x_62021 & x_62022;
assign x_62024 = x_62020 & x_62023;
assign x_62025 = x_30738 & x_30739;
assign x_62026 = x_30740 & x_30741;
assign x_62027 = x_62025 & x_62026;
assign x_62028 = x_30742 & x_30743;
assign x_62029 = x_30744 & x_30745;
assign x_62030 = x_62028 & x_62029;
assign x_62031 = x_62027 & x_62030;
assign x_62032 = x_62024 & x_62031;
assign x_62033 = x_62017 & x_62032;
assign x_62034 = x_62003 & x_62033;
assign x_62035 = x_30747 & x_30748;
assign x_62036 = x_30746 & x_62035;
assign x_62037 = x_30749 & x_30750;
assign x_62038 = x_30751 & x_30752;
assign x_62039 = x_62037 & x_62038;
assign x_62040 = x_62036 & x_62039;
assign x_62041 = x_30753 & x_30754;
assign x_62042 = x_30755 & x_30756;
assign x_62043 = x_62041 & x_62042;
assign x_62044 = x_30757 & x_30758;
assign x_62045 = x_30759 & x_30760;
assign x_62046 = x_62044 & x_62045;
assign x_62047 = x_62043 & x_62046;
assign x_62048 = x_62040 & x_62047;
assign x_62049 = x_30761 & x_30762;
assign x_62050 = x_30763 & x_30764;
assign x_62051 = x_62049 & x_62050;
assign x_62052 = x_30765 & x_30766;
assign x_62053 = x_30767 & x_30768;
assign x_62054 = x_62052 & x_62053;
assign x_62055 = x_62051 & x_62054;
assign x_62056 = x_30769 & x_30770;
assign x_62057 = x_30771 & x_30772;
assign x_62058 = x_62056 & x_62057;
assign x_62059 = x_30773 & x_30774;
assign x_62060 = x_30775 & x_30776;
assign x_62061 = x_62059 & x_62060;
assign x_62062 = x_62058 & x_62061;
assign x_62063 = x_62055 & x_62062;
assign x_62064 = x_62048 & x_62063;
assign x_62065 = x_30778 & x_30779;
assign x_62066 = x_30777 & x_62065;
assign x_62067 = x_30780 & x_30781;
assign x_62068 = x_30782 & x_30783;
assign x_62069 = x_62067 & x_62068;
assign x_62070 = x_62066 & x_62069;
assign x_62071 = x_30784 & x_30785;
assign x_62072 = x_30786 & x_30787;
assign x_62073 = x_62071 & x_62072;
assign x_62074 = x_30788 & x_30789;
assign x_62075 = x_30790 & x_30791;
assign x_62076 = x_62074 & x_62075;
assign x_62077 = x_62073 & x_62076;
assign x_62078 = x_62070 & x_62077;
assign x_62079 = x_30792 & x_30793;
assign x_62080 = x_30794 & x_30795;
assign x_62081 = x_62079 & x_62080;
assign x_62082 = x_30796 & x_30797;
assign x_62083 = x_30798 & x_30799;
assign x_62084 = x_62082 & x_62083;
assign x_62085 = x_62081 & x_62084;
assign x_62086 = x_30800 & x_30801;
assign x_62087 = x_30802 & x_30803;
assign x_62088 = x_62086 & x_62087;
assign x_62089 = x_30804 & x_30805;
assign x_62090 = x_30806 & x_30807;
assign x_62091 = x_62089 & x_62090;
assign x_62092 = x_62088 & x_62091;
assign x_62093 = x_62085 & x_62092;
assign x_62094 = x_62078 & x_62093;
assign x_62095 = x_62064 & x_62094;
assign x_62096 = x_62034 & x_62095;
assign x_62097 = x_61974 & x_62096;
assign x_62098 = x_61853 & x_62097;
assign x_62099 = x_30809 & x_30810;
assign x_62100 = x_30808 & x_62099;
assign x_62101 = x_30811 & x_30812;
assign x_62102 = x_30813 & x_30814;
assign x_62103 = x_62101 & x_62102;
assign x_62104 = x_62100 & x_62103;
assign x_62105 = x_30815 & x_30816;
assign x_62106 = x_30817 & x_30818;
assign x_62107 = x_62105 & x_62106;
assign x_62108 = x_30819 & x_30820;
assign x_62109 = x_30821 & x_30822;
assign x_62110 = x_62108 & x_62109;
assign x_62111 = x_62107 & x_62110;
assign x_62112 = x_62104 & x_62111;
assign x_62113 = x_30824 & x_30825;
assign x_62114 = x_30823 & x_62113;
assign x_62115 = x_30826 & x_30827;
assign x_62116 = x_30828 & x_30829;
assign x_62117 = x_62115 & x_62116;
assign x_62118 = x_62114 & x_62117;
assign x_62119 = x_30830 & x_30831;
assign x_62120 = x_30832 & x_30833;
assign x_62121 = x_62119 & x_62120;
assign x_62122 = x_30834 & x_30835;
assign x_62123 = x_30836 & x_30837;
assign x_62124 = x_62122 & x_62123;
assign x_62125 = x_62121 & x_62124;
assign x_62126 = x_62118 & x_62125;
assign x_62127 = x_62112 & x_62126;
assign x_62128 = x_30839 & x_30840;
assign x_62129 = x_30838 & x_62128;
assign x_62130 = x_30841 & x_30842;
assign x_62131 = x_30843 & x_30844;
assign x_62132 = x_62130 & x_62131;
assign x_62133 = x_62129 & x_62132;
assign x_62134 = x_30845 & x_30846;
assign x_62135 = x_30847 & x_30848;
assign x_62136 = x_62134 & x_62135;
assign x_62137 = x_30849 & x_30850;
assign x_62138 = x_30851 & x_30852;
assign x_62139 = x_62137 & x_62138;
assign x_62140 = x_62136 & x_62139;
assign x_62141 = x_62133 & x_62140;
assign x_62142 = x_30853 & x_30854;
assign x_62143 = x_30855 & x_30856;
assign x_62144 = x_62142 & x_62143;
assign x_62145 = x_30857 & x_30858;
assign x_62146 = x_30859 & x_30860;
assign x_62147 = x_62145 & x_62146;
assign x_62148 = x_62144 & x_62147;
assign x_62149 = x_30861 & x_30862;
assign x_62150 = x_30863 & x_30864;
assign x_62151 = x_62149 & x_62150;
assign x_62152 = x_30865 & x_30866;
assign x_62153 = x_30867 & x_30868;
assign x_62154 = x_62152 & x_62153;
assign x_62155 = x_62151 & x_62154;
assign x_62156 = x_62148 & x_62155;
assign x_62157 = x_62141 & x_62156;
assign x_62158 = x_62127 & x_62157;
assign x_62159 = x_30870 & x_30871;
assign x_62160 = x_30869 & x_62159;
assign x_62161 = x_30872 & x_30873;
assign x_62162 = x_30874 & x_30875;
assign x_62163 = x_62161 & x_62162;
assign x_62164 = x_62160 & x_62163;
assign x_62165 = x_30876 & x_30877;
assign x_62166 = x_30878 & x_30879;
assign x_62167 = x_62165 & x_62166;
assign x_62168 = x_30880 & x_30881;
assign x_62169 = x_30882 & x_30883;
assign x_62170 = x_62168 & x_62169;
assign x_62171 = x_62167 & x_62170;
assign x_62172 = x_62164 & x_62171;
assign x_62173 = x_30885 & x_30886;
assign x_62174 = x_30884 & x_62173;
assign x_62175 = x_30887 & x_30888;
assign x_62176 = x_30889 & x_30890;
assign x_62177 = x_62175 & x_62176;
assign x_62178 = x_62174 & x_62177;
assign x_62179 = x_30891 & x_30892;
assign x_62180 = x_30893 & x_30894;
assign x_62181 = x_62179 & x_62180;
assign x_62182 = x_30895 & x_30896;
assign x_62183 = x_30897 & x_30898;
assign x_62184 = x_62182 & x_62183;
assign x_62185 = x_62181 & x_62184;
assign x_62186 = x_62178 & x_62185;
assign x_62187 = x_62172 & x_62186;
assign x_62188 = x_30900 & x_30901;
assign x_62189 = x_30899 & x_62188;
assign x_62190 = x_30902 & x_30903;
assign x_62191 = x_30904 & x_30905;
assign x_62192 = x_62190 & x_62191;
assign x_62193 = x_62189 & x_62192;
assign x_62194 = x_30906 & x_30907;
assign x_62195 = x_30908 & x_30909;
assign x_62196 = x_62194 & x_62195;
assign x_62197 = x_30910 & x_30911;
assign x_62198 = x_30912 & x_30913;
assign x_62199 = x_62197 & x_62198;
assign x_62200 = x_62196 & x_62199;
assign x_62201 = x_62193 & x_62200;
assign x_62202 = x_30914 & x_30915;
assign x_62203 = x_30916 & x_30917;
assign x_62204 = x_62202 & x_62203;
assign x_62205 = x_30918 & x_30919;
assign x_62206 = x_30920 & x_30921;
assign x_62207 = x_62205 & x_62206;
assign x_62208 = x_62204 & x_62207;
assign x_62209 = x_30922 & x_30923;
assign x_62210 = x_30924 & x_30925;
assign x_62211 = x_62209 & x_62210;
assign x_62212 = x_30926 & x_30927;
assign x_62213 = x_30928 & x_30929;
assign x_62214 = x_62212 & x_62213;
assign x_62215 = x_62211 & x_62214;
assign x_62216 = x_62208 & x_62215;
assign x_62217 = x_62201 & x_62216;
assign x_62218 = x_62187 & x_62217;
assign x_62219 = x_62158 & x_62218;
assign x_62220 = x_30931 & x_30932;
assign x_62221 = x_30930 & x_62220;
assign x_62222 = x_30933 & x_30934;
assign x_62223 = x_30935 & x_30936;
assign x_62224 = x_62222 & x_62223;
assign x_62225 = x_62221 & x_62224;
assign x_62226 = x_30937 & x_30938;
assign x_62227 = x_30939 & x_30940;
assign x_62228 = x_62226 & x_62227;
assign x_62229 = x_30941 & x_30942;
assign x_62230 = x_30943 & x_30944;
assign x_62231 = x_62229 & x_62230;
assign x_62232 = x_62228 & x_62231;
assign x_62233 = x_62225 & x_62232;
assign x_62234 = x_30946 & x_30947;
assign x_62235 = x_30945 & x_62234;
assign x_62236 = x_30948 & x_30949;
assign x_62237 = x_30950 & x_30951;
assign x_62238 = x_62236 & x_62237;
assign x_62239 = x_62235 & x_62238;
assign x_62240 = x_30952 & x_30953;
assign x_62241 = x_30954 & x_30955;
assign x_62242 = x_62240 & x_62241;
assign x_62243 = x_30956 & x_30957;
assign x_62244 = x_30958 & x_30959;
assign x_62245 = x_62243 & x_62244;
assign x_62246 = x_62242 & x_62245;
assign x_62247 = x_62239 & x_62246;
assign x_62248 = x_62233 & x_62247;
assign x_62249 = x_30961 & x_30962;
assign x_62250 = x_30960 & x_62249;
assign x_62251 = x_30963 & x_30964;
assign x_62252 = x_30965 & x_30966;
assign x_62253 = x_62251 & x_62252;
assign x_62254 = x_62250 & x_62253;
assign x_62255 = x_30967 & x_30968;
assign x_62256 = x_30969 & x_30970;
assign x_62257 = x_62255 & x_62256;
assign x_62258 = x_30971 & x_30972;
assign x_62259 = x_30973 & x_30974;
assign x_62260 = x_62258 & x_62259;
assign x_62261 = x_62257 & x_62260;
assign x_62262 = x_62254 & x_62261;
assign x_62263 = x_30975 & x_30976;
assign x_62264 = x_30977 & x_30978;
assign x_62265 = x_62263 & x_62264;
assign x_62266 = x_30979 & x_30980;
assign x_62267 = x_30981 & x_30982;
assign x_62268 = x_62266 & x_62267;
assign x_62269 = x_62265 & x_62268;
assign x_62270 = x_30983 & x_30984;
assign x_62271 = x_30985 & x_30986;
assign x_62272 = x_62270 & x_62271;
assign x_62273 = x_30987 & x_30988;
assign x_62274 = x_30989 & x_30990;
assign x_62275 = x_62273 & x_62274;
assign x_62276 = x_62272 & x_62275;
assign x_62277 = x_62269 & x_62276;
assign x_62278 = x_62262 & x_62277;
assign x_62279 = x_62248 & x_62278;
assign x_62280 = x_30992 & x_30993;
assign x_62281 = x_30991 & x_62280;
assign x_62282 = x_30994 & x_30995;
assign x_62283 = x_30996 & x_30997;
assign x_62284 = x_62282 & x_62283;
assign x_62285 = x_62281 & x_62284;
assign x_62286 = x_30998 & x_30999;
assign x_62287 = x_31000 & x_31001;
assign x_62288 = x_62286 & x_62287;
assign x_62289 = x_31002 & x_31003;
assign x_62290 = x_31004 & x_31005;
assign x_62291 = x_62289 & x_62290;
assign x_62292 = x_62288 & x_62291;
assign x_62293 = x_62285 & x_62292;
assign x_62294 = x_31006 & x_31007;
assign x_62295 = x_31008 & x_31009;
assign x_62296 = x_62294 & x_62295;
assign x_62297 = x_31010 & x_31011;
assign x_62298 = x_31012 & x_31013;
assign x_62299 = x_62297 & x_62298;
assign x_62300 = x_62296 & x_62299;
assign x_62301 = x_31014 & x_31015;
assign x_62302 = x_31016 & x_31017;
assign x_62303 = x_62301 & x_62302;
assign x_62304 = x_31018 & x_31019;
assign x_62305 = x_31020 & x_31021;
assign x_62306 = x_62304 & x_62305;
assign x_62307 = x_62303 & x_62306;
assign x_62308 = x_62300 & x_62307;
assign x_62309 = x_62293 & x_62308;
assign x_62310 = x_31023 & x_31024;
assign x_62311 = x_31022 & x_62310;
assign x_62312 = x_31025 & x_31026;
assign x_62313 = x_31027 & x_31028;
assign x_62314 = x_62312 & x_62313;
assign x_62315 = x_62311 & x_62314;
assign x_62316 = x_31029 & x_31030;
assign x_62317 = x_31031 & x_31032;
assign x_62318 = x_62316 & x_62317;
assign x_62319 = x_31033 & x_31034;
assign x_62320 = x_31035 & x_31036;
assign x_62321 = x_62319 & x_62320;
assign x_62322 = x_62318 & x_62321;
assign x_62323 = x_62315 & x_62322;
assign x_62324 = x_31037 & x_31038;
assign x_62325 = x_31039 & x_31040;
assign x_62326 = x_62324 & x_62325;
assign x_62327 = x_31041 & x_31042;
assign x_62328 = x_31043 & x_31044;
assign x_62329 = x_62327 & x_62328;
assign x_62330 = x_62326 & x_62329;
assign x_62331 = x_31045 & x_31046;
assign x_62332 = x_31047 & x_31048;
assign x_62333 = x_62331 & x_62332;
assign x_62334 = x_31049 & x_31050;
assign x_62335 = x_31051 & x_31052;
assign x_62336 = x_62334 & x_62335;
assign x_62337 = x_62333 & x_62336;
assign x_62338 = x_62330 & x_62337;
assign x_62339 = x_62323 & x_62338;
assign x_62340 = x_62309 & x_62339;
assign x_62341 = x_62279 & x_62340;
assign x_62342 = x_62219 & x_62341;
assign x_62343 = x_31054 & x_31055;
assign x_62344 = x_31053 & x_62343;
assign x_62345 = x_31056 & x_31057;
assign x_62346 = x_31058 & x_31059;
assign x_62347 = x_62345 & x_62346;
assign x_62348 = x_62344 & x_62347;
assign x_62349 = x_31060 & x_31061;
assign x_62350 = x_31062 & x_31063;
assign x_62351 = x_62349 & x_62350;
assign x_62352 = x_31064 & x_31065;
assign x_62353 = x_31066 & x_31067;
assign x_62354 = x_62352 & x_62353;
assign x_62355 = x_62351 & x_62354;
assign x_62356 = x_62348 & x_62355;
assign x_62357 = x_31069 & x_31070;
assign x_62358 = x_31068 & x_62357;
assign x_62359 = x_31071 & x_31072;
assign x_62360 = x_31073 & x_31074;
assign x_62361 = x_62359 & x_62360;
assign x_62362 = x_62358 & x_62361;
assign x_62363 = x_31075 & x_31076;
assign x_62364 = x_31077 & x_31078;
assign x_62365 = x_62363 & x_62364;
assign x_62366 = x_31079 & x_31080;
assign x_62367 = x_31081 & x_31082;
assign x_62368 = x_62366 & x_62367;
assign x_62369 = x_62365 & x_62368;
assign x_62370 = x_62362 & x_62369;
assign x_62371 = x_62356 & x_62370;
assign x_62372 = x_31084 & x_31085;
assign x_62373 = x_31083 & x_62372;
assign x_62374 = x_31086 & x_31087;
assign x_62375 = x_31088 & x_31089;
assign x_62376 = x_62374 & x_62375;
assign x_62377 = x_62373 & x_62376;
assign x_62378 = x_31090 & x_31091;
assign x_62379 = x_31092 & x_31093;
assign x_62380 = x_62378 & x_62379;
assign x_62381 = x_31094 & x_31095;
assign x_62382 = x_31096 & x_31097;
assign x_62383 = x_62381 & x_62382;
assign x_62384 = x_62380 & x_62383;
assign x_62385 = x_62377 & x_62384;
assign x_62386 = x_31098 & x_31099;
assign x_62387 = x_31100 & x_31101;
assign x_62388 = x_62386 & x_62387;
assign x_62389 = x_31102 & x_31103;
assign x_62390 = x_31104 & x_31105;
assign x_62391 = x_62389 & x_62390;
assign x_62392 = x_62388 & x_62391;
assign x_62393 = x_31106 & x_31107;
assign x_62394 = x_31108 & x_31109;
assign x_62395 = x_62393 & x_62394;
assign x_62396 = x_31110 & x_31111;
assign x_62397 = x_31112 & x_31113;
assign x_62398 = x_62396 & x_62397;
assign x_62399 = x_62395 & x_62398;
assign x_62400 = x_62392 & x_62399;
assign x_62401 = x_62385 & x_62400;
assign x_62402 = x_62371 & x_62401;
assign x_62403 = x_31115 & x_31116;
assign x_62404 = x_31114 & x_62403;
assign x_62405 = x_31117 & x_31118;
assign x_62406 = x_31119 & x_31120;
assign x_62407 = x_62405 & x_62406;
assign x_62408 = x_62404 & x_62407;
assign x_62409 = x_31121 & x_31122;
assign x_62410 = x_31123 & x_31124;
assign x_62411 = x_62409 & x_62410;
assign x_62412 = x_31125 & x_31126;
assign x_62413 = x_31127 & x_31128;
assign x_62414 = x_62412 & x_62413;
assign x_62415 = x_62411 & x_62414;
assign x_62416 = x_62408 & x_62415;
assign x_62417 = x_31130 & x_31131;
assign x_62418 = x_31129 & x_62417;
assign x_62419 = x_31132 & x_31133;
assign x_62420 = x_31134 & x_31135;
assign x_62421 = x_62419 & x_62420;
assign x_62422 = x_62418 & x_62421;
assign x_62423 = x_31136 & x_31137;
assign x_62424 = x_31138 & x_31139;
assign x_62425 = x_62423 & x_62424;
assign x_62426 = x_31140 & x_31141;
assign x_62427 = x_31142 & x_31143;
assign x_62428 = x_62426 & x_62427;
assign x_62429 = x_62425 & x_62428;
assign x_62430 = x_62422 & x_62429;
assign x_62431 = x_62416 & x_62430;
assign x_62432 = x_31145 & x_31146;
assign x_62433 = x_31144 & x_62432;
assign x_62434 = x_31147 & x_31148;
assign x_62435 = x_31149 & x_31150;
assign x_62436 = x_62434 & x_62435;
assign x_62437 = x_62433 & x_62436;
assign x_62438 = x_31151 & x_31152;
assign x_62439 = x_31153 & x_31154;
assign x_62440 = x_62438 & x_62439;
assign x_62441 = x_31155 & x_31156;
assign x_62442 = x_31157 & x_31158;
assign x_62443 = x_62441 & x_62442;
assign x_62444 = x_62440 & x_62443;
assign x_62445 = x_62437 & x_62444;
assign x_62446 = x_31159 & x_31160;
assign x_62447 = x_31161 & x_31162;
assign x_62448 = x_62446 & x_62447;
assign x_62449 = x_31163 & x_31164;
assign x_62450 = x_31165 & x_31166;
assign x_62451 = x_62449 & x_62450;
assign x_62452 = x_62448 & x_62451;
assign x_62453 = x_31167 & x_31168;
assign x_62454 = x_31169 & x_31170;
assign x_62455 = x_62453 & x_62454;
assign x_62456 = x_31171 & x_31172;
assign x_62457 = x_31173 & x_31174;
assign x_62458 = x_62456 & x_62457;
assign x_62459 = x_62455 & x_62458;
assign x_62460 = x_62452 & x_62459;
assign x_62461 = x_62445 & x_62460;
assign x_62462 = x_62431 & x_62461;
assign x_62463 = x_62402 & x_62462;
assign x_62464 = x_31176 & x_31177;
assign x_62465 = x_31175 & x_62464;
assign x_62466 = x_31178 & x_31179;
assign x_62467 = x_31180 & x_31181;
assign x_62468 = x_62466 & x_62467;
assign x_62469 = x_62465 & x_62468;
assign x_62470 = x_31182 & x_31183;
assign x_62471 = x_31184 & x_31185;
assign x_62472 = x_62470 & x_62471;
assign x_62473 = x_31186 & x_31187;
assign x_62474 = x_31188 & x_31189;
assign x_62475 = x_62473 & x_62474;
assign x_62476 = x_62472 & x_62475;
assign x_62477 = x_62469 & x_62476;
assign x_62478 = x_31191 & x_31192;
assign x_62479 = x_31190 & x_62478;
assign x_62480 = x_31193 & x_31194;
assign x_62481 = x_31195 & x_31196;
assign x_62482 = x_62480 & x_62481;
assign x_62483 = x_62479 & x_62482;
assign x_62484 = x_31197 & x_31198;
assign x_62485 = x_31199 & x_31200;
assign x_62486 = x_62484 & x_62485;
assign x_62487 = x_31201 & x_31202;
assign x_62488 = x_31203 & x_31204;
assign x_62489 = x_62487 & x_62488;
assign x_62490 = x_62486 & x_62489;
assign x_62491 = x_62483 & x_62490;
assign x_62492 = x_62477 & x_62491;
assign x_62493 = x_31206 & x_31207;
assign x_62494 = x_31205 & x_62493;
assign x_62495 = x_31208 & x_31209;
assign x_62496 = x_31210 & x_31211;
assign x_62497 = x_62495 & x_62496;
assign x_62498 = x_62494 & x_62497;
assign x_62499 = x_31212 & x_31213;
assign x_62500 = x_31214 & x_31215;
assign x_62501 = x_62499 & x_62500;
assign x_62502 = x_31216 & x_31217;
assign x_62503 = x_31218 & x_31219;
assign x_62504 = x_62502 & x_62503;
assign x_62505 = x_62501 & x_62504;
assign x_62506 = x_62498 & x_62505;
assign x_62507 = x_31220 & x_31221;
assign x_62508 = x_31222 & x_31223;
assign x_62509 = x_62507 & x_62508;
assign x_62510 = x_31224 & x_31225;
assign x_62511 = x_31226 & x_31227;
assign x_62512 = x_62510 & x_62511;
assign x_62513 = x_62509 & x_62512;
assign x_62514 = x_31228 & x_31229;
assign x_62515 = x_31230 & x_31231;
assign x_62516 = x_62514 & x_62515;
assign x_62517 = x_31232 & x_31233;
assign x_62518 = x_31234 & x_31235;
assign x_62519 = x_62517 & x_62518;
assign x_62520 = x_62516 & x_62519;
assign x_62521 = x_62513 & x_62520;
assign x_62522 = x_62506 & x_62521;
assign x_62523 = x_62492 & x_62522;
assign x_62524 = x_31237 & x_31238;
assign x_62525 = x_31236 & x_62524;
assign x_62526 = x_31239 & x_31240;
assign x_62527 = x_31241 & x_31242;
assign x_62528 = x_62526 & x_62527;
assign x_62529 = x_62525 & x_62528;
assign x_62530 = x_31243 & x_31244;
assign x_62531 = x_31245 & x_31246;
assign x_62532 = x_62530 & x_62531;
assign x_62533 = x_31247 & x_31248;
assign x_62534 = x_31249 & x_31250;
assign x_62535 = x_62533 & x_62534;
assign x_62536 = x_62532 & x_62535;
assign x_62537 = x_62529 & x_62536;
assign x_62538 = x_31251 & x_31252;
assign x_62539 = x_31253 & x_31254;
assign x_62540 = x_62538 & x_62539;
assign x_62541 = x_31255 & x_31256;
assign x_62542 = x_31257 & x_31258;
assign x_62543 = x_62541 & x_62542;
assign x_62544 = x_62540 & x_62543;
assign x_62545 = x_31259 & x_31260;
assign x_62546 = x_31261 & x_31262;
assign x_62547 = x_62545 & x_62546;
assign x_62548 = x_31263 & x_31264;
assign x_62549 = x_31265 & x_31266;
assign x_62550 = x_62548 & x_62549;
assign x_62551 = x_62547 & x_62550;
assign x_62552 = x_62544 & x_62551;
assign x_62553 = x_62537 & x_62552;
assign x_62554 = x_31268 & x_31269;
assign x_62555 = x_31267 & x_62554;
assign x_62556 = x_31270 & x_31271;
assign x_62557 = x_31272 & x_31273;
assign x_62558 = x_62556 & x_62557;
assign x_62559 = x_62555 & x_62558;
assign x_62560 = x_31274 & x_31275;
assign x_62561 = x_31276 & x_31277;
assign x_62562 = x_62560 & x_62561;
assign x_62563 = x_31278 & x_31279;
assign x_62564 = x_31280 & x_31281;
assign x_62565 = x_62563 & x_62564;
assign x_62566 = x_62562 & x_62565;
assign x_62567 = x_62559 & x_62566;
assign x_62568 = x_31282 & x_31283;
assign x_62569 = x_31284 & x_31285;
assign x_62570 = x_62568 & x_62569;
assign x_62571 = x_31286 & x_31287;
assign x_62572 = x_31288 & x_31289;
assign x_62573 = x_62571 & x_62572;
assign x_62574 = x_62570 & x_62573;
assign x_62575 = x_31290 & x_31291;
assign x_62576 = x_31292 & x_31293;
assign x_62577 = x_62575 & x_62576;
assign x_62578 = x_31294 & x_31295;
assign x_62579 = x_31296 & x_31297;
assign x_62580 = x_62578 & x_62579;
assign x_62581 = x_62577 & x_62580;
assign x_62582 = x_62574 & x_62581;
assign x_62583 = x_62567 & x_62582;
assign x_62584 = x_62553 & x_62583;
assign x_62585 = x_62523 & x_62584;
assign x_62586 = x_62463 & x_62585;
assign x_62587 = x_62342 & x_62586;
assign x_62588 = x_62098 & x_62587;
assign x_62589 = x_61610 & x_62588;
assign x_62590 = x_60633 & x_62589;
assign x_62591 = x_58678 & x_62590;
assign x_62592 = x_54767 & x_62591;
assign x_62593 = x_46944 & x_62592;
assign o_1 = x_62593;
endmodule
