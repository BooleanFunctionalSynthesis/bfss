// Verilog file written by procedure writeCombinationalCircuitInVerilog
//Skolem functions to be generated for i_ variables
module bobtuint30neg_all_bit_differing_from_cycle ( i_1, i_2, i_3, i_4, i_5, i_6, i_7, i_8, i_9, i_10, i_11, i_12, i_13, i_14, i_15, i_16, i_17, i_18, i_19, i_20, i_21, i_22, i_23, i_24, i_25, i_26, i_27, i_28, i_29, i_30, i_31, i_32, i_33, i_34, i_35, i_36, i_37, i_38, i_39, i_40, i_41, i_42, i_43, i_44, i_45, i_46, i_47, i_48, i_49, i_50, i_51, i_52, i_53, i_54, i_55, i_56, i_57, i_58, i_59, i_60, i_61, i_62, i_63, i_64, i_65, i_66, i_67, i_68, i_69, i_70, i_71, i_72, i_73, i_74, i_75, i_76, i_77, i_78, i_79, i_80, i_81, i_82, i_83, i_84, i_85, i_86, i_87, i_88, i_89, i_90, i_91, i_92, i_93, i_94, i_95, i_96, i_97, i_98, i_99, i_100, i_101, i_102, i_103, i_104, i_105, i_106, i_107, i_108, i_109, i_110, i_111, i_112, i_113, i_114, i_115, i_116, i_117, i_118, i_119, i_120, i_121, i_122, i_123, i_124, i_125, i_126, i_127, i_128, i_129, i_130, i_131, i_132, i_133, i_134, i_135, i_136, i_137, i_138, i_139, i_140, i_141, i_142, i_143, i_144, i_145, i_146, i_147, i_148, i_149, i_150, i_151, i_152, i_153, i_154, i_155, i_156, i_157, i_158, i_159, i_160, i_161, i_162, i_163, i_164, i_165, i_166, i_167, i_168, i_169, i_170, i_171, i_172, i_173, i_174, i_175, i_176, i_177, i_178, i_179, i_180, i_181, i_182, i_183, i_184, i_185, i_186, i_187, i_188, i_189, i_190, i_191, i_192, i_193, i_194, i_195, i_196, i_197, i_198, i_199, i_200, i_201, i_202, i_203, i_204, i_205, i_206, i_207, i_208, i_209, i_210, i_211, i_212, i_213, x_214, x_215, x_216, x_217, x_218, x_219, x_220, x_221, x_222, x_223, x_224, x_225, x_226, x_227, x_228, x_229, x_230, x_231, x_232, x_233, x_234, x_235, x_236, x_237, x_238, x_239, x_240, x_241, x_242, x_243, x_244, x_245, x_246, x_247, x_248, x_249, x_250, x_251, x_252, x_253, x_254, x_255, x_256, x_257, x_258, x_259, x_260, x_261, x_262, x_263, x_264, x_265, x_266, x_267, x_268, x_269, x_270, x_271, x_272, x_273, x_274, x_275, x_276, x_277, x_278, x_279, x_280, x_281, x_282, x_283, x_284, x_285, x_286, x_287, x_288, x_289, x_290, x_291, x_292, x_293, x_294, x_295, x_296, x_297, x_298, x_299, x_300, x_301, x_302, x_303, x_304, x_305, x_306, x_307, x_308, x_309, x_310, x_311, x_312, x_313, x_314, x_315, x_316, x_317, x_318, x_319, x_320, x_321, x_322, x_323, x_324, x_325, x_326, x_327, x_328, x_329, x_330, x_331, x_332, x_333, x_334, x_335, x_336, x_337, x_338, x_339, x_340, x_341, x_342, x_343, x_344, x_345, x_346, x_347, x_348, x_349, x_350, x_351, x_352, x_353, x_354, x_355, x_356, x_357, x_358, x_359, x_360, x_361, x_362, x_363, x_364, x_365, x_366, x_367, x_368, x_369, x_370, x_371, x_372, x_373, x_374, x_375, x_376, x_377, x_378, x_379, x_380, x_381, x_382, x_383, x_384, x_385, x_386, x_387, x_388, x_389, x_390, x_391, x_392, x_393, x_394, x_395, x_396, x_397, x_398, x_399, x_400, x_401, x_402, x_403, x_404, x_405, x_406, x_407, x_408, x_409, x_410, x_411, x_412, x_413, x_414, x_415, x_416, x_417, x_418, x_419, x_420, x_421, x_422, x_423, x_424, x_425, x_426, x_427, x_428, x_429, x_430, x_431, x_432, x_433, x_434, x_435, x_436, x_437, x_438, x_439, x_440, x_441, x_442, x_443, x_444, x_445, x_446, x_447, x_448, x_449, x_450, x_451, x_452, x_453, x_454, x_455, x_456, x_457, x_458, x_459, x_460, x_461, x_462, x_463, x_464, x_465, x_466, x_467, x_468, x_469, x_470, x_471, x_472, x_473, x_474, x_475, x_476, x_477, x_478, x_479, x_480, x_481, x_482, x_483, x_484, x_485, x_486, x_487, x_488, x_489, x_490, x_491, x_492, x_493, x_494, x_495, x_496, x_497, x_498, x_499, x_500, x_501, x_502, x_503, x_504, x_505, x_506, x_507, x_508, x_509, x_510, x_511, x_512, x_513, x_514, x_515, x_516, x_517, x_518, x_519, x_520, x_521, x_522, x_523, x_524, x_525, x_526, x_527, x_528, x_529, x_530, x_531, x_532, x_533, x_534, x_535, x_536, x_537, x_538, x_539, x_540, x_541, x_542, x_543, x_544, x_545, x_546, x_547, x_548, x_549, x_550, x_551, x_552, x_553, x_554, x_555, x_556, x_557, x_558, x_559, x_560, x_561, x_562, x_563, x_564, x_565, x_566, x_567, x_568, x_569, x_570, x_571, x_572, x_573, x_574, x_575, x_576, x_577, x_578, x_579, x_580, x_581, x_582, x_583, x_584, x_585, x_586, x_587, x_588, x_589, x_590, x_591, x_592, x_593, x_594, x_595, x_596, x_597, x_598, x_599, x_600, x_601, x_602, x_603, x_604, x_605, x_606, x_607, x_608, x_609, x_610, x_611, x_612, x_613, x_614, x_615, x_616, x_617, x_618, x_619, x_620, x_621, x_622, x_623, x_624, x_625, x_626, x_627, x_628, x_629, x_630, x_631, x_632, x_633, x_634, x_635, x_636, x_637, o_1 );
input i_1;
input i_2;
input i_3;
input i_4;
input i_5;
input i_6;
input i_7;
input i_8;
input i_9;
input i_10;
input i_11;
input i_12;
input i_13;
input i_14;
input i_15;
input i_16;
input i_17;
input i_18;
input i_19;
input i_20;
input i_21;
input i_22;
input i_23;
input i_24;
input i_25;
input i_26;
input i_27;
input i_28;
input i_29;
input i_30;
input i_31;
input i_32;
input i_33;
input i_34;
input i_35;
input i_36;
input i_37;
input i_38;
input i_39;
input i_40;
input i_41;
input i_42;
input i_43;
input i_44;
input i_45;
input i_46;
input i_47;
input i_48;
input i_49;
input i_50;
input i_51;
input i_52;
input i_53;
input i_54;
input i_55;
input i_56;
input i_57;
input i_58;
input i_59;
input i_60;
input i_61;
input i_62;
input i_63;
input i_64;
input i_65;
input i_66;
input i_67;
input i_68;
input i_69;
input i_70;
input i_71;
input i_72;
input i_73;
input i_74;
input i_75;
input i_76;
input i_77;
input i_78;
input i_79;
input i_80;
input i_81;
input i_82;
input i_83;
input i_84;
input i_85;
input i_86;
input i_87;
input i_88;
input i_89;
input i_90;
input i_91;
input i_92;
input i_93;
input i_94;
input i_95;
input i_96;
input i_97;
input i_98;
input i_99;
input i_100;
input i_101;
input i_102;
input i_103;
input i_104;
input i_105;
input i_106;
input i_107;
input i_108;
input i_109;
input i_110;
input i_111;
input i_112;
input i_113;
input i_114;
input i_115;
input i_116;
input i_117;
input i_118;
input i_119;
input i_120;
input i_121;
input i_122;
input i_123;
input i_124;
input i_125;
input i_126;
input i_127;
input i_128;
input i_129;
input i_130;
input i_131;
input i_132;
input i_133;
input i_134;
input i_135;
input i_136;
input i_137;
input i_138;
input i_139;
input i_140;
input i_141;
input i_142;
input i_143;
input i_144;
input i_145;
input i_146;
input i_147;
input i_148;
input i_149;
input i_150;
input i_151;
input i_152;
input i_153;
input i_154;
input i_155;
input i_156;
input i_157;
input i_158;
input i_159;
input i_160;
input i_161;
input i_162;
input i_163;
input i_164;
input i_165;
input i_166;
input i_167;
input i_168;
input i_169;
input i_170;
input i_171;
input i_172;
input i_173;
input i_174;
input i_175;
input i_176;
input i_177;
input i_178;
input i_179;
input i_180;
input i_181;
input i_182;
input i_183;
input i_184;
input i_185;
input i_186;
input i_187;
input i_188;
input i_189;
input i_190;
input i_191;
input i_192;
input i_193;
input i_194;
input i_195;
input i_196;
input i_197;
input i_198;
input i_199;
input i_200;
input i_201;
input i_202;
input i_203;
input i_204;
input i_205;
input i_206;
input i_207;
input i_208;
input i_209;
input i_210;
input i_211;
input i_212;
input i_213;
input x_214;
input x_215;
input x_216;
input x_217;
input x_218;
input x_219;
input x_220;
input x_221;
input x_222;
input x_223;
input x_224;
input x_225;
input x_226;
input x_227;
input x_228;
input x_229;
input x_230;
input x_231;
input x_232;
input x_233;
input x_234;
input x_235;
input x_236;
input x_237;
input x_238;
input x_239;
input x_240;
input x_241;
input x_242;
input x_243;
input x_244;
input x_245;
input x_246;
input x_247;
input x_248;
input x_249;
input x_250;
input x_251;
input x_252;
input x_253;
input x_254;
input x_255;
input x_256;
input x_257;
input x_258;
input x_259;
input x_260;
input x_261;
input x_262;
input x_263;
input x_264;
input x_265;
input x_266;
input x_267;
input x_268;
input x_269;
input x_270;
input x_271;
input x_272;
input x_273;
input x_274;
input x_275;
input x_276;
input x_277;
input x_278;
input x_279;
input x_280;
input x_281;
input x_282;
input x_283;
input x_284;
input x_285;
input x_286;
input x_287;
input x_288;
input x_289;
input x_290;
input x_291;
input x_292;
input x_293;
input x_294;
input x_295;
input x_296;
input x_297;
input x_298;
input x_299;
input x_300;
input x_301;
input x_302;
input x_303;
input x_304;
input x_305;
input x_306;
input x_307;
input x_308;
input x_309;
input x_310;
input x_311;
input x_312;
input x_313;
input x_314;
input x_315;
input x_316;
input x_317;
input x_318;
input x_319;
input x_320;
input x_321;
input x_322;
input x_323;
input x_324;
input x_325;
input x_326;
input x_327;
input x_328;
input x_329;
input x_330;
input x_331;
input x_332;
input x_333;
input x_334;
input x_335;
input x_336;
input x_337;
input x_338;
input x_339;
input x_340;
input x_341;
input x_342;
input x_343;
input x_344;
input x_345;
input x_346;
input x_347;
input x_348;
input x_349;
input x_350;
input x_351;
input x_352;
input x_353;
input x_354;
input x_355;
input x_356;
input x_357;
input x_358;
input x_359;
input x_360;
input x_361;
input x_362;
input x_363;
input x_364;
input x_365;
input x_366;
input x_367;
input x_368;
input x_369;
input x_370;
input x_371;
input x_372;
input x_373;
input x_374;
input x_375;
input x_376;
input x_377;
input x_378;
input x_379;
input x_380;
input x_381;
input x_382;
input x_383;
input x_384;
input x_385;
input x_386;
input x_387;
input x_388;
input x_389;
input x_390;
input x_391;
input x_392;
input x_393;
input x_394;
input x_395;
input x_396;
input x_397;
input x_398;
input x_399;
input x_400;
input x_401;
input x_402;
input x_403;
input x_404;
input x_405;
input x_406;
input x_407;
input x_408;
input x_409;
input x_410;
input x_411;
input x_412;
input x_413;
input x_414;
input x_415;
input x_416;
input x_417;
input x_418;
input x_419;
input x_420;
input x_421;
input x_422;
input x_423;
input x_424;
input x_425;
input x_426;
input x_427;
input x_428;
input x_429;
input x_430;
input x_431;
input x_432;
input x_433;
input x_434;
input x_435;
input x_436;
input x_437;
input x_438;
input x_439;
input x_440;
input x_441;
input x_442;
input x_443;
input x_444;
input x_445;
input x_446;
input x_447;
input x_448;
input x_449;
input x_450;
input x_451;
input x_452;
input x_453;
input x_454;
input x_455;
input x_456;
input x_457;
input x_458;
input x_459;
input x_460;
input x_461;
input x_462;
input x_463;
input x_464;
input x_465;
input x_466;
input x_467;
input x_468;
input x_469;
input x_470;
input x_471;
input x_472;
input x_473;
input x_474;
input x_475;
input x_476;
input x_477;
input x_478;
input x_479;
input x_480;
input x_481;
input x_482;
input x_483;
input x_484;
input x_485;
input x_486;
input x_487;
input x_488;
input x_489;
input x_490;
input x_491;
input x_492;
input x_493;
input x_494;
input x_495;
input x_496;
input x_497;
input x_498;
input x_499;
input x_500;
input x_501;
input x_502;
input x_503;
input x_504;
input x_505;
input x_506;
input x_507;
input x_508;
input x_509;
input x_510;
input x_511;
input x_512;
input x_513;
input x_514;
input x_515;
input x_516;
input x_517;
input x_518;
input x_519;
input x_520;
input x_521;
input x_522;
input x_523;
input x_524;
input x_525;
input x_526;
input x_527;
input x_528;
input x_529;
input x_530;
input x_531;
input x_532;
input x_533;
input x_534;
input x_535;
input x_536;
input x_537;
input x_538;
input x_539;
input x_540;
input x_541;
input x_542;
input x_543;
input x_544;
input x_545;
input x_546;
input x_547;
input x_548;
input x_549;
input x_550;
input x_551;
input x_552;
input x_553;
input x_554;
input x_555;
input x_556;
input x_557;
input x_558;
input x_559;
input x_560;
input x_561;
input x_562;
input x_563;
input x_564;
input x_565;
input x_566;
input x_567;
input x_568;
input x_569;
input x_570;
input x_571;
input x_572;
input x_573;
input x_574;
input x_575;
input x_576;
input x_577;
input x_578;
input x_579;
input x_580;
input x_581;
input x_582;
input x_583;
input x_584;
input x_585;
input x_586;
input x_587;
input x_588;
input x_589;
input x_590;
input x_591;
input x_592;
input x_593;
input x_594;
input x_595;
input x_596;
input x_597;
input x_598;
input x_599;
input x_600;
input x_601;
input x_602;
input x_603;
input x_604;
input x_605;
input x_606;
input x_607;
input x_608;
input x_609;
input x_610;
input x_611;
input x_612;
input x_613;
input x_614;
input x_615;
input x_616;
input x_617;
input x_618;
input x_619;
input x_620;
input x_621;
input x_622;
input x_623;
input x_624;
input x_625;
input x_626;
input x_627;
input x_628;
input x_629;
input x_630;
input x_631;
input x_632;
input x_633;
input x_634;
input x_635;
input x_636;
input x_637;
output o_1;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_12;
wire n_13;
wire n_14;
wire n_15;
wire n_16;
wire n_17;
wire n_18;
wire n_19;
wire n_20;
wire n_21;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_27;
wire n_28;
wire n_29;
wire n_30;
wire n_31;
wire n_32;
wire n_33;
wire n_34;
wire n_35;
wire n_36;
wire n_37;
wire n_38;
wire n_39;
wire n_40;
wire n_41;
wire n_42;
wire n_43;
wire n_44;
wire n_45;
wire n_46;
wire n_47;
wire n_48;
wire n_49;
wire n_50;
wire n_51;
wire n_52;
wire n_53;
wire n_54;
wire n_55;
wire n_56;
wire n_57;
wire n_58;
wire n_59;
wire n_60;
wire n_61;
wire n_62;
wire n_63;
wire n_64;
wire n_65;
wire n_66;
wire n_67;
wire n_68;
wire n_69;
wire n_70;
wire n_71;
wire n_72;
wire n_73;
wire n_74;
wire n_75;
wire n_76;
wire n_77;
wire n_78;
wire n_79;
wire n_80;
wire n_81;
wire n_82;
wire n_83;
wire n_84;
wire n_85;
wire n_86;
wire n_87;
wire n_88;
wire n_89;
wire n_90;
wire n_91;
wire n_92;
wire n_93;
wire n_94;
wire n_95;
wire n_96;
wire n_97;
wire n_98;
wire n_99;
wire n_100;
wire n_101;
wire n_102;
wire n_103;
wire n_104;
wire n_105;
wire n_106;
wire n_107;
wire n_108;
wire n_109;
wire n_110;
wire n_111;
wire n_112;
wire n_113;
wire n_114;
wire n_115;
wire n_116;
wire n_117;
wire n_118;
wire n_119;
wire n_120;
wire n_121;
wire n_122;
wire n_123;
wire n_124;
wire n_125;
wire n_126;
wire n_127;
wire n_128;
wire n_129;
wire n_130;
wire n_131;
wire n_132;
wire n_133;
wire n_134;
wire n_135;
wire n_136;
wire n_137;
wire n_138;
wire n_139;
wire n_140;
wire n_141;
wire n_142;
wire n_143;
wire n_144;
wire n_145;
wire n_146;
wire n_147;
wire n_148;
wire n_149;
wire n_150;
wire n_151;
wire n_152;
wire n_153;
wire n_154;
wire n_155;
wire n_156;
wire n_157;
wire n_158;
wire n_159;
wire n_160;
wire n_161;
wire n_162;
wire n_163;
wire n_164;
wire n_165;
wire n_166;
wire n_167;
wire n_168;
wire n_169;
wire n_170;
wire n_171;
wire n_172;
wire n_173;
wire n_174;
wire n_175;
wire n_176;
wire n_177;
wire n_178;
wire n_179;
wire n_180;
wire n_181;
wire n_182;
wire n_183;
wire n_184;
wire n_185;
wire n_186;
wire n_187;
wire n_188;
wire n_189;
wire n_190;
wire n_191;
wire n_192;
wire n_193;
wire n_194;
wire n_195;
wire n_196;
wire n_197;
wire n_198;
wire n_199;
wire n_200;
wire n_201;
wire n_202;
wire n_203;
wire n_204;
wire n_205;
wire n_206;
wire n_207;
wire n_208;
wire n_209;
wire n_210;
wire n_211;
wire n_212;
wire n_213;
wire n_214;
wire n_215;
wire n_216;
wire n_217;
wire n_218;
wire n_219;
wire n_220;
wire n_221;
wire n_222;
wire n_223;
wire n_224;
wire n_225;
wire n_226;
wire n_227;
wire n_228;
wire n_229;
wire n_230;
wire n_231;
wire n_232;
wire n_233;
wire n_234;
wire n_235;
wire n_236;
wire n_237;
wire n_238;
wire n_239;
wire n_240;
wire n_241;
wire n_242;
wire n_243;
wire n_244;
wire n_245;
wire n_246;
wire n_247;
wire n_248;
wire n_249;
wire n_250;
wire n_251;
wire n_252;
wire n_253;
wire n_254;
wire n_255;
wire n_256;
wire n_257;
wire n_258;
wire n_259;
wire n_260;
wire n_261;
wire n_262;
wire n_263;
wire n_264;
wire n_265;
wire n_266;
wire n_267;
wire n_268;
wire n_269;
wire n_270;
wire n_271;
wire n_272;
wire n_273;
wire n_274;
wire n_275;
wire n_276;
wire n_277;
wire n_278;
wire n_279;
wire n_280;
wire n_281;
wire n_282;
wire n_283;
wire n_284;
wire n_285;
wire n_286;
wire n_287;
wire n_288;
wire n_289;
wire n_290;
wire n_291;
wire n_292;
wire n_293;
wire n_294;
wire n_295;
wire n_296;
wire n_297;
wire n_298;
wire n_299;
wire n_300;
wire n_301;
wire n_302;
wire n_303;
wire n_304;
wire n_305;
wire n_306;
wire n_307;
wire n_308;
wire n_309;
wire n_310;
wire n_311;
wire n_312;
wire n_313;
wire n_314;
wire n_315;
wire n_316;
wire n_317;
wire n_318;
wire n_319;
wire n_320;
wire n_321;
wire n_322;
wire n_323;
wire n_324;
wire n_325;
wire n_326;
wire n_327;
wire n_328;
wire n_329;
wire n_330;
wire n_331;
wire n_332;
wire n_333;
wire n_334;
wire n_335;
wire n_336;
wire n_337;
wire n_338;
wire n_339;
wire n_340;
wire n_341;
wire n_342;
wire n_343;
wire n_344;
wire n_345;
wire n_346;
wire n_347;
wire n_348;
wire n_349;
wire n_350;
wire n_351;
wire n_352;
wire n_353;
wire n_354;
wire n_355;
wire n_356;
wire n_357;
wire n_358;
wire n_359;
wire n_360;
wire n_361;
wire n_362;
wire n_363;
wire n_364;
wire n_365;
wire n_366;
wire n_367;
wire n_368;
wire n_369;
wire n_370;
wire n_371;
wire n_372;
wire n_373;
wire n_374;
wire n_375;
wire n_376;
wire n_377;
wire n_378;
wire n_379;
wire n_380;
wire n_381;
wire n_382;
wire n_383;
wire n_384;
wire n_385;
wire n_386;
wire n_387;
wire n_388;
wire n_389;
wire n_390;
wire n_391;
wire n_392;
wire n_393;
wire n_394;
wire n_395;
wire n_396;
wire n_397;
wire n_398;
wire n_399;
wire n_400;
wire n_401;
wire n_402;
wire n_403;
wire n_404;
wire n_405;
wire n_406;
wire n_407;
wire n_408;
wire n_409;
wire n_410;
wire n_411;
wire n_412;
wire n_413;
wire n_414;
wire n_415;
wire n_416;
wire n_417;
wire n_418;
wire n_419;
wire n_420;
wire n_421;
wire n_422;
wire n_423;
wire n_424;
wire n_425;
wire n_426;
wire n_427;
wire n_428;
wire n_429;
wire n_430;
wire n_431;
wire n_432;
wire n_433;
wire n_434;
wire n_435;
wire n_436;
wire n_437;
wire n_438;
wire n_439;
wire n_440;
wire n_441;
wire n_442;
wire n_443;
wire n_444;
wire n_445;
wire n_446;
wire n_447;
wire n_448;
wire n_449;
wire n_450;
wire n_451;
wire n_452;
wire n_453;
wire n_454;
wire n_455;
wire n_456;
wire n_457;
wire n_458;
wire n_459;
wire n_460;
wire n_461;
wire n_462;
wire n_463;
wire n_464;
wire n_465;
wire n_466;
wire n_467;
wire n_468;
wire n_469;
wire n_470;
wire n_471;
wire n_472;
wire n_473;
wire n_474;
wire n_475;
wire n_476;
wire n_477;
wire n_478;
wire n_479;
wire n_480;
wire n_481;
wire n_482;
wire n_483;
wire n_484;
wire n_485;
wire n_486;
wire n_487;
wire n_488;
wire n_489;
wire n_490;
wire n_491;
wire n_492;
wire n_493;
wire n_494;
wire n_495;
wire n_496;
wire n_497;
wire n_498;
wire n_499;
wire n_500;
wire n_501;
wire n_502;
wire n_503;
wire n_504;
wire n_505;
wire n_506;
wire n_507;
wire n_508;
wire n_509;
wire n_510;
wire n_511;
wire n_512;
wire n_513;
wire n_514;
wire n_515;
wire n_516;
wire n_517;
wire n_518;
wire n_519;
wire n_520;
wire n_521;
wire n_522;
wire n_523;
wire n_524;
wire n_525;
wire n_526;
wire n_527;
wire n_528;
wire n_529;
wire n_530;
wire n_531;
wire n_532;
wire n_533;
wire n_534;
wire n_535;
wire n_536;
wire n_537;
wire n_538;
wire n_539;
wire n_540;
wire n_541;
wire n_542;
wire n_543;
wire n_544;
wire n_545;
wire n_546;
wire n_547;
wire n_548;
wire n_549;
wire n_550;
wire n_551;
wire n_552;
wire n_553;
wire n_554;
wire n_555;
wire n_556;
wire n_557;
wire n_558;
wire n_559;
wire n_560;
wire n_561;
wire n_562;
wire n_563;
wire n_564;
wire n_565;
wire n_566;
wire n_567;
wire n_568;
wire n_569;
wire n_570;
wire n_571;
wire n_572;
wire n_573;
wire n_574;
wire n_575;
wire n_576;
wire n_577;
wire n_578;
wire n_579;
wire n_580;
wire n_581;
wire n_582;
wire n_583;
wire n_584;
wire n_585;
wire n_586;
wire n_587;
wire n_588;
wire n_589;
wire n_590;
wire n_591;
wire n_592;
wire n_593;
wire n_594;
wire n_595;
wire n_596;
wire n_597;
wire n_598;
wire n_599;
wire n_600;
wire n_601;
wire n_602;
wire n_603;
wire n_604;
wire n_605;
wire n_606;
wire n_607;
wire n_608;
wire n_609;
wire n_610;
wire n_611;
wire n_612;
wire n_613;
wire n_614;
wire n_615;
wire n_616;
wire n_617;
wire n_618;
wire n_619;
wire n_620;
wire n_621;
wire n_622;
wire n_623;
wire n_624;
wire n_625;
wire n_626;
wire n_627;
wire n_628;
wire n_629;
wire n_630;
wire n_631;
wire n_632;
wire n_633;
wire n_634;
wire n_635;
wire n_636;
wire n_637;
wire n_638;
wire n_639;
wire n_640;
wire n_641;
wire n_642;
wire n_643;
wire n_644;
wire n_645;
wire n_646;
wire n_647;
wire n_648;
wire n_649;
wire n_650;
wire n_651;
wire n_652;
wire n_653;
wire n_654;
wire n_655;
wire n_656;
wire n_657;
wire n_658;
wire n_659;
wire n_660;
wire n_661;
wire n_662;
wire n_663;
wire n_664;
wire n_665;
wire n_666;
wire n_667;
wire n_668;
wire n_669;
wire n_670;
wire n_671;
wire n_672;
wire n_673;
wire n_674;
wire n_675;
wire n_676;
wire n_677;
wire n_678;
wire n_679;
wire n_680;
wire n_681;
wire n_682;
wire n_683;
wire n_684;
wire n_685;
wire n_686;
wire n_687;
wire n_688;
wire n_689;
wire n_690;
wire n_691;
wire n_692;
wire n_693;
wire n_694;
wire n_695;
wire n_696;
wire n_697;
wire n_698;
wire n_699;
wire n_700;
wire n_701;
wire n_702;
wire n_703;
wire n_704;
wire n_705;
wire n_706;
wire n_707;
wire n_708;
wire n_709;
wire n_710;
wire n_711;
wire n_712;
wire n_713;
wire n_714;
wire n_715;
wire n_716;
wire n_717;
wire n_718;
wire n_719;
wire n_720;
wire n_721;
wire n_722;
wire n_723;
wire n_724;
wire n_725;
wire n_726;
wire n_727;
wire n_728;
wire n_729;
wire n_730;
wire n_731;
wire n_732;
wire n_733;
wire n_734;
wire n_735;
wire n_736;
wire n_737;
wire n_738;
wire n_739;
wire n_740;
wire n_741;
wire n_742;
wire n_743;
wire n_744;
wire n_745;
wire n_746;
wire n_747;
wire n_748;
wire n_749;
wire n_750;
wire n_751;
wire n_752;
wire n_753;
wire n_754;
wire n_755;
wire n_756;
wire n_757;
wire n_758;
wire n_759;
wire n_760;
wire n_761;
wire n_762;
wire n_763;
wire n_764;
wire n_765;
wire n_766;
wire n_767;
wire n_768;
wire n_769;
wire n_770;
wire n_771;
wire n_772;
wire n_773;
wire n_774;
wire n_775;
wire n_776;
wire n_777;
wire n_778;
wire n_779;
wire n_780;
wire n_781;
wire n_782;
wire n_783;
wire n_784;
wire n_785;
wire n_786;
wire n_787;
wire n_788;
wire n_789;
wire n_790;
wire n_791;
wire n_792;
wire n_793;
wire n_794;
wire n_795;
wire n_796;
wire n_797;
wire n_798;
wire n_799;
wire n_800;
wire n_801;
wire n_802;
wire n_803;
wire n_804;
wire n_805;
wire n_806;
wire n_807;
wire n_808;
wire n_809;
wire n_810;
wire n_811;
wire n_812;
wire n_813;
wire n_814;
wire n_815;
wire n_816;
wire n_817;
wire n_818;
wire n_819;
wire n_820;
wire n_821;
wire n_822;
wire n_823;
wire n_824;
wire n_825;
wire n_826;
wire n_827;
wire n_828;
wire n_829;
wire n_830;
wire n_831;
wire n_832;
wire n_833;
wire n_834;
wire n_835;
wire n_836;
wire n_837;
wire n_838;
wire n_839;
wire n_840;
wire n_841;
wire n_842;
wire n_843;
wire n_844;
wire n_845;
wire n_846;
wire n_847;
wire n_848;
wire n_849;
wire n_850;
wire n_851;
wire n_852;
wire n_853;
wire n_854;
wire n_855;
wire n_856;
wire n_857;
wire n_858;
wire n_859;
wire n_860;
wire n_861;
wire n_862;
wire n_863;
wire n_864;
wire n_865;
wire n_866;
wire n_867;
wire n_868;
wire n_869;
wire n_870;
wire n_871;
wire n_872;
wire n_873;
wire n_874;
wire n_875;
wire n_876;
wire n_877;
wire n_878;
wire n_879;
wire n_880;
wire n_881;
wire n_882;
wire n_883;
wire n_884;
wire n_885;
wire n_886;
wire n_887;
wire n_888;
wire n_889;
wire n_890;
wire n_891;
wire n_892;
wire n_893;
wire n_894;
wire n_895;
wire n_896;
wire n_897;
wire n_898;
wire n_899;
wire n_900;
wire n_901;
wire n_902;
wire n_903;
wire n_904;
wire n_905;
wire n_906;
wire n_907;
wire n_908;
wire n_909;
wire n_910;
wire n_911;
wire n_912;
wire n_913;
wire n_914;
wire n_915;
wire n_916;
wire n_917;
wire n_918;
wire n_919;
wire n_920;
wire n_921;
wire n_922;
wire n_923;
wire n_924;
wire n_925;
wire n_926;
wire n_927;
wire n_928;
wire n_929;
wire n_930;
wire n_931;
wire n_932;
wire n_933;
wire n_934;
wire n_935;
wire n_936;
wire n_937;
wire n_938;
wire n_939;
wire n_940;
wire n_941;
wire n_942;
wire n_943;
wire n_944;
wire n_945;
wire n_946;
wire n_947;
wire n_948;
wire n_949;
wire n_950;
wire n_951;
wire n_952;
wire n_953;
wire n_954;
wire n_955;
wire n_956;
wire n_957;
wire n_958;
wire n_959;
wire n_960;
wire n_961;
wire n_962;
wire n_963;
wire n_964;
wire n_965;
wire n_966;
wire n_967;
wire n_968;
wire n_969;
wire n_970;
wire n_971;
wire n_972;
wire n_973;
wire n_974;
wire n_975;
wire n_976;
wire n_977;
wire n_978;
wire n_979;
wire n_980;
wire n_981;
wire n_982;
wire n_983;
wire n_984;
wire n_985;
wire n_986;
wire n_987;
wire n_988;
wire n_989;
wire n_990;
wire n_991;
wire n_992;
wire n_993;
wire n_994;
wire n_995;
wire n_996;
wire n_997;
wire n_998;
wire n_999;
wire n_1000;
wire n_1001;
wire n_1002;
wire n_1003;
wire n_1004;
wire n_1005;
wire n_1006;
wire n_1007;
wire n_1008;
wire n_1009;
wire n_1010;
wire n_1011;
wire n_1012;
wire n_1013;
wire n_1014;
wire n_1015;
wire n_1016;
wire n_1017;
wire n_1018;
wire n_1019;
wire n_1020;
wire n_1021;
wire n_1022;
wire n_1023;
wire n_1024;
wire n_1025;
wire n_1026;
wire n_1027;
wire n_1028;
wire n_1029;
wire n_1030;
wire n_1031;
wire n_1032;
wire n_1033;
wire n_1034;
wire n_1035;
wire n_1036;
wire n_1037;
wire n_1038;
wire n_1039;
wire n_1040;
wire n_1041;
wire n_1042;
wire n_1043;
wire n_1044;
wire n_1045;
wire n_1046;
wire n_1047;
wire n_1048;
wire n_1049;
wire n_1050;
wire n_1051;
wire n_1052;
wire n_1053;
wire n_1054;
wire n_1055;
wire n_1056;
wire n_1057;
wire n_1058;
wire n_1059;
wire n_1060;
wire n_1061;
wire n_1062;
wire n_1063;
wire n_1064;
wire n_1065;
wire n_1066;
wire n_1067;
wire n_1068;
wire n_1069;
wire n_1070;
wire n_1071;
wire n_1072;
wire n_1073;
wire n_1074;
wire n_1075;
wire n_1076;
wire n_1077;
wire n_1078;
wire n_1079;
wire n_1080;
wire n_1081;
wire n_1082;
wire n_1083;
wire n_1084;
wire n_1085;
wire n_1086;
wire n_1087;
wire n_1088;
wire n_1089;
wire n_1090;
wire n_1091;
wire n_1092;
wire n_1093;
wire n_1094;
wire n_1095;
wire n_1096;
wire n_1097;
wire n_1098;
wire n_1099;
wire n_1100;
wire n_1101;
wire n_1102;
wire n_1103;
wire n_1104;
wire n_1105;
wire n_1106;
wire n_1107;
wire n_1108;
wire n_1109;
wire n_1110;
wire n_1111;
wire n_1112;
wire n_1113;
wire n_1114;
wire n_1115;
wire n_1116;
wire n_1117;
wire n_1118;
wire n_1119;
wire n_1120;
wire n_1121;
wire n_1122;
wire n_1123;
wire n_1124;
wire n_1125;
wire n_1126;
wire n_1127;
wire n_1128;
wire n_1129;
wire n_1130;
wire n_1131;
wire n_1132;
wire n_1133;
wire n_1134;
wire n_1135;
wire n_1136;
wire n_1137;
wire n_1138;
wire n_1139;
wire n_1140;
wire n_1141;
wire n_1142;
wire n_1143;
wire n_1144;
wire n_1145;
wire n_1146;
wire n_1147;
wire n_1148;
wire n_1149;
wire n_1150;
wire n_1151;
wire n_1152;
wire n_1153;
wire n_1154;
wire n_1155;
wire n_1156;
wire n_1157;
wire n_1158;
wire n_1159;
wire n_1160;
wire n_1161;
wire n_1162;
wire n_1163;
wire n_1164;
wire n_1165;
wire n_1166;
wire n_1167;
wire n_1168;
wire n_1169;
wire n_1170;
wire n_1171;
wire n_1172;
wire n_1173;
wire n_1174;
wire n_1175;
wire n_1176;
wire n_1177;
wire n_1178;
wire n_1179;
wire n_1180;
wire n_1181;
wire n_1182;
wire n_1183;
wire n_1184;
wire n_1185;
wire n_1186;
wire n_1187;
wire n_1188;
wire n_1189;
wire n_1190;
wire n_1191;
wire n_1192;
wire n_1193;
wire n_1194;
wire n_1195;
wire n_1196;
wire n_1197;
wire n_1198;
wire n_1199;
wire n_1200;
wire n_1201;
wire n_1202;
wire n_1203;
wire n_1204;
wire n_1205;
wire n_1206;
wire n_1207;
wire n_1208;
wire n_1209;
wire n_1210;
wire n_1211;
wire n_1212;
wire n_1213;
wire n_1214;
wire n_1215;
wire n_1216;
wire n_1217;
wire n_1218;
wire n_1219;
wire n_1220;
wire n_1221;
wire n_1222;
wire n_1223;
wire n_1224;
wire n_1225;
wire n_1226;
wire n_1227;
wire n_1228;
wire n_1229;
wire n_1230;
wire n_1231;
wire n_1232;
wire n_1233;
wire n_1234;
wire n_1235;
wire n_1236;
wire n_1237;
wire n_1238;
wire n_1239;
wire n_1240;
wire n_1241;
wire n_1242;
wire n_1243;
wire n_1244;
wire n_1245;
wire n_1246;
wire n_1247;
wire n_1248;
wire n_1249;
wire n_1250;
wire n_1251;
wire n_1252;
wire n_1253;
wire n_1254;
wire n_1255;
wire n_1256;
wire n_1257;
wire n_1258;
wire n_1259;
wire n_1260;
wire n_1261;
wire n_1262;
wire n_1263;
wire n_1264;
wire n_1265;
wire n_1266;
wire n_1267;
wire n_1268;
wire n_1269;
wire n_1270;
wire n_1271;
wire n_1272;
wire n_1273;
wire n_1274;
wire n_1275;
wire n_1276;
wire n_1277;
wire n_1278;
wire n_1279;
wire n_1280;
wire n_1281;
wire n_1282;
wire n_1283;
wire n_1284;
wire n_1285;
wire n_1286;
wire n_1287;
wire n_1288;
wire n_1289;
wire n_1290;
wire n_1291;
wire n_1292;
wire n_1293;
wire n_1294;
wire n_1295;
wire n_1296;
wire n_1297;
wire n_1298;
wire n_1299;
wire n_1300;
wire n_1301;
wire n_1302;
wire n_1303;
wire n_1304;
wire n_1305;
wire n_1306;
wire n_1307;
wire n_1308;
wire n_1309;
wire n_1310;
wire n_1311;
wire n_1312;
wire n_1313;
wire n_1314;
wire n_1315;
wire n_1316;
wire n_1317;
wire n_1318;
wire n_1319;
wire n_1320;
wire n_1321;
wire n_1322;
wire n_1323;
wire n_1324;
wire n_1325;
wire n_1326;
wire n_1327;
wire n_1328;
wire n_1329;
wire n_1330;
wire n_1331;
wire n_1332;
wire n_1333;
wire n_1334;
wire n_1335;
wire n_1336;
wire n_1337;
wire n_1338;
wire n_1339;
wire n_1340;
wire n_1341;
wire n_1342;
wire n_1343;
wire n_1344;
wire n_1345;
wire n_1346;
wire n_1347;
wire n_1348;
wire n_1349;
wire n_1350;
wire n_1351;
wire n_1352;
wire n_1353;
wire n_1354;
wire n_1355;
wire n_1356;
wire n_1357;
wire n_1358;
wire n_1359;
wire n_1360;
wire n_1361;
wire n_1362;
wire n_1363;
wire n_1364;
wire n_1365;
wire n_1366;
wire n_1367;
wire n_1368;
wire n_1369;
wire n_1370;
wire n_1371;
wire n_1372;
wire n_1373;
wire n_1374;
wire n_1375;
wire n_1376;
wire n_1377;
wire n_1378;
wire n_1379;
wire n_1380;
wire n_1381;
wire n_1382;
wire n_1383;
wire n_1384;
wire n_1385;
wire n_1386;
wire n_1387;
wire n_1388;
wire n_1389;
wire n_1390;
wire n_1391;
wire n_1392;
wire n_1393;
wire n_1394;
wire n_1395;
wire n_1396;
wire n_1397;
wire n_1398;
wire n_1399;
wire n_1400;
wire n_1401;
wire n_1402;
wire n_1403;
wire n_1404;
wire n_1405;
wire n_1406;
wire n_1407;
wire n_1408;
wire n_1409;
wire n_1410;
wire n_1411;
wire n_1412;
wire n_1413;
wire n_1414;
wire n_1415;
wire n_1416;
wire n_1417;
wire n_1418;
wire n_1419;
wire n_1420;
wire n_1421;
wire n_1422;
wire n_1423;
wire n_1424;
wire n_1425;
wire n_1426;
wire n_1427;
wire n_1428;
wire n_1429;
wire n_1430;
wire n_1431;
wire n_1432;
wire n_1433;
wire n_1434;
wire n_1435;
wire n_1436;
wire n_1437;
wire n_1438;
wire n_1439;
wire n_1440;
wire n_1441;
wire n_1442;
wire n_1443;
wire n_1444;
wire n_1445;
wire n_1446;
wire n_1447;
wire n_1448;
wire n_1449;
wire n_1450;
wire n_1451;
wire n_1452;
wire n_1453;
wire n_1454;
wire n_1455;
wire n_1456;
wire n_1457;
wire n_1458;
wire n_1459;
wire n_1460;
wire n_1461;
wire n_1462;
wire n_1463;
wire n_1464;
wire n_1465;
wire n_1466;
wire n_1467;
wire n_1468;
wire n_1469;
wire n_1470;
wire n_1471;
wire n_1472;
wire n_1473;
wire n_1474;
wire n_1475;
wire n_1476;
wire n_1477;
wire n_1478;
wire n_1479;
wire n_1480;
wire n_1481;
wire n_1482;
wire n_1483;
wire n_1484;
wire n_1485;
wire n_1486;
wire n_1487;
wire n_1488;
wire n_1489;
wire n_1490;
wire n_1491;
wire n_1492;
wire n_1493;
wire n_1494;
wire n_1495;
wire n_1496;
wire n_1497;
wire n_1498;
wire n_1499;
wire n_1500;
wire n_1501;
wire n_1502;
wire n_1503;
wire n_1504;
wire n_1505;
wire n_1506;
wire n_1507;
wire n_1508;
wire n_1509;
wire n_1510;
wire n_1511;
wire n_1512;
wire n_1513;
wire n_1514;
wire n_1515;
wire n_1516;
wire n_1517;
wire n_1518;
wire n_1519;
wire n_1520;
wire n_1521;
wire n_1522;
wire n_1523;
wire n_1524;
wire n_1525;
wire n_1526;
wire n_1527;
wire n_1528;
wire n_1529;
wire n_1530;
wire n_1531;
wire n_1532;
wire n_1533;
wire n_1534;
wire n_1535;
wire n_1536;
wire n_1537;
wire n_1538;
wire n_1539;
wire n_1540;
wire n_1541;
wire n_1542;
wire n_1543;
wire n_1544;
wire n_1545;
wire n_1546;
wire n_1547;
wire n_1548;
wire n_1549;
wire n_1550;
wire n_1551;
wire n_1552;
wire n_1553;
wire n_1554;
wire n_1555;
wire n_1556;
wire n_1557;
wire n_1558;
wire n_1559;
wire n_1560;
wire n_1561;
wire n_1562;
wire n_1563;
wire n_1564;
wire n_1565;
wire n_1566;
wire n_1567;
wire n_1568;
wire n_1569;
wire n_1570;
wire n_1571;
wire n_1572;
wire n_1573;
wire n_1574;
wire n_1575;
wire n_1576;
wire n_1577;
wire n_1578;
wire n_1579;
wire n_1580;
wire n_1581;
wire n_1582;
wire n_1583;
wire n_1584;
wire n_1585;
wire n_1586;
wire n_1587;
wire n_1588;
wire n_1589;
wire n_1590;
wire n_1591;
wire n_1592;
wire n_1593;
wire n_1594;
wire n_1595;
wire n_1596;
wire n_1597;
wire n_1598;
wire n_1599;
wire n_1600;
wire n_1601;
wire n_1602;
wire n_1603;
wire n_1604;
wire n_1605;
wire n_1606;
wire n_1607;
wire n_1608;
wire n_1609;
wire n_1610;
wire n_1611;
wire n_1612;
wire n_1613;
wire n_1614;
wire n_1615;
wire n_1616;
wire n_1617;
wire n_1618;
wire n_1619;
wire n_1620;
wire n_1621;
wire n_1622;
wire n_1623;
wire n_1624;
wire n_1625;
wire n_1626;
wire n_1627;
wire n_1628;
wire n_1629;
wire n_1630;
wire n_1631;
wire n_1632;
wire n_1633;
wire n_1634;
wire n_1635;
wire n_1636;
wire n_1637;
wire n_1638;
wire n_1639;
wire n_1640;
wire n_1641;
wire n_1642;
wire n_1643;
wire n_1644;
wire n_1645;
wire n_1646;
wire n_1647;
wire n_1648;
wire n_1649;
wire n_1650;
wire n_1651;
wire n_1652;
wire n_1653;
wire n_1654;
wire n_1655;
wire n_1656;
wire n_1657;
wire n_1658;
wire n_1659;
wire n_1660;
wire n_1661;
wire n_1662;
wire n_1663;
wire n_1664;
wire n_1665;
wire n_1666;
wire n_1667;
wire n_1668;
wire n_1669;
wire n_1670;
wire n_1671;
wire n_1672;
wire n_1673;
wire n_1674;
wire n_1675;
wire n_1676;
wire n_1677;
wire n_1678;
wire n_1679;
wire n_1680;
wire n_1681;
wire n_1682;
wire n_1683;
wire n_1684;
wire n_1685;
wire n_1686;
wire n_1687;
wire n_1688;
wire n_1689;
wire n_1690;
wire n_1691;
wire n_1692;
wire n_1693;
wire n_1694;
wire n_1695;
wire n_1696;
wire n_1697;
wire n_1698;
wire n_1699;
wire n_1700;
wire n_1701;
wire n_1702;
wire n_1703;
wire n_1704;
wire n_1705;
wire n_1706;
wire n_1707;
wire n_1708;
wire n_1709;
wire n_1710;
wire n_1711;
wire n_1712;
wire n_1713;
wire n_1714;
wire n_1715;
wire n_1716;
wire n_1717;
wire n_1718;
wire n_1719;
wire n_1720;
wire n_1721;
wire n_1722;
wire n_1723;
wire n_1724;
wire n_1725;
wire n_1726;
wire n_1727;
wire n_1728;
wire n_1729;
wire n_1730;
wire n_1731;
wire n_1732;
wire n_1733;
wire n_1734;
wire n_1735;
wire n_1736;
wire n_1737;
wire n_1738;
wire n_1739;
wire n_1740;
wire n_1741;
wire n_1742;
wire n_1743;
wire n_1744;
wire n_1745;
wire n_1746;
wire n_1747;
wire n_1748;
wire n_1749;
wire n_1750;
wire n_1751;
wire n_1752;
wire n_1753;
wire n_1754;
wire n_1755;
wire n_1756;
wire n_1757;
wire n_1758;
wire n_1759;
wire n_1760;
wire n_1761;
wire n_1762;
wire n_1763;
wire n_1764;
wire n_1765;
wire n_1766;
wire n_1767;
wire n_1768;
wire n_1769;
wire n_1770;
wire n_1771;
wire n_1772;
wire n_1773;
wire n_1774;
wire n_1775;
wire n_1776;
wire n_1777;
wire n_1778;
wire n_1779;
wire n_1780;
wire n_1781;
wire n_1782;
wire n_1783;
wire n_1784;
wire n_1785;
wire n_1786;
wire n_1787;
wire n_1788;
wire n_1789;
wire n_1790;
wire n_1791;
wire n_1792;
wire n_1793;
wire n_1794;
wire n_1795;
wire n_1796;
wire n_1797;
wire n_1798;
wire n_1799;
wire n_1800;
wire n_1801;
wire n_1802;
wire n_1803;
wire n_1804;
wire n_1805;
wire n_1806;
wire n_1807;
wire n_1808;
wire n_1809;
wire n_1810;
wire n_1811;
wire n_1812;
wire n_1813;
wire n_1814;
wire n_1815;
wire n_1816;
wire n_1817;
wire n_1818;
wire n_1819;
wire n_1820;
wire n_1821;
wire n_1822;
wire n_1823;
wire n_1824;
wire n_1825;
wire n_1826;
wire n_1827;
wire n_1828;
wire n_1829;
wire n_1830;
wire n_1831;
wire n_1832;
wire n_1833;
wire n_1834;
wire n_1835;
wire n_1836;
wire n_1837;
wire n_1838;
wire n_1839;
wire n_1840;
wire n_1841;
wire n_1842;
wire n_1843;
wire n_1844;
wire n_1845;
wire n_1846;
wire n_1847;
wire n_1848;
wire n_1849;
wire n_1850;
wire n_1851;
wire n_1852;
wire n_1853;
wire n_1854;
wire n_1855;
wire n_1856;
wire n_1857;
wire n_1858;
wire n_1859;
wire n_1860;
wire n_1861;
wire n_1862;
wire n_1863;
wire n_1864;
wire n_1865;
wire n_1866;
wire n_1867;
wire n_1868;
wire n_1869;
wire n_1870;
wire n_1871;
wire n_1872;
wire n_1873;
wire n_1874;
wire n_1875;
wire n_1876;
wire n_1877;
wire n_1878;
wire n_1879;
wire n_1880;
wire n_1881;
wire n_1882;
wire n_1883;
wire n_1884;
wire n_1885;
wire n_1886;
wire n_1887;
wire n_1888;
wire n_1889;
wire n_1890;
wire n_1891;
wire n_1892;
wire n_1893;
wire n_1894;
wire n_1895;
wire n_1896;
wire n_1897;
wire n_1898;
wire n_1899;
wire n_1900;
wire n_1901;
wire n_1902;
wire n_1903;
wire n_1904;
wire n_1905;
wire n_1906;
wire n_1907;
wire n_1908;
wire n_1909;
wire n_1910;
wire n_1911;
wire n_1912;
wire n_1913;
wire n_1914;
wire n_1915;
wire n_1916;
wire n_1917;
wire n_1918;
wire n_1919;
wire n_1920;
wire n_1921;
wire n_1922;
wire n_1923;
wire n_1924;
wire n_1925;
wire n_1926;
wire n_1927;
wire n_1928;
wire n_1929;
wire n_1930;
wire n_1931;
wire n_1932;
wire n_1933;
wire n_1934;
wire n_1935;
wire n_1936;
wire n_1937;
wire n_1938;
wire n_1939;
wire n_1940;
wire n_1941;
wire n_1942;
wire n_1943;
wire n_1944;
wire n_1945;
wire n_1946;
wire n_1947;
wire n_1948;
wire n_1949;
wire n_1950;
wire n_1951;
wire n_1952;
wire n_1953;
wire n_1954;
wire n_1955;
wire n_1956;
wire n_1957;
wire n_1958;
wire n_1959;
wire n_1960;
wire n_1961;
wire n_1962;
wire n_1963;
wire n_1964;
wire n_1965;
wire n_1966;
wire n_1967;
wire n_1968;
wire n_1969;
wire n_1970;
wire n_1971;
wire n_1972;
wire n_1973;
wire n_1974;
wire n_1975;
wire n_1976;
wire n_1977;
wire n_1978;
wire n_1979;
wire n_1980;
wire n_1981;
wire n_1982;
wire n_1983;
wire n_1984;
wire n_1985;
wire n_1986;
wire n_1987;
wire n_1988;
wire n_1989;
wire n_1990;
wire n_1991;
wire n_1992;
wire n_1993;
wire n_1994;
wire n_1995;
wire n_1996;
wire n_1997;
wire n_1998;
wire n_1999;
wire n_2000;
wire n_2001;
wire n_2002;
wire n_2003;
wire n_2004;
wire n_2005;
wire n_2006;
wire n_2007;
wire n_2008;
wire n_2009;
wire n_2010;
wire n_2011;
wire n_2012;
wire n_2013;
wire n_2014;
wire n_2015;
wire n_2016;
wire n_2017;
wire n_2018;
wire n_2019;
wire n_2020;
wire n_2021;
wire n_2022;
wire n_2023;
wire n_2024;
wire n_2025;
wire n_2026;
wire n_2027;
wire n_2028;
wire n_2029;
wire n_2030;
wire n_2031;
wire n_2032;
wire n_2033;
wire n_2034;
wire n_2035;
wire n_2036;
wire n_2037;
wire n_2038;
wire n_2039;
wire n_2040;
wire n_2041;
wire n_2042;
wire n_2043;
wire n_2044;
wire n_2045;
wire n_2046;
wire n_2047;
wire n_2048;
wire n_2049;
wire n_2050;
wire n_2051;
wire n_2052;
wire n_2053;
wire n_2054;
wire n_2055;
wire n_2056;
wire n_2057;
wire n_2058;
wire n_2059;
wire n_2060;
wire n_2061;
wire n_2062;
wire n_2063;
wire n_2064;
wire n_2065;
wire n_2066;
wire n_2067;
wire n_2068;
wire n_2069;
wire n_2070;
wire n_2071;
wire n_2072;
wire n_2073;
wire n_2074;
wire n_2075;
wire n_2076;
wire n_2077;
wire n_2078;
wire n_2079;
wire n_2080;
wire n_2081;
wire n_2082;
wire n_2083;
wire n_2084;
wire n_2085;
wire n_2086;
wire n_2087;
wire n_2088;
wire n_2089;
wire n_2090;
wire n_2091;
wire n_2092;
wire n_2093;
wire n_2094;
wire n_2095;
wire n_2096;
wire n_2097;
wire n_2098;
wire n_2099;
wire n_2100;
wire n_2101;
wire n_2102;
wire n_2103;
wire n_2104;
wire n_2105;
wire n_2106;
wire n_2107;
wire n_2108;
wire n_2109;
wire n_2110;
wire n_2111;
wire n_2112;
wire n_2113;
wire n_2114;
wire n_2115;
wire n_2116;
wire n_2117;
wire n_2118;
wire n_2119;
wire n_2120;
wire n_2121;
wire n_2122;
wire n_2123;
wire n_2124;
wire n_2125;
wire n_2126;
wire n_2127;
wire n_2128;
wire n_2129;
wire n_2130;
wire n_2131;
wire n_2132;
wire n_2133;
wire n_2134;
wire n_2135;
wire n_2136;
wire n_2137;
wire n_2138;
wire n_2139;
wire n_2140;
wire n_2141;
wire n_2142;
wire n_2143;
wire n_2144;
wire n_2145;
wire n_2146;
wire n_2147;
wire n_2148;
wire n_2149;
wire n_2150;
wire n_2151;
wire n_2152;
wire n_2153;
wire n_2154;
wire n_2155;
wire n_2156;
wire n_2157;
wire n_2158;
wire n_2159;
wire n_2160;
wire n_2161;
wire n_2162;
wire n_2163;
wire n_2164;
wire n_2165;
wire n_2166;
wire n_2167;
wire n_2168;
wire n_2169;
wire n_2170;
wire n_2171;
wire n_2172;
wire n_2173;
wire n_2174;
wire n_2175;
wire n_2176;
wire n_2177;
wire n_2178;
wire n_2179;
wire n_2180;
wire n_2181;
wire n_2182;
wire n_2183;
wire n_2184;
wire n_2185;
wire n_2186;
wire n_2187;
wire n_2188;
wire n_2189;
wire n_2190;
wire n_2191;
wire n_2192;
wire n_2193;
wire n_2194;
wire n_2195;
wire n_2196;
wire n_2197;
wire n_2198;
wire n_2199;
wire n_2200;
wire n_2201;
wire n_2202;
wire n_2203;
wire n_2204;
wire n_2205;
wire n_2206;
wire n_2207;
wire n_2208;
wire n_2209;
wire n_2210;
wire n_2211;
wire n_2212;
wire n_2213;
wire n_2214;
wire n_2215;
wire n_2216;
wire n_2217;
wire n_2218;
wire n_2219;
wire n_2220;
wire n_2221;
wire n_2222;
wire n_2223;
wire n_2224;
wire n_2225;
wire n_2226;
wire n_2227;
wire n_2228;
wire n_2229;
wire n_2230;
wire n_2231;
wire n_2232;
wire n_2233;
wire n_2234;
wire n_2235;
wire n_2236;
wire n_2237;
wire n_2238;
wire n_2239;
wire n_2240;
wire n_2241;
wire n_2242;
wire n_2243;
wire n_2244;
wire n_2245;
wire n_2246;
wire n_2247;
wire n_2248;
wire n_2249;
wire n_2250;
wire n_2251;
wire n_2252;
wire n_2253;
wire n_2254;
wire n_2255;
wire n_2256;
wire n_2257;
wire n_2258;
wire n_2259;
wire n_2260;
wire n_2261;
wire n_2262;
wire n_2263;
wire n_2264;
wire n_2265;
wire n_2266;
wire n_2267;
wire n_2268;
wire n_2269;
wire n_2270;
wire n_2271;
wire n_2272;
wire n_2273;
wire n_2274;
wire n_2275;
wire n_2276;
wire n_2277;
wire n_2278;
wire n_2279;
wire n_2280;
wire n_2281;
wire n_2282;
wire n_2283;
wire n_2284;
wire n_2285;
wire n_2286;
wire n_2287;
wire n_2288;
wire n_2289;
wire n_2290;
wire n_2291;
wire n_2292;
wire n_2293;
wire n_2294;
wire n_2295;
wire n_2296;
wire n_2297;
wire n_2298;
wire n_2299;
wire n_2300;
wire n_2301;
wire n_2302;
wire n_2303;
wire n_2304;
wire n_2305;
wire n_2306;
wire n_2307;
wire n_2308;
wire n_2309;
wire n_2310;
wire n_2311;
wire n_2312;
wire n_2313;
wire n_2314;
wire n_2315;
wire n_2316;
wire n_2317;
wire n_2318;
wire n_2319;
wire n_2320;
wire n_2321;
wire n_2322;
wire n_2323;
wire n_2324;
wire n_2325;
wire n_2326;
wire n_2327;
wire n_2328;
wire n_2329;
wire n_2330;
wire n_2331;
wire n_2332;
wire n_2333;
wire n_2334;
wire n_2335;
wire n_2336;
wire n_2337;
wire n_2338;
wire n_2339;
wire n_2340;
wire n_2341;
wire n_2342;
wire n_2343;
wire n_2344;
wire n_2345;
wire n_2346;
wire n_2347;
wire n_2348;
wire n_2349;
wire n_2350;
wire n_2351;
wire n_2352;
wire n_2353;
wire n_2354;
wire n_2355;
wire n_2356;
wire n_2357;
wire n_2358;
wire n_2359;
wire n_2360;
wire n_2361;
wire n_2362;
wire n_2363;
wire n_2364;
wire n_2365;
wire n_2366;
wire n_2367;
wire n_2368;
wire n_2369;
wire n_2370;
wire n_2371;
wire n_2372;
wire n_2373;
wire n_2374;
wire n_2375;
wire n_2376;
wire n_2377;
wire n_2378;
wire n_2379;
wire n_2380;
wire n_2381;
wire n_2382;
wire n_2383;
wire n_2384;
wire n_2385;
wire n_2386;
wire n_2387;
wire n_2388;
wire n_2389;
wire n_2390;
wire n_2391;
wire n_2392;
wire n_2393;
wire n_2394;
wire n_2395;
wire n_2396;
wire n_2397;
wire n_2398;
wire n_2399;
wire n_2400;
wire n_2401;
wire n_2402;
wire n_2403;
wire n_2404;
wire n_2405;
wire n_2406;
wire n_2407;
wire n_2408;
wire n_2409;
wire n_2410;
wire n_2411;
wire n_2412;
wire n_2413;
wire n_2414;
wire n_2415;
wire n_2416;
wire n_2417;
wire n_2418;
wire n_2419;
wire n_2420;
wire n_2421;
wire n_2422;
wire n_2423;
wire n_2424;
wire n_2425;
wire n_2426;
wire n_2427;
wire n_2428;
wire n_2429;
wire n_2430;
wire n_2431;
wire n_2432;
wire n_2433;
wire n_2434;
wire n_2435;
wire n_2436;
wire n_2437;
wire n_2438;
wire n_2439;
wire n_2440;
wire n_2441;
wire n_2442;
wire n_2443;
wire n_2444;
wire n_2445;
wire n_2446;
wire n_2447;
wire n_2448;
wire n_2449;
wire n_2450;
wire n_2451;
wire n_2452;
wire n_2453;
wire n_2454;
wire n_2455;
wire n_2456;
wire n_2457;
wire n_2458;
wire n_2459;
wire n_2460;
wire n_2461;
wire n_2462;
wire n_2463;
wire n_2464;
wire n_2465;
wire n_2466;
wire n_2467;
wire n_2468;
wire n_2469;
wire n_2470;
wire n_2471;
wire n_2472;
wire n_2473;
wire n_2474;
wire n_2475;
wire n_2476;
wire n_2477;
wire n_2478;
wire n_2479;
wire n_2480;
wire n_2481;
wire n_2482;
wire n_2483;
wire n_2484;
wire n_2485;
wire n_2486;
wire n_2487;
wire n_2488;
wire n_2489;
wire n_2490;
wire n_2491;
wire n_2492;
wire n_2493;
wire n_2494;
wire n_2495;
wire n_2496;
wire n_2497;
wire n_2498;
wire n_2499;
wire n_2500;
wire n_2501;
wire n_2502;
wire n_2503;
wire n_2504;
wire n_2505;
wire n_2506;
wire n_2507;
wire n_2508;
wire n_2509;
wire n_2510;
wire n_2511;
wire n_2512;
wire n_2513;
wire n_2514;
wire n_2515;
wire n_2516;
wire n_2517;
wire n_2518;
wire n_2519;
wire n_2520;
wire n_2521;
wire n_2522;
wire n_2523;
wire n_2524;
wire n_2525;
wire n_2526;
wire n_2527;
wire n_2528;
wire n_2529;
wire n_2530;
wire n_2531;
wire n_2532;
wire n_2533;
wire n_2534;
wire n_2535;
wire n_2536;
wire n_2537;
wire n_2538;
wire n_2539;
wire n_2540;
wire n_2541;
wire n_2542;
wire n_2543;
wire n_2544;
wire n_2545;
wire n_2546;
wire n_2547;
wire n_2548;
wire n_2549;
wire n_2550;
wire n_2551;
wire n_2552;
wire n_2553;
wire n_2554;
wire n_2555;
wire n_2556;
wire n_2557;
wire n_2558;
wire n_2559;
wire n_2560;
wire n_2561;
wire n_2562;
wire n_2563;
wire n_2564;
wire n_2565;
wire n_2566;
wire n_2567;
wire n_2568;
wire n_2569;
wire n_2570;
wire n_2571;
wire n_2572;
wire n_2573;
wire n_2574;
wire n_2575;
wire n_2576;
wire n_2577;
wire n_2578;
wire n_2579;
wire n_2580;
wire n_2581;
wire n_2582;
wire n_2583;
wire n_2584;
wire n_2585;
wire n_2586;
wire n_2587;
wire n_2588;
wire n_2589;
wire n_2590;
wire n_2591;
wire n_2592;
wire n_2593;
wire n_2594;
wire n_2595;
wire n_2596;
wire n_2597;
wire n_2598;
wire n_2599;
wire n_2600;
wire n_2601;
wire n_2602;
wire n_2603;
wire n_2604;
wire n_2605;
wire n_2606;
wire n_2607;
wire n_2608;
wire n_2609;
wire n_2610;
wire n_2611;
wire n_2612;
wire n_2613;
wire n_2614;
wire n_2615;
wire n_2616;
wire n_2617;
wire n_2618;
wire n_2619;
wire n_2620;
wire n_2621;
wire n_2622;
wire n_2623;
wire n_2624;
wire n_2625;
wire n_2626;
wire n_2627;
wire n_2628;
wire n_2629;
wire n_2630;
wire n_2631;
wire n_2632;
wire n_2633;
wire n_2634;
wire n_2635;
wire n_2636;
wire n_2637;
wire n_2638;
wire n_2639;
wire n_2640;
wire n_2641;
wire n_2642;
wire n_2643;
wire n_2644;
wire n_2645;
wire n_2646;
wire n_2647;
wire n_2648;
wire n_2649;
wire n_2650;
wire n_2651;
wire n_2652;
wire n_2653;
wire n_2654;
wire n_2655;
wire n_2656;
wire n_2657;
wire n_2658;
wire n_2659;
wire n_2660;
wire n_2661;
wire n_2662;
wire n_2663;
wire n_2664;
wire n_2665;
wire n_2666;
wire n_2667;
wire n_2668;
wire n_2669;
wire n_2670;
wire n_2671;
wire n_2672;
wire n_2673;
wire n_2674;
wire n_2675;
wire n_2676;
wire n_2677;
wire n_2678;
wire n_2679;
wire n_2680;
wire n_2681;
wire n_2682;
wire n_2683;
wire n_2684;
wire n_2685;
wire n_2686;
wire n_2687;
wire n_2688;
wire n_2689;
wire n_2690;
wire n_2691;
wire n_2692;
wire n_2693;
wire n_2694;
wire n_2695;
wire n_2696;
wire n_2697;
wire n_2698;
wire n_2699;
wire n_2700;
wire n_2701;
wire n_2702;
wire n_2703;
wire n_2704;
wire n_2705;
wire n_2706;
wire n_2707;
wire n_2708;
wire n_2709;
wire n_2710;
wire n_2711;
wire n_2712;
wire n_2713;
wire n_2714;
wire n_2715;
wire n_2716;
wire n_2717;
wire n_2718;
wire n_2719;
wire n_2720;
wire n_2721;
wire n_2722;
wire n_2723;
wire n_2724;
wire n_2725;
wire n_2726;
wire n_2727;
wire n_2728;
wire n_2729;
wire n_2730;
wire n_2731;
wire n_2732;
wire n_2733;
wire n_2734;
wire n_2735;
wire n_2736;
wire n_2737;
wire n_2738;
wire n_2739;
wire n_2740;
wire n_2741;
wire n_2742;
wire n_2743;
wire n_2744;
wire n_2745;
wire n_2746;
wire n_2747;
wire n_2748;
wire n_2749;
wire n_2750;
wire n_2751;
wire n_2752;
wire n_2753;
wire n_2754;
wire n_2755;
wire n_2756;
wire n_2757;
wire n_2758;
wire n_2759;
wire n_2760;
wire n_2761;
wire n_2762;
wire n_2763;
wire n_2764;
wire n_2765;
wire n_2766;
wire n_2767;
wire n_2768;
assign n_1 = ~x_305 & ~x_400;
assign n_2 = ~x_244 &  x_263;
assign n_3 =  x_270 & ~n_2;
assign n_4 =  n_1 & ~n_3;
assign n_5 = ~x_227 & ~n_4;
assign n_6 = ~x_283 & ~n_5;
assign n_7 = ~x_262 &  x_400;
assign n_8 = ~x_402 &  n_7;
assign n_9 =  x_311 & ~n_8;
assign n_10 =  x_364 & ~n_8;
assign n_11 = ~n_9 & ~n_10;
assign n_12 = ~n_6 &  n_11;
assign n_13 =  x_368 &  n_12;
assign n_14 = ~x_311 &  x_420;
assign n_15 = ~x_423 &  n_14;
assign n_16 =  x_421 &  n_15;
assign n_17 = ~x_311 &  x_424;
assign n_18 = ~x_422 &  n_17;
assign n_19 =  n_16 &  n_18;
assign n_20 = ~x_420 & ~x_421;
assign n_21 = ~x_311 &  x_423;
assign n_22 =  n_20 &  n_21;
assign n_23 = ~x_423 &  n_20;
assign n_24 = ~n_22 & ~n_23;
assign n_25 = ~n_16 &  n_24;
assign n_26 = ~x_424 & ~n_25;
assign n_27 = ~x_421 &  n_15;
assign n_28 =  x_421 & ~n_14;
assign n_29 = ~n_21 &  n_28;
assign n_30 = ~n_27 & ~n_29;
assign n_31 = ~n_26 &  n_30;
assign n_32 =  x_422 & ~n_31;
assign n_33 = ~x_420 &  x_423;
assign n_34 =  x_420 &  x_421;
assign n_35 = ~n_20 & ~n_34;
assign n_36 =  x_422 & ~n_35;
assign n_37 = ~n_33 & ~n_36;
assign n_38 =  x_424 & ~n_37;
assign n_39 = ~x_421 & ~x_424;
assign n_40 =  x_420 &  x_422;
assign n_41 = ~n_39 &  n_40;
assign n_42 =  x_423 & ~n_20;
assign n_43 = ~n_41 &  n_42;
assign n_44 = ~n_38 & ~n_43;
assign n_45 = ~n_32 &  n_44;
assign n_46 = ~x_311 & ~n_45;
assign n_47 = ~n_6 & ~n_11;
assign n_48 = ~x_311 &  x_422;
assign n_49 = ~n_48 & ~n_17;
assign n_50 =  n_49 &  n_22;
assign n_51 =  n_47 & ~n_50;
assign n_52 = ~n_46 &  n_51;
assign n_53 = ~n_19 &  n_52;
assign n_54 =  n_49 &  n_16;
assign n_55 =  n_53 & ~n_54;
assign n_56 =  n_27 &  n_18;
assign n_57 =  n_55 &  n_56;
assign n_58 = ~n_13 & ~n_57;
assign n_59 =  x_368 & ~n_58;
assign n_60 = ~x_368 &  n_58;
assign n_61 = ~n_59 & ~n_60;
assign n_62 =  x_367 &  n_12;
assign n_63 =  n_53 &  n_54;
assign n_64 = ~n_62 & ~n_63;
assign n_65 =  x_367 & ~n_64;
assign n_66 = ~x_367 &  n_64;
assign n_67 = ~n_65 & ~n_66;
assign n_68 =  x_366 &  n_12;
assign n_69 = ~i_205 & ~x_425;
assign n_70 =  i_204 &  i_206;
assign n_71 = ~n_69 &  n_70;
assign n_72 =  i_207 & ~n_71;
assign n_73 =  i_206 & ~i_207;
assign n_74 =  i_204 &  i_205;
assign n_75 =  x_425 &  n_74;
assign n_76 = ~n_73 & ~n_75;
assign n_77 = ~n_72 &  n_76;
assign n_78 = ~x_311 & ~n_77;
assign n_79 =  n_47 & ~n_78;
assign n_80 = ~i_207 & ~x_311;
assign n_81 =  i_204 &  n_80;
assign n_82 =  i_206 & ~x_311;
assign n_83 = ~x_311 &  x_425;
assign n_84 = ~n_82 & ~n_83;
assign n_85 =  i_205 &  n_84;
assign n_86 =  n_81 &  n_85;
assign n_87 =  n_79 &  n_86;
assign n_88 = ~n_68 & ~n_87;
assign n_89 =  x_366 & ~n_88;
assign n_90 = ~x_366 &  n_88;
assign n_91 = ~n_89 & ~n_90;
assign n_92 =  x_310 &  x_324;
assign n_93 =  i_3 & ~x_325;
assign n_94 = ~n_5 &  n_93;
assign n_95 =  x_245 & ~x_327;
assign n_96 =  x_261 &  n_95;
assign n_97 =  x_271 & ~n_96;
assign n_98 =  x_416 & ~n_95;
assign n_99 =  n_97 & ~n_98;
assign n_100 = ~i_172 & ~n_95;
assign n_101 = ~x_227 & ~n_100;
assign n_102 = ~x_326 & ~x_341;
assign n_103 = ~x_249 & ~x_417;
assign n_104 =  n_102 &  n_103;
assign n_105 = ~x_270 & ~x_418;
assign n_106 =  n_104 &  n_105;
assign n_107 =  x_272 &  n_106;
assign n_108 = ~n_101 &  n_107;
assign n_109 = ~n_99 & ~n_108;
assign n_110 =  n_94 & ~n_109;
assign n_111 =  n_92 &  n_110;
assign n_112 = ~x_263 &  x_270;
assign n_113 =  x_365 & ~n_112;
assign n_114 =  n_5 &  n_113;
assign n_115 = ~n_111 & ~n_114;
assign n_116 =  x_365 & ~n_115;
assign n_117 = ~x_365 &  n_115;
assign n_118 = ~n_116 & ~n_117;
assign n_119 = ~x_228 & ~x_232;
assign n_120 =  i_146 &  x_424;
assign n_121 = ~i_199 &  x_420;
assign n_122 = ~i_146 & ~x_424;
assign n_123 = ~n_121 & ~n_122;
assign n_124 = ~n_120 &  n_123;
assign n_125 = ~i_200 & ~x_421;
assign n_126 =  i_200 &  x_421;
assign n_127 = ~n_125 & ~n_126;
assign n_128 =  i_199 & ~x_420;
assign n_129 =  i_147 & ~x_422;
assign n_130 = ~n_128 &  n_129;
assign n_131 = ~i_198 &  x_423;
assign n_132 =  i_198 & ~x_423;
assign n_133 = ~n_131 & ~n_132;
assign n_134 =  n_130 &  n_133;
assign n_135 = ~n_127 &  n_134;
assign n_136 =  n_124 &  n_135;
assign n_137 = ~i_49 &  i_144;
assign n_138 = ~i_47 &  i_142;
assign n_139 = ~n_137 & ~n_138;
assign n_140 =  i_48 & ~i_143;
assign n_141 =  i_50 & ~i_145;
assign n_142 = ~n_140 & ~n_141;
assign n_143 =  n_139 &  n_142;
assign n_144 = ~i_48 &  i_143;
assign n_145 =  i_49 & ~i_144;
assign n_146 = ~n_144 & ~n_145;
assign n_147 = ~i_50 &  i_145;
assign n_148 =  i_47 & ~i_142;
assign n_149 = ~n_147 & ~n_148;
assign n_150 =  n_146 &  n_149;
assign n_151 =  n_143 &  n_150;
assign n_152 = ~i_46 &  n_151;
assign n_153 = ~i_202 &  x_420;
assign n_154 = ~i_139 & ~x_424;
assign n_155 =  i_202 & ~x_420;
assign n_156 = ~n_154 & ~n_155;
assign n_157 = ~n_153 &  n_156;
assign n_158 = ~i_201 & ~x_423;
assign n_159 =  i_201 &  x_423;
assign n_160 = ~n_158 & ~n_159;
assign n_161 = ~i_203 & ~x_421;
assign n_162 =  i_203 &  x_421;
assign n_163 = ~n_161 & ~n_162;
assign n_164 =  i_139 &  x_424;
assign n_165 =  i_140 & ~x_422;
assign n_166 = ~n_164 &  n_165;
assign n_167 = ~n_163 &  n_166;
assign n_168 = ~n_160 &  n_167;
assign n_169 =  n_157 &  n_168;
assign n_170 = ~n_152 & ~n_169;
assign n_171 = ~n_136 &  n_170;
assign n_172 = ~i_201 &  i_207;
assign n_173 =  i_139 &  x_425;
assign n_174 =  i_201 & ~i_207;
assign n_175 = ~n_173 & ~n_174;
assign n_176 = ~n_172 &  n_175;
assign n_177 = ~i_203 & ~i_205;
assign n_178 =  i_203 &  i_205;
assign n_179 = ~n_177 & ~n_178;
assign n_180 = ~i_139 & ~x_425;
assign n_181 =  i_140 & ~i_206;
assign n_182 = ~n_180 &  n_181;
assign n_183 =  i_202 & ~i_204;
assign n_184 = ~i_202 &  i_204;
assign n_185 = ~n_183 & ~n_184;
assign n_186 =  n_182 &  n_185;
assign n_187 = ~n_179 &  n_186;
assign n_188 =  n_176 &  n_187;
assign n_189 = ~i_46 & ~i_141;
assign n_190 =  i_46 &  i_141;
assign n_191 = ~n_189 & ~n_190;
assign n_192 =  n_151 & ~n_191;
assign n_193 = ~i_199 &  i_204;
assign n_194 = ~i_146 & ~x_425;
assign n_195 =  i_199 & ~i_204;
assign n_196 = ~n_194 & ~n_195;
assign n_197 = ~n_193 &  n_196;
assign n_198 = ~i_198 & ~i_207;
assign n_199 =  i_198 &  i_207;
assign n_200 = ~n_198 & ~n_199;
assign n_201 = ~i_200 & ~i_205;
assign n_202 =  i_200 &  i_205;
assign n_203 = ~n_201 & ~n_202;
assign n_204 =  i_146 &  x_425;
assign n_205 =  i_147 & ~i_206;
assign n_206 = ~n_204 &  n_205;
assign n_207 = ~n_203 &  n_206;
assign n_208 = ~n_200 &  n_207;
assign n_209 =  n_197 &  n_208;
assign n_210 = ~n_192 & ~n_209;
assign n_211 = ~n_188 &  n_210;
assign n_212 =  n_171 &  n_211;
assign n_213 = ~x_283 & ~x_312;
assign n_214 = ~x_304 & ~x_311;
assign n_215 = ~n_213 &  n_214;
assign n_216 = ~n_212 &  n_215;
assign n_217 = ~x_419 & ~n_216;
assign n_218 = ~x_313 & ~x_314;
assign n_219 =  x_419 &  n_218;
assign n_220 = ~n_8 & ~n_219;
assign n_221 = ~n_217 &  n_220;
assign n_222 =  x_364 & ~n_221;
assign n_223 =  x_304 & ~n_8;
assign n_224 =  i_165 &  x_307;
assign n_225 = ~n_223 & ~n_224;
assign n_226 = ~n_222 &  n_225;
assign n_227 =  n_119 & ~n_226;
assign n_228 =  x_364 &  n_227;
assign n_229 = ~x_364 & ~n_227;
assign n_230 = ~n_228 & ~n_229;
assign n_231 =  x_363 &  n_12;
assign n_232 =  n_49 &  n_27;
assign n_233 =  n_55 & ~n_56;
assign n_234 =  n_232 &  n_233;
assign n_235 = ~n_231 & ~n_234;
assign n_236 =  x_363 & ~n_235;
assign n_237 = ~x_363 &  n_235;
assign n_238 = ~n_236 & ~n_237;
assign n_239 = ~x_228 & ~n_6;
assign n_240 = ~n_9 & ~n_112;
assign n_241 =  x_362 &  n_240;
assign n_242 =  n_239 &  n_241;
assign n_243 = ~n_10 & ~n_242;
assign n_244 =  x_362 & ~n_243;
assign n_245 = ~x_362 &  n_243;
assign n_246 = ~n_244 & ~n_245;
assign n_247 =  x_361 &  n_12;
assign n_248 = ~i_205 &  n_81;
assign n_249 =  n_84 &  n_248;
assign n_250 = ~i_206 &  n_83;
assign n_251 =  n_248 &  n_250;
assign n_252 =  n_79 & ~n_251;
assign n_253 =  n_249 &  n_252;
assign n_254 = ~n_247 & ~n_253;
assign n_255 =  x_361 & ~n_254;
assign n_256 = ~x_361 &  n_254;
assign n_257 = ~n_255 & ~n_256;
assign n_258 = ~x_311 &  x_312;
assign n_259 = ~n_171 &  n_258;
assign n_260 =  x_314 &  x_419;
assign n_261 = ~n_260 &  n_10;
assign n_262 = ~n_259 &  n_261;
assign n_263 =  i_171 &  n_8;
assign n_264 =  x_360 & ~n_10;
assign n_265 = ~n_263 &  n_264;
assign n_266 =  n_240 &  n_265;
assign n_267 =  n_239 &  n_266;
assign n_268 = ~n_262 & ~n_267;
assign n_269 =  x_360 & ~n_268;
assign n_270 = ~x_360 &  n_268;
assign n_271 = ~n_269 & ~n_270;
assign n_272 =  x_365 &  n_9;
assign n_273 =  x_359 &  n_240;
assign n_274 = ~n_272 & ~n_273;
assign n_275 =  n_5 & ~n_274;
assign n_276 = ~n_92 &  n_110;
assign n_277 = ~n_275 & ~n_276;
assign n_278 = ~x_228 & ~n_277;
assign n_279 =  x_359 &  n_278;
assign n_280 = ~x_359 & ~n_278;
assign n_281 = ~n_279 & ~n_280;
assign n_282 =  x_358 &  n_8;
assign n_283 = ~x_228 & ~n_8;
assign n_284 =  x_362 &  x_363;
assign n_285 =  x_360 &  x_361;
assign n_286 =  i_170 &  x_359;
assign n_287 = ~n_285 & ~n_286;
assign n_288 = ~n_284 &  n_287;
assign n_289 = ~n_3 & ~n_288;
assign n_290 =  n_283 &  n_289;
assign n_291 = ~n_282 & ~n_290;
assign n_292 =  x_358 & ~n_291;
assign n_293 = ~x_358 &  n_291;
assign n_294 = ~n_292 & ~n_293;
assign n_295 =  x_357 &  n_8;
assign n_296 =  x_362 &  x_367;
assign n_297 =  x_360 &  x_366;
assign n_298 =  i_173 &  x_359;
assign n_299 = ~n_297 & ~n_298;
assign n_300 = ~n_296 &  n_299;
assign n_301 = ~n_3 & ~n_300;
assign n_302 =  n_283 &  n_301;
assign n_303 = ~n_295 & ~n_302;
assign n_304 =  x_357 & ~n_303;
assign n_305 = ~x_357 &  n_303;
assign n_306 = ~n_304 & ~n_305;
assign n_307 =  x_356 &  n_8;
assign n_308 =  x_362 &  x_368;
assign n_309 =  i_175 &  x_360;
assign n_310 =  i_174 &  x_359;
assign n_311 = ~n_309 & ~n_310;
assign n_312 = ~n_308 &  n_311;
assign n_313 = ~n_3 & ~n_312;
assign n_314 =  n_283 &  n_313;
assign n_315 = ~n_307 & ~n_314;
assign n_316 =  x_356 & ~n_315;
assign n_317 = ~x_356 &  n_315;
assign n_318 = ~n_316 & ~n_317;
assign n_319 =  x_355 &  n_8;
assign n_320 =  x_362 &  x_370;
assign n_321 =  x_360 &  x_369;
assign n_322 =  i_176 &  x_359;
assign n_323 = ~n_321 & ~n_322;
assign n_324 = ~n_320 &  n_323;
assign n_325 = ~n_3 & ~n_324;
assign n_326 =  n_283 &  n_325;
assign n_327 = ~n_319 & ~n_326;
assign n_328 =  x_355 & ~n_327;
assign n_329 = ~x_355 &  n_327;
assign n_330 = ~n_328 & ~n_329;
assign n_331 =  x_354 &  n_8;
assign n_332 =  x_362 &  x_371;
assign n_333 =  i_178 &  x_360;
assign n_334 =  i_177 &  x_359;
assign n_335 = ~n_333 & ~n_334;
assign n_336 = ~n_332 &  n_335;
assign n_337 = ~n_3 & ~n_336;
assign n_338 =  n_283 &  n_337;
assign n_339 = ~n_331 & ~n_338;
assign n_340 =  x_354 & ~n_339;
assign n_341 = ~x_354 &  n_339;
assign n_342 = ~n_340 & ~n_341;
assign n_343 =  x_353 &  n_8;
assign n_344 =  x_362 &  x_374;
assign n_345 =  x_360 &  x_373;
assign n_346 =  x_359 &  x_372;
assign n_347 = ~n_345 & ~n_346;
assign n_348 = ~n_344 &  n_347;
assign n_349 = ~n_3 & ~n_348;
assign n_350 =  n_283 &  n_349;
assign n_351 = ~n_343 & ~n_350;
assign n_352 =  x_353 & ~n_351;
assign n_353 = ~x_353 &  n_351;
assign n_354 = ~n_352 & ~n_353;
assign n_355 =  x_352 &  n_8;
assign n_356 =  x_362 &  x_377;
assign n_357 =  x_360 &  x_376;
assign n_358 =  x_359 &  x_375;
assign n_359 = ~n_357 & ~n_358;
assign n_360 = ~n_356 &  n_359;
assign n_361 = ~n_3 & ~n_360;
assign n_362 =  n_283 &  n_361;
assign n_363 = ~n_355 & ~n_362;
assign n_364 =  x_352 & ~n_363;
assign n_365 = ~x_352 &  n_363;
assign n_366 = ~n_364 & ~n_365;
assign n_367 =  x_351 &  n_8;
assign n_368 =  x_214 & ~x_379;
assign n_369 =  x_362 & ~n_368;
assign n_370 = ~i_179 &  x_214;
assign n_371 =  x_360 & ~n_370;
assign n_372 =  x_214 & ~x_378;
assign n_373 =  x_359 & ~n_372;
assign n_374 = ~n_371 & ~n_373;
assign n_375 = ~n_369 &  n_374;
assign n_376 = ~n_3 & ~n_375;
assign n_377 =  n_376 &  n_283;
assign n_378 = ~n_367 & ~n_377;
assign n_379 =  x_351 & ~n_378;
assign n_380 = ~x_351 &  n_378;
assign n_381 = ~n_379 & ~n_380;
assign n_382 =  x_351 &  n_283;
assign n_383 = ~n_376 &  n_382;
assign n_384 =  x_350 &  n_383;
assign n_385 = ~x_350 & ~n_383;
assign n_386 = ~n_384 & ~n_385;
assign n_387 =  x_349 &  n_5;
assign n_388 =  x_272 &  n_98;
assign n_389 = ~n_99 & ~n_388;
assign n_390 = ~n_389 &  n_94;
assign n_391 = ~n_387 & ~n_390;
assign n_392 =  x_349 & ~n_391;
assign n_393 = ~x_349 &  n_391;
assign n_394 = ~n_392 & ~n_393;
assign n_395 = ~i_156 &  x_308;
assign n_396 = ~x_308 &  x_348;
assign n_397 = ~n_395 & ~n_396;
assign n_398 =  x_348 & ~n_397;
assign n_399 = ~x_348 &  n_397;
assign n_400 = ~n_398 & ~n_399;
assign n_401 =  i_163 &  x_308;
assign n_402 = ~x_308 &  x_347;
assign n_403 = ~n_401 & ~n_402;
assign n_404 =  x_347 & ~n_403;
assign n_405 = ~x_347 &  n_403;
assign n_406 = ~n_404 & ~n_405;
assign n_407 =  i_160 &  x_308;
assign n_408 = ~x_308 &  x_346;
assign n_409 = ~n_407 & ~n_408;
assign n_410 =  x_346 & ~n_409;
assign n_411 = ~x_346 &  n_409;
assign n_412 = ~n_410 & ~n_411;
assign n_413 =  i_158 &  x_308;
assign n_414 = ~x_308 &  x_345;
assign n_415 = ~n_413 & ~n_414;
assign n_416 =  x_345 & ~n_415;
assign n_417 = ~x_345 &  n_415;
assign n_418 = ~n_416 & ~n_417;
assign n_419 = ~x_308 & ~x_344;
assign n_420 = ~n_395 & ~n_419;
assign n_421 =  x_344 &  n_420;
assign n_422 = ~x_344 & ~n_420;
assign n_423 = ~n_421 & ~n_422;
assign n_424 = ~i_7 & ~x_231;
assign n_425 =  x_343 &  n_424;
assign n_426 = ~x_228 & ~n_425;
assign n_427 =  x_343 & ~n_426;
assign n_428 = ~x_343 &  n_426;
assign n_429 = ~n_427 & ~n_428;
assign n_430 =  x_335 &  x_342;
assign n_431 = ~x_335 & ~x_342;
assign n_432 = ~n_430 & ~n_431;
assign n_433 = ~x_228 &  x_249;
assign n_434 =  x_341 &  n_433;
assign n_435 = ~x_341 & ~n_433;
assign n_436 = ~n_434 & ~n_435;
assign n_437 = ~x_303 & ~x_400;
assign n_438 = ~x_402 &  n_437;
assign n_439 =  x_268 &  x_269;
assign n_440 =  n_438 &  n_439;
assign n_441 =  i_2 &  n_440;
assign n_442 = ~x_243 & ~x_259;
assign n_443 = ~x_339 &  n_442;
assign n_444 = ~i_153 & ~x_229;
assign n_445 = ~x_230 & ~x_231;
assign n_446 =  n_444 &  n_445;
assign n_447 =  n_119 &  n_446;
assign n_448 =  n_443 &  n_447;
assign n_449 =  n_441 &  n_448;
assign n_450 =  x_340 &  n_449;
assign n_451 = ~x_340 & ~n_449;
assign n_452 = ~n_450 & ~n_451;
assign n_453 =  i_7 &  x_343;
assign n_454 =  x_338 & ~n_453;
assign n_455 = ~x_260 & ~n_454;
assign n_456 =  i_8 & ~x_337;
assign n_457 = ~n_453 &  n_456;
assign n_458 =  n_443 &  n_457;
assign n_459 = ~n_455 &  n_458;
assign n_460 =  x_339 &  n_459;
assign n_461 = ~x_339 & ~n_459;
assign n_462 = ~n_460 & ~n_461;
assign n_463 =  x_338 & ~n_455;
assign n_464 = ~x_338 &  n_455;
assign n_465 = ~n_463 & ~n_464;
assign n_466 =  x_337 &  n_453;
assign n_467 = ~x_337 & ~n_453;
assign n_468 = ~n_466 & ~n_467;
assign n_469 =  x_332 &  x_333;
assign n_470 =  x_334 &  n_469;
assign n_471 = ~x_334 & ~n_469;
assign n_472 = ~n_470 & ~n_471;
assign n_473 =  i_150 & ~n_472;
assign n_474 = ~i_150 &  n_472;
assign n_475 =  i_149 &  i_213;
assign n_476 = ~i_149 & ~i_213;
assign n_477 = ~x_332 & ~x_333;
assign n_478 = ~n_469 & ~n_477;
assign n_479 = ~n_476 & ~n_478;
assign n_480 = ~n_475 & ~n_479;
assign n_481 = ~n_474 & ~n_480;
assign n_482 = ~n_473 & ~n_481;
assign n_483 =  i_151 & ~n_482;
assign n_484 = ~i_151 &  n_482;
assign n_485 = ~n_483 & ~n_484;
assign n_486 =  i_152 & ~n_470;
assign n_487 = ~i_152 &  n_470;
assign n_488 = ~n_486 & ~n_487;
assign n_489 = ~n_485 & ~n_488;
assign n_490 =  n_485 &  n_488;
assign n_491 =  i_4 & ~n_490;
assign n_492 = ~n_489 &  n_491;
assign n_493 =  i_6 &  n_492;
assign n_494 = ~x_225 & ~x_242;
assign n_495 = ~x_257 & ~x_336;
assign n_496 =  n_494 &  n_495;
assign n_497 =  n_493 &  n_496;
assign n_498 =  x_336 &  n_497;
assign n_499 = ~x_336 & ~n_497;
assign n_500 = ~n_498 & ~n_499;
assign n_501 =  x_335 &  n_493;
assign n_502 = ~x_335 & ~n_493;
assign n_503 = ~n_501 & ~n_502;
assign n_504 = ~i_16 &  n_492;
assign n_505 = ~i_17 &  n_504;
assign n_506 = ~x_329 & ~x_330;
assign n_507 = ~x_331 &  n_506;
assign n_508 =  x_215 &  n_507;
assign n_509 =  n_505 & ~n_508;
assign n_510 = ~n_472 &  n_509;
assign n_511 =  i_16 &  n_492;
assign n_512 = ~i_17 &  n_511;
assign n_513 = ~x_334 & ~n_509;
assign n_514 = ~n_512 & ~n_513;
assign n_515 = ~n_510 &  n_514;
assign n_516 =  i_17 &  n_504;
assign n_517 = ~x_215 &  x_330;
assign n_518 =  x_329 &  x_330;
assign n_519 = ~x_331 & ~n_518;
assign n_520 = ~n_517 &  n_519;
assign n_521 = ~x_334 &  n_520;
assign n_522 = ~n_472 & ~n_520;
assign n_523 = ~n_521 & ~n_522;
assign n_524 =  n_512 &  n_523;
assign n_525 = ~n_516 & ~n_524;
assign n_526 = ~n_515 &  n_525;
assign n_527 =  i_17 &  n_511;
assign n_528 =  x_331 & ~n_506;
assign n_529 = ~n_472 &  n_528;
assign n_530 = ~x_334 & ~n_528;
assign n_531 =  x_215 & ~n_530;
assign n_532 = ~n_529 &  n_531;
assign n_533 =  x_331 &  n_469;
assign n_534 =  x_334 &  n_533;
assign n_535 = ~x_334 & ~n_533;
assign n_536 = ~x_215 & ~n_535;
assign n_537 = ~n_534 &  n_536;
assign n_538 = ~n_532 & ~n_537;
assign n_539 =  n_516 &  n_538;
assign n_540 = ~n_527 & ~n_539;
assign n_541 = ~n_526 &  n_540;
assign n_542 =  x_215 &  n_527;
assign n_543 =  x_331 &  n_518;
assign n_544 = ~x_334 & ~n_543;
assign n_545 =  n_542 & ~n_544;
assign n_546 = ~x_215 &  n_527;
assign n_547 =  x_330 &  x_331;
assign n_548 = ~x_334 & ~n_547;
assign n_549 =  n_546 & ~n_548;
assign n_550 = ~n_545 & ~n_549;
assign n_551 = ~x_329 &  n_545;
assign n_552 = ~n_472 &  n_547;
assign n_553 = ~n_551 &  n_552;
assign n_554 = ~n_550 & ~n_553;
assign n_555 = ~n_541 & ~n_554;
assign n_556 = ~x_225 & ~n_555;
assign n_557 =  i_21 &  x_225;
assign n_558 = ~n_556 & ~n_557;
assign n_559 =  x_334 & ~n_558;
assign n_560 = ~x_334 &  n_558;
assign n_561 = ~n_559 & ~n_560;
assign n_562 = ~i_22 &  x_225;
assign n_563 =  n_478 &  n_509;
assign n_564 =  x_333 & ~n_509;
assign n_565 = ~n_512 & ~n_564;
assign n_566 = ~n_563 &  n_565;
assign n_567 = ~x_330 & ~x_331;
assign n_568 =  x_332 & ~n_567;
assign n_569 = ~x_215 & ~n_568;
assign n_570 =  x_332 & ~n_519;
assign n_571 =  x_215 & ~n_570;
assign n_572 = ~n_569 & ~n_571;
assign n_573 =  x_333 & ~n_572;
assign n_574 = ~x_333 &  n_572;
assign n_575 = ~n_573 & ~n_574;
assign n_576 =  n_512 &  n_575;
assign n_577 = ~n_566 & ~n_576;
assign n_578 = ~n_516 & ~n_577;
assign n_579 =  x_331 &  x_332;
assign n_580 = ~x_333 & ~n_579;
assign n_581 = ~n_580 & ~n_533;
assign n_582 = ~x_215 & ~n_581;
assign n_583 =  x_333 & ~n_528;
assign n_584 =  n_478 &  n_528;
assign n_585 =  x_215 & ~n_584;
assign n_586 = ~n_583 &  n_585;
assign n_587 = ~n_582 & ~n_586;
assign n_588 =  n_516 & ~n_587;
assign n_589 = ~n_546 & ~n_588;
assign n_590 = ~n_578 &  n_589;
assign n_591 = ~x_333 & ~n_547;
assign n_592 = ~n_478 &  n_547;
assign n_593 = ~n_591 & ~n_592;
assign n_594 =  n_527 &  n_593;
assign n_595 = ~n_590 & ~n_594;
assign n_596 = ~n_542 & ~n_595;
assign n_597 = ~x_333 & ~n_543;
assign n_598 = ~n_478 &  n_543;
assign n_599 = ~n_597 & ~n_598;
assign n_600 =  n_542 &  n_599;
assign n_601 = ~x_225 & ~n_600;
assign n_602 = ~n_596 &  n_601;
assign n_603 = ~n_562 & ~n_602;
assign n_604 =  x_333 &  n_603;
assign n_605 = ~x_333 & ~n_603;
assign n_606 = ~n_604 & ~n_605;
assign n_607 = ~i_23 &  x_225;
assign n_608 = ~x_332 & ~n_547;
assign n_609 =  x_330 &  n_579;
assign n_610 = ~x_215 & ~n_609;
assign n_611 = ~n_608 &  n_610;
assign n_612 =  n_527 & ~n_611;
assign n_613 = ~x_331 & ~x_332;
assign n_614 = ~x_215 & ~n_579;
assign n_615 = ~n_613 &  n_614;
assign n_616 =  n_516 & ~n_615;
assign n_617 =  x_332 &  n_509;
assign n_618 = ~x_332 & ~n_509;
assign n_619 = ~n_512 & ~n_618;
assign n_620 = ~n_617 &  n_619;
assign n_621 =  x_215 &  n_512;
assign n_622 = ~n_518 &  n_613;
assign n_623 = ~n_570 & ~n_622;
assign n_624 =  n_621 &  n_623;
assign n_625 = ~x_215 &  n_516;
assign n_626 = ~x_332 &  n_567;
assign n_627 =  n_569 & ~n_626;
assign n_628 =  n_512 &  n_627;
assign n_629 = ~n_625 & ~n_628;
assign n_630 = ~n_624 &  n_629;
assign n_631 = ~n_620 &  n_630;
assign n_632 = ~n_616 & ~n_631;
assign n_633 =  x_215 &  n_516;
assign n_634 = ~x_332 & ~n_528;
assign n_635 =  x_332 &  n_528;
assign n_636 = ~n_634 & ~n_635;
assign n_637 =  n_633 &  n_636;
assign n_638 = ~n_546 & ~n_637;
assign n_639 = ~n_632 &  n_638;
assign n_640 = ~n_612 & ~n_639;
assign n_641 = ~x_332 & ~n_543;
assign n_642 =  x_329 &  n_609;
assign n_643 = ~n_641 & ~n_642;
assign n_644 =  n_542 &  n_643;
assign n_645 = ~x_225 & ~n_644;
assign n_646 = ~n_640 &  n_645;
assign n_647 = ~n_607 & ~n_646;
assign n_648 =  x_332 &  n_647;
assign n_649 = ~x_332 & ~n_647;
assign n_650 = ~n_648 & ~n_649;
assign n_651 =  i_24 &  x_225;
assign n_652 = ~n_547 & ~n_567;
assign n_653 = ~x_215 & ~n_652;
assign n_654 =  n_527 & ~n_653;
assign n_655 = ~x_215 &  x_331;
assign n_656 =  n_516 & ~n_655;
assign n_657 = ~x_215 &  n_512;
assign n_658 =  x_215 &  n_505;
assign n_659 =  x_331 & ~n_658;
assign n_660 = ~n_657 &  n_659;
assign n_661 = ~n_528 & ~n_507;
assign n_662 =  n_658 & ~n_661;
assign n_663 = ~x_215 &  n_652;
assign n_664 =  n_512 & ~n_663;
assign n_665 = ~n_662 & ~n_664;
assign n_666 = ~n_660 &  n_665;
assign n_667 = ~n_543 & ~n_519;
assign n_668 =  n_667 &  n_621;
assign n_669 = ~n_516 & ~n_668;
assign n_670 = ~n_666 &  n_669;
assign n_671 = ~n_656 & ~n_670;
assign n_672 =  n_633 & ~n_661;
assign n_673 = ~n_527 & ~n_672;
assign n_674 = ~n_671 &  n_673;
assign n_675 = ~n_654 & ~n_674;
assign n_676 = ~n_667 &  n_542;
assign n_677 = ~x_225 & ~n_676;
assign n_678 = ~n_675 &  n_677;
assign n_679 = ~n_651 & ~n_678;
assign n_680 =  x_331 & ~n_679;
assign n_681 = ~x_331 &  n_679;
assign n_682 = ~n_680 & ~n_681;
assign n_683 = ~i_25 &  x_225;
assign n_684 = ~n_518 & ~n_506;
assign n_685 =  n_684 &  n_658;
assign n_686 = ~x_330 & ~n_658;
assign n_687 = ~n_512 & ~n_686;
assign n_688 = ~n_685 &  n_687;
assign n_689 =  x_215 & ~n_684;
assign n_690 = ~n_517 & ~n_689;
assign n_691 =  n_512 &  n_690;
assign n_692 = ~n_633 & ~n_691;
assign n_693 = ~n_688 &  n_692;
assign n_694 =  n_684 &  n_633;
assign n_695 = ~n_527 & ~n_694;
assign n_696 = ~n_693 &  n_695;
assign n_697 =  n_690 &  n_527;
assign n_698 = ~x_225 & ~n_697;
assign n_699 = ~n_696 &  n_698;
assign n_700 = ~n_683 & ~n_699;
assign n_701 =  x_330 &  n_700;
assign n_702 = ~x_330 & ~n_700;
assign n_703 = ~n_701 & ~n_702;
assign n_704 =  i_26 &  x_225;
assign n_705 =  x_215 &  n_492;
assign n_706 = ~x_329 & ~n_705;
assign n_707 =  x_329 &  n_705;
assign n_708 = ~x_225 & ~n_707;
assign n_709 = ~n_706 &  n_708;
assign n_710 = ~n_704 & ~n_709;
assign n_711 =  x_329 & ~n_710;
assign n_712 = ~x_329 &  n_710;
assign n_713 = ~n_711 & ~n_712;
assign n_714 =  x_328 &  n_492;
assign n_715 = ~x_328 & ~n_492;
assign n_716 = ~n_714 & ~n_715;
assign n_717 = ~x_227 & ~n_1;
assign n_718 =  x_327 &  n_717;
assign n_719 = ~x_327 & ~n_717;
assign n_720 = ~n_718 & ~n_719;
assign n_721 = ~x_228 &  x_341;
assign n_722 =  x_326 &  n_721;
assign n_723 = ~x_326 & ~n_721;
assign n_724 = ~n_722 & ~n_723;
assign n_725 = ~x_228 & ~n_3;
assign n_726 =  x_272 &  n_1;
assign n_727 =  n_725 &  n_726;
assign n_728 =  x_325 & ~n_727;
assign n_729 = ~x_232 & ~n_728;
assign n_730 =  x_325 & ~n_729;
assign n_731 = ~x_325 &  n_729;
assign n_732 = ~n_730 & ~n_731;
assign n_733 = ~n_389 & ~n_93;
assign n_734 = ~n_5 &  n_733;
assign n_735 =  x_324 &  n_5;
assign n_736 = ~n_734 & ~n_735;
assign n_737 =  x_324 & ~n_736;
assign n_738 = ~x_324 &  n_736;
assign n_739 = ~n_737 & ~n_738;
assign n_740 =  i_148 &  x_308;
assign n_741 = ~x_308 &  x_323;
assign n_742 = ~n_740 & ~n_741;
assign n_743 =  x_323 & ~n_742;
assign n_744 = ~x_323 &  n_742;
assign n_745 = ~n_743 & ~n_744;
assign n_746 =  x_322 &  n_8;
assign n_747 =  x_312 & ~n_8;
assign n_748 =  i_138 &  n_747;
assign n_749 = ~n_746 & ~n_748;
assign n_750 =  x_322 & ~n_749;
assign n_751 = ~x_322 &  n_749;
assign n_752 = ~n_750 & ~n_751;
assign n_753 = ~x_315 & ~x_322;
assign n_754 = ~n_8 & ~n_753;
assign n_755 =  x_246 & ~n_223;
assign n_756 = ~n_754 & ~n_755;
assign n_757 =  x_321 & ~n_756;
assign n_758 = ~x_321 &  n_756;
assign n_759 = ~n_757 & ~n_758;
assign n_760 =  x_320 &  n_441;
assign n_761 = ~x_320 & ~n_441;
assign n_762 = ~n_760 & ~n_761;
assign n_763 = ~x_228 & ~x_244;
assign n_764 =  x_319 & ~n_763;
assign n_765 = ~x_319 &  n_763;
assign n_766 = ~n_764 & ~n_765;
assign n_767 = ~x_228 & ~x_319;
assign n_768 =  x_318 & ~n_767;
assign n_769 = ~x_318 &  n_767;
assign n_770 = ~n_768 & ~n_769;
assign n_771 = ~x_228 & ~x_318;
assign n_772 =  x_317 & ~n_771;
assign n_773 = ~x_317 &  n_771;
assign n_774 = ~n_772 & ~n_773;
assign n_775 = ~x_228 & ~x_317;
assign n_776 =  x_316 &  n_775;
assign n_777 = ~x_316 & ~n_775;
assign n_778 = ~n_776 & ~n_777;
assign n_779 =  x_315 &  n_8;
assign n_780 =  i_137 &  n_747;
assign n_781 = ~n_779 & ~n_780;
assign n_782 =  x_315 & ~n_781;
assign n_783 = ~x_315 &  n_781;
assign n_784 = ~n_782 & ~n_783;
assign n_785 =  i_20 &  x_300;
assign n_786 = ~x_300 &  x_314;
assign n_787 = ~n_785 & ~n_786;
assign n_788 =  x_314 & ~n_787;
assign n_789 = ~x_314 &  n_787;
assign n_790 = ~n_788 & ~n_789;
assign n_791 =  i_27 &  x_300;
assign n_792 = ~x_300 &  x_313;
assign n_793 = ~n_791 & ~n_792;
assign n_794 =  x_313 & ~n_793;
assign n_795 = ~x_313 &  n_793;
assign n_796 = ~n_794 & ~n_795;
assign n_797 =  x_312 & ~n_9;
assign n_798 = ~x_283 & ~n_223;
assign n_799 = ~n_797 &  n_798;
assign n_800 =  n_119 & ~n_799;
assign n_801 =  x_312 &  n_800;
assign n_802 = ~x_312 & ~n_800;
assign n_803 = ~n_801 & ~n_802;
assign n_804 =  x_311 &  n_8;
assign n_805 = ~n_213 &  n_221;
assign n_806 = ~n_804 & ~n_805;
assign n_807 =  x_311 & ~n_806;
assign n_808 = ~x_311 &  n_806;
assign n_809 = ~n_807 & ~n_808;
assign n_810 =  x_310 & ~n_3;
assign n_811 =  n_717 &  n_810;
assign n_812 =  n_98 & ~n_106;
assign n_813 = ~n_5 & ~n_812;
assign n_814 = ~n_389 &  n_813;
assign n_815 = ~n_811 & ~n_814;
assign n_816 = ~x_228 & ~n_815;
assign n_817 =  x_310 &  n_816;
assign n_818 = ~x_310 & ~n_816;
assign n_819 = ~n_817 & ~n_818;
assign n_820 =  x_221 &  x_300;
assign n_821 = ~x_309 & ~n_820;
assign n_822 = ~x_307 & ~n_821;
assign n_823 =  x_309 &  n_822;
assign n_824 = ~x_309 & ~n_822;
assign n_825 = ~n_823 & ~n_824;
assign n_826 =  x_308 &  n_820;
assign n_827 = ~x_308 & ~n_820;
assign n_828 = ~n_826 & ~n_827;
assign n_829 = ~i_136 & ~x_309;
assign n_830 =  x_228 & ~n_829;
assign n_831 = ~x_307 & ~n_830;
assign n_832 =  x_307 &  n_830;
assign n_833 = ~n_831 & ~n_832;
assign n_834 = ~x_306 & ~n_223;
assign n_835 =  x_306 &  n_223;
assign n_836 = ~n_834 & ~n_835;
assign n_837 =  x_304 &  n_8;
assign n_838 = ~x_283 & ~x_305;
assign n_839 = ~n_8 &  n_838;
assign n_840 = ~i_1 &  x_309;
assign n_841 = ~x_307 &  n_92;
assign n_842 = ~n_840 &  n_841;
assign n_843 =  n_839 &  n_842;
assign n_844 =  n_725 &  n_843;
assign n_845 = ~n_837 & ~n_844;
assign n_846 =  n_119 & ~n_845;
assign n_847 = ~n_8 &  n_846;
assign n_848 =  x_305 & ~n_9;
assign n_849 = ~x_283 & ~n_848;
assign n_850 = ~n_847 &  n_849;
assign n_851 =  n_119 & ~n_850;
assign n_852 =  x_305 &  n_851;
assign n_853 = ~x_305 & ~n_851;
assign n_854 = ~n_852 & ~n_853;
assign n_855 =  x_304 &  n_846;
assign n_856 = ~x_304 & ~n_846;
assign n_857 = ~n_855 & ~n_856;
assign n_858 =  x_303 &  n_8;
assign n_859 = ~x_283 & ~n_858;
assign n_860 =  x_303 & ~n_859;
assign n_861 = ~x_303 &  n_859;
assign n_862 = ~n_860 & ~n_861;
assign n_863 = ~x_381 &  x_382;
assign n_864 =  x_380 &  n_863;
assign n_865 =  x_384 &  n_864;
assign n_866 =  x_381 &  x_382;
assign n_867 = ~x_380 &  n_866;
assign n_868 =  x_390 &  n_867;
assign n_869 = ~n_865 & ~n_868;
assign n_870 =  x_381 & ~x_382;
assign n_871 =  x_380 &  n_870;
assign n_872 =  x_385 &  n_871;
assign n_873 =  x_380 &  n_866;
assign n_874 =  x_383 &  n_873;
assign n_875 = ~n_872 & ~n_874;
assign n_876 =  n_869 &  n_875;
assign n_877 = ~x_380 &  n_870;
assign n_878 =  x_389 &  n_877;
assign n_879 = ~x_381 & ~x_382;
assign n_880 =  x_380 &  n_879;
assign n_881 =  x_387 &  n_880;
assign n_882 = ~n_878 & ~n_881;
assign n_883 = ~x_380 &  n_879;
assign n_884 =  x_386 &  n_883;
assign n_885 = ~x_380 &  n_863;
assign n_886 =  x_388 &  n_885;
assign n_887 = ~n_884 & ~n_886;
assign n_888 =  n_882 &  n_887;
assign n_889 =  n_876 &  n_888;
assign n_890 =  i_187 &  n_880;
assign n_891 =  i_191 &  n_877;
assign n_892 = ~n_890 & ~n_891;
assign n_893 =  i_188 &  n_883;
assign n_894 =  i_190 &  n_885;
assign n_895 = ~n_893 & ~n_894;
assign n_896 =  n_892 &  n_895;
assign n_897 =  i_186 &  n_867;
assign n_898 =  i_185 &  n_864;
assign n_899 = ~n_897 & ~n_898;
assign n_900 =  i_189 &  n_871;
assign n_901 =  i_184 &  n_873;
assign n_902 = ~n_900 & ~n_901;
assign n_903 =  n_899 &  n_902;
assign n_904 =  n_896 &  n_903;
assign n_905 =  n_889 &  n_904;
assign n_906 =  x_352 &  n_864;
assign n_907 =  x_358 &  n_867;
assign n_908 = ~n_906 & ~n_907;
assign n_909 =  x_353 &  n_871;
assign n_910 =  x_351 &  n_873;
assign n_911 = ~n_909 & ~n_910;
assign n_912 =  n_908 &  n_911;
assign n_913 =  x_357 &  n_877;
assign n_914 =  x_355 &  n_880;
assign n_915 = ~n_913 & ~n_914;
assign n_916 =  x_354 &  n_883;
assign n_917 =  x_356 &  n_885;
assign n_918 = ~n_916 & ~n_917;
assign n_919 =  n_915 &  n_918;
assign n_920 =  n_912 &  n_919;
assign n_921 =  n_4 &  n_92;
assign n_922 = ~x_228 &  n_921;
assign n_923 = ~n_920 &  n_922;
assign n_924 = ~n_905 &  n_923;
assign n_925 =  x_302 &  n_924;
assign n_926 = ~x_302 & ~n_924;
assign n_927 = ~n_925 & ~n_926;
assign n_928 = ~i_42 & ~i_64;
assign n_929 =  i_42 &  i_64;
assign n_930 = ~n_928 & ~n_929;
assign n_931 = ~i_40 & ~i_63;
assign n_932 =  i_40 &  i_63;
assign n_933 = ~n_931 & ~n_932;
assign n_934 = ~i_43 & ~i_62;
assign n_935 =  i_43 &  i_62;
assign n_936 = ~n_934 & ~n_935;
assign n_937 = ~n_933 & ~n_936;
assign n_938 = ~n_930 &  n_937;
assign n_939 = ~i_39 &  i_61;
assign n_940 = ~i_41 &  i_65;
assign n_941 =  i_39 & ~i_61;
assign n_942 = ~n_940 & ~n_941;
assign n_943 = ~n_939 &  n_942;
assign n_944 = ~i_44 &  i_66;
assign n_945 = ~i_45 & ~i_67;
assign n_946 = ~n_944 & ~n_945;
assign n_947 =  i_45 &  i_67;
assign n_948 =  i_41 & ~i_65;
assign n_949 = ~n_947 & ~n_948;
assign n_950 =  n_946 &  n_949;
assign n_951 =  x_225 & ~x_249;
assign n_952 =  x_272 &  n_951;
assign n_953 =  i_44 & ~i_66;
assign n_954 =  n_119 & ~n_953;
assign n_955 =  n_952 &  n_954;
assign n_956 =  n_950 &  n_955;
assign n_957 =  n_943 &  n_956;
assign n_958 =  n_938 &  n_957;
assign n_959 = ~x_228 &  x_326;
assign n_960 = ~x_232 & ~n_959;
assign n_961 = ~n_3 &  n_960;
assign n_962 = ~n_958 &  n_961;
assign n_963 =  x_301 & ~n_962;
assign n_964 = ~x_301 &  n_962;
assign n_965 = ~n_963 & ~n_964;
assign n_966 = ~x_284 & ~x_300;
assign n_967 = ~x_232 & ~n_966;
assign n_968 =  x_218 &  x_316;
assign n_969 =  n_119 &  n_968;
assign n_970 = ~n_967 &  n_969;
assign n_971 =  x_300 &  n_970;
assign n_972 = ~x_300 & ~n_970;
assign n_973 = ~n_971 & ~n_972;
assign n_974 =  x_302 &  n_119;
assign n_975 =  x_350 &  n_873;
assign n_976 =  x_413 &  n_883;
assign n_977 = ~n_975 & ~n_976;
assign n_978 =  x_412 &  n_871;
assign n_979 =  x_409 &  n_885;
assign n_980 = ~n_978 & ~n_979;
assign n_981 =  n_977 &  n_980;
assign n_982 =  x_408 &  n_880;
assign n_983 =  x_410 &  n_877;
assign n_984 = ~n_982 & ~n_983;
assign n_985 =  x_414 &  n_864;
assign n_986 =  x_411 &  n_867;
assign n_987 = ~n_985 & ~n_986;
assign n_988 =  n_984 &  n_987;
assign n_989 =  n_981 &  n_988;
assign n_990 = ~n_905 & ~n_989;
assign n_991 =  n_920 & ~n_990;
assign n_992 = ~n_991 &  n_922;
assign n_993 = ~n_974 & ~n_992;
assign n_994 =  x_299 & ~n_993;
assign n_995 = ~x_299 &  n_993;
assign n_996 = ~n_994 & ~n_995;
assign n_997 =  x_349 &  n_920;
assign n_998 = ~x_400 & ~n_3;
assign n_999 = ~x_349 & ~x_351;
assign n_1000 =  n_998 & ~n_999;
assign n_1001 = ~n_997 &  n_1000;
assign n_1002 =  x_298 &  n_1001;
assign n_1003 = ~x_298 & ~n_1001;
assign n_1004 = ~n_1002 & ~n_1003;
assign n_1005 = ~x_232 & ~x_284;
assign n_1006 =  x_297 &  n_1005;
assign n_1007 = ~x_297 & ~n_1005;
assign n_1008 = ~n_1006 & ~n_1007;
assign n_1009 = ~x_226 & ~x_235;
assign n_1010 =  x_250 &  n_1009;
assign n_1011 = ~x_225 &  n_1010;
assign n_1012 = ~x_274 & ~x_293;
assign n_1013 =  x_274 &  x_293;
assign n_1014 = ~n_1012 & ~n_1013;
assign n_1015 = ~x_273 & ~x_285;
assign n_1016 =  x_273 &  x_285;
assign n_1017 = ~n_1015 & ~n_1016;
assign n_1018 =  i_59 & ~x_292;
assign n_1019 = ~i_59 &  x_292;
assign n_1020 = ~n_1018 & ~n_1019;
assign n_1021 = ~n_1017 &  n_1020;
assign n_1022 = ~n_1014 &  n_1021;
assign n_1023 = ~x_282 &  x_295;
assign n_1024 = ~i_60 &  x_294;
assign n_1025 = ~n_1023 & ~n_1024;
assign n_1026 =  x_275 & ~x_291;
assign n_1027 = ~x_275 &  x_291;
assign n_1028 = ~n_1026 & ~n_1027;
assign n_1029 =  n_1025 &  n_1028;
assign n_1030 =  i_128 & ~x_276;
assign n_1031 = ~i_128 &  x_276;
assign n_1032 = ~n_1030 & ~n_1031;
assign n_1033 =  x_282 & ~x_295;
assign n_1034 =  i_60 & ~x_294;
assign n_1035 = ~n_1033 & ~n_1034;
assign n_1036 =  n_1032 &  n_1035;
assign n_1037 =  n_1029 &  n_1036;
assign n_1038 =  n_1022 &  n_1037;
assign n_1039 = ~n_1011 &  n_1038;
assign n_1040 = ~x_296 &  x_297;
assign n_1041 = ~n_2 &  n_1040;
assign n_1042 =  n_1011 &  n_1041;
assign n_1043 =  i_18 &  i_19;
assign n_1044 =  x_217 &  n_1043;
assign n_1045 =  n_1042 &  n_1044;
assign n_1046 = ~n_1039 & ~n_1045;
assign n_1047 =  x_296 &  n_1046;
assign n_1048 = ~x_296 & ~n_1046;
assign n_1049 = ~n_1047 & ~n_1048;
assign n_1050 = ~i_18 & ~x_217;
assign n_1051 = ~i_19 &  n_1050;
assign n_1052 =  x_294 &  n_1051;
assign n_1053 = ~x_294 & ~n_1051;
assign n_1054 =  i_19 &  n_1050;
assign n_1055 = ~i_19 & ~n_1050;
assign n_1056 = ~n_1054 & ~n_1055;
assign n_1057 =  x_293 & ~n_1056;
assign n_1058 = ~x_293 &  n_1056;
assign n_1059 = ~n_1057 & ~n_1058;
assign n_1060 =  x_217 &  x_291;
assign n_1061 = ~i_18 &  n_1060;
assign n_1062 =  i_18 &  x_217;
assign n_1063 = ~x_291 &  n_1062;
assign n_1064 =  i_128 & ~n_1050;
assign n_1065 = ~n_1063 &  n_1064;
assign n_1066 = ~n_1061 & ~n_1065;
assign n_1067 =  n_1059 & ~n_1066;
assign n_1068 = ~n_1057 & ~n_1067;
assign n_1069 = ~n_1053 & ~n_1068;
assign n_1070 = ~n_1052 & ~n_1069;
assign n_1071 = ~x_295 &  n_1070;
assign n_1072 =  x_295 & ~n_1070;
assign n_1073 =  n_1010 &  n_494;
assign n_1074 = ~n_1072 &  n_1073;
assign n_1075 = ~n_1071 &  n_1074;
assign n_1076 =  i_130 &  x_242;
assign n_1077 = ~x_242 & ~n_1011;
assign n_1078 =  x_295 &  n_1077;
assign n_1079 = ~n_1076 & ~n_1078;
assign n_1080 = ~n_1075 &  n_1079;
assign n_1081 =  x_295 & ~n_1080;
assign n_1082 = ~x_295 &  n_1080;
assign n_1083 = ~n_1081 & ~n_1082;
assign n_1084 =  n_1053 &  n_1068;
assign n_1085 =  n_1073 & ~n_1084;
assign n_1086 =  n_1070 &  n_1085;
assign n_1087 = ~i_135 &  x_242;
assign n_1088 =  x_294 &  n_1077;
assign n_1089 = ~n_1087 & ~n_1088;
assign n_1090 = ~n_1086 &  n_1089;
assign n_1091 =  x_294 & ~n_1090;
assign n_1092 = ~x_294 &  n_1090;
assign n_1093 = ~n_1091 & ~n_1092;
assign n_1094 = ~n_1059 &  n_1066;
assign n_1095 = ~n_1067 &  n_1073;
assign n_1096 = ~n_1094 &  n_1095;
assign n_1097 =  i_134 &  x_242;
assign n_1098 =  x_293 &  n_1077;
assign n_1099 = ~n_1097 & ~n_1098;
assign n_1100 = ~n_1096 &  n_1099;
assign n_1101 =  x_293 & ~n_1100;
assign n_1102 = ~x_293 &  n_1100;
assign n_1103 = ~n_1101 & ~n_1102;
assign n_1104 = ~x_292 & ~n_1072;
assign n_1105 =  x_292 &  n_1072;
assign n_1106 = ~n_1105 &  n_1073;
assign n_1107 = ~n_1104 &  n_1106;
assign n_1108 =  i_132 &  x_242;
assign n_1109 =  x_292 &  n_1077;
assign n_1110 = ~n_1108 & ~n_1109;
assign n_1111 = ~n_1107 &  n_1110;
assign n_1112 =  x_292 & ~n_1111;
assign n_1113 = ~x_292 &  n_1111;
assign n_1114 = ~n_1112 & ~n_1113;
assign n_1115 =  x_291 &  n_1077;
assign n_1116 =  i_133 &  x_242;
assign n_1117 = ~x_217 & ~x_291;
assign n_1118 = ~n_1060 & ~n_1117;
assign n_1119 =  n_1118 &  n_1073;
assign n_1120 = ~n_1116 & ~n_1119;
assign n_1121 = ~n_1115 &  n_1120;
assign n_1122 =  x_291 & ~n_1121;
assign n_1123 = ~x_291 &  n_1121;
assign n_1124 = ~n_1122 & ~n_1123;
assign n_1125 = ~i_83 &  x_286;
assign n_1126 = ~x_289 &  n_1125;
assign n_1127 = ~x_292 &  n_1126;
assign n_1128 = ~i_74 & ~i_123;
assign n_1129 = ~i_107 &  n_1128;
assign n_1130 = ~i_128 & ~x_293;
assign n_1131 = ~i_74 & ~i_115;
assign n_1132 =  x_291 & ~x_295;
assign n_1133 =  n_1131 &  n_1132;
assign n_1134 =  n_1130 &  n_1133;
assign n_1135 =  n_1129 &  n_1134;
assign n_1136 =  n_1052 &  n_1135;
assign n_1137 = ~x_291 &  n_1130;
assign n_1138 =  n_1044 &  n_1137;
assign n_1139 =  x_295 &  n_1138;
assign n_1140 =  n_1084 &  n_1139;
assign n_1141 = ~n_1136 & ~n_1140;
assign n_1142 =  n_1127 & ~n_1141;
assign n_1143 =  x_294 & ~n_1051;
assign n_1144 = ~i_86 & ~i_94;
assign n_1145 = ~i_102 &  n_1144;
assign n_1146 = ~i_78 & ~i_115;
assign n_1147 =  n_1128 &  n_1146;
assign n_1148 =  n_1145 &  n_1147;
assign n_1149 = ~i_107 &  n_1148;
assign n_1150 = ~i_128 &  x_293;
assign n_1151 =  x_291 &  n_1150;
assign n_1152 =  n_1054 &  n_1151;
assign n_1153 =  n_1149 &  n_1152;
assign n_1154 =  i_128 & ~x_293;
assign n_1155 = ~i_19 &  n_1154;
assign n_1156 =  i_18 & ~x_217;
assign n_1157 =  x_291 &  n_1156;
assign n_1158 =  n_1155 &  n_1157;
assign n_1159 = ~i_19 &  n_1150;
assign n_1160 =  n_1063 &  n_1159;
assign n_1161 = ~i_94 &  n_1160;
assign n_1162 = ~n_1158 & ~n_1161;
assign n_1163 = ~i_91 & ~i_99;
assign n_1164 = ~i_86 &  n_1163;
assign n_1165 =  n_1126 &  n_1164;
assign n_1166 = ~n_1162 &  n_1165;
assign n_1167 = ~n_1153 & ~n_1166;
assign n_1168 = ~x_292 & ~x_295;
assign n_1169 = ~i_74 & ~i_78;
assign n_1170 =  n_1168 &  n_1169;
assign n_1171 = ~n_1167 &  n_1170;
assign n_1172 =  i_19 &  n_1156;
assign n_1173 =  i_128 &  x_293;
assign n_1174 =  x_291 &  n_1173;
assign n_1175 =  n_1172 &  n_1174;
assign n_1176 = ~i_110 & ~i_118;
assign n_1177 = ~x_295 &  n_1176;
assign n_1178 =  n_1175 &  n_1177;
assign n_1179 =  n_1127 &  n_1178;
assign n_1180 =  n_1149 &  n_1179;
assign n_1181 = ~n_1171 & ~n_1180;
assign n_1182 =  n_1143 & ~n_1181;
assign n_1183 =  n_1163 &  n_1146;
assign n_1184 =  n_1129 &  n_1183;
assign n_1185 = ~i_83 & ~x_291;
assign n_1186 =  n_1184 &  n_1185;
assign n_1187 = ~i_18 &  i_19;
assign n_1188 =  x_217 &  n_1187;
assign n_1189 =  x_286 &  n_1188;
assign n_1190 = ~i_118 & ~i_126;
assign n_1191 =  n_1189 & ~n_1190;
assign n_1192 = ~i_18 & ~i_19;
assign n_1193 =  x_217 &  n_1192;
assign n_1194 =  x_294 &  n_1154;
assign n_1195 =  n_1125 &  n_1168;
assign n_1196 =  n_1194 &  n_1195;
assign n_1197 =  n_1193 &  n_1196;
assign n_1198 = ~n_1191 & ~n_1197;
assign n_1199 =  n_1186 & ~n_1198;
assign n_1200 = ~n_1182 & ~n_1199;
assign n_1201 = ~n_1142 &  n_1200;
assign n_1202 =  n_1073 & ~n_1201;
assign n_1203 =  x_290 &  n_1077;
assign n_1204 = ~i_131 & ~i_132;
assign n_1205 =  n_1204 &  n_1116;
assign n_1206 = ~i_134 &  i_135;
assign n_1207 =  n_1206 &  n_1076;
assign n_1208 =  n_1205 &  n_1207;
assign n_1209 = ~n_1203 & ~n_1208;
assign n_1210 = ~n_1202 &  n_1209;
assign n_1211 =  x_290 & ~n_1210;
assign n_1212 = ~x_290 &  n_1210;
assign n_1213 = ~n_1211 & ~n_1212;
assign n_1214 = ~i_73 & ~i_85;
assign n_1215 = ~i_93 & ~i_101;
assign n_1216 = ~x_290 &  n_1215;
assign n_1217 =  n_1214 &  n_1216;
assign n_1218 = ~i_110 &  n_1217;
assign n_1219 = ~i_118 &  n_1218;
assign n_1220 =  n_1145 &  n_1219;
assign n_1221 = ~i_70 & ~i_106;
assign n_1222 = ~i_114 &  n_1221;
assign n_1223 = ~i_90 & ~i_98;
assign n_1224 = ~i_122 &  n_1223;
assign n_1225 =  n_1222 &  n_1224;
assign n_1226 = ~i_76 & ~i_126;
assign n_1227 =  x_286 &  n_1226;
assign n_1228 =  n_1184 &  n_1227;
assign n_1229 =  n_1225 &  n_1228;
assign n_1230 =  n_1220 &  n_1229;
assign n_1231 = ~i_109 & ~i_117;
assign n_1232 = ~i_125 &  n_1231;
assign n_1233 = ~i_75 & ~i_79;
assign n_1234 = ~i_87 & ~i_95;
assign n_1235 =  n_1233 &  n_1234;
assign n_1236 =  n_1232 &  n_1235;
assign n_1237 = ~i_113 & ~i_119;
assign n_1238 = ~i_127 & ~x_287;
assign n_1239 =  n_1237 &  n_1238;
assign n_1240 = ~i_69 & ~i_103;
assign n_1241 = ~i_105 & ~i_111;
assign n_1242 =  n_1240 &  n_1241;
assign n_1243 = ~i_72 & ~i_77;
assign n_1244 = ~i_89 & ~i_97;
assign n_1245 =  n_1243 &  n_1244;
assign n_1246 =  n_1242 &  n_1245;
assign n_1247 =  n_1239 &  n_1246;
assign n_1248 =  n_1236 &  n_1247;
assign n_1249 =  x_292 &  x_295;
assign n_1250 =  x_294 &  n_1249;
assign n_1251 = ~n_1130 &  n_1250;
assign n_1252 =  n_1251 & ~n_1173;
assign n_1253 = ~i_71 & ~i_116;
assign n_1254 = ~i_124 &  n_1253;
assign n_1255 = ~i_82 & ~i_108;
assign n_1256 = ~x_288 &  n_1255;
assign n_1257 =  n_1254 &  n_1256;
assign n_1258 = ~i_100 &  n_1257;
assign n_1259 = ~i_84 & ~i_92;
assign n_1260 = ~i_81 & ~i_121;
assign n_1261 =  n_1259 &  n_1260;
assign n_1262 = ~n_1051 &  n_1261;
assign n_1263 =  n_1258 &  n_1262;
assign n_1264 = ~n_1252 &  n_1263;
assign n_1265 =  n_1248 &  n_1264;
assign n_1266 =  n_1230 &  n_1265;
assign n_1267 =  i_112 &  n_1266;
assign n_1268 =  n_1267 &  n_1188;
assign n_1269 = ~i_83 & ~i_112;
assign n_1270 = ~x_289 &  n_1269;
assign n_1271 =  n_1266 &  n_1270;
assign n_1272 =  n_1172 &  n_1271;
assign n_1273 =  x_292 &  n_1243;
assign n_1274 = ~i_100 &  n_1259;
assign n_1275 =  n_1273 &  n_1274;
assign n_1276 =  n_1225 &  n_1257;
assign n_1277 =  n_1275 &  n_1276;
assign n_1278 =  n_1154 &  n_1190;
assign n_1279 =  n_1145 &  n_1274;
assign n_1280 =  n_1278 &  n_1279;
assign n_1281 = ~i_103 &  x_295;
assign n_1282 = ~i_108 & ~i_111;
assign n_1283 =  n_1281 &  n_1282;
assign n_1284 =  n_1254 &  n_1283;
assign n_1285 =  n_1236 &  n_1284;
assign n_1286 =  n_1280 &  n_1285;
assign n_1287 =  n_1218 &  n_1186;
assign n_1288 =  n_1286 &  n_1287;
assign n_1289 =  n_1277 &  n_1288;
assign n_1290 =  n_1230 &  n_1289;
assign n_1291 = ~i_121 &  n_1143;
assign n_1292 = ~i_76 & ~i_81;
assign n_1293 =  n_1244 &  n_1292;
assign n_1294 = ~i_105 &  n_1193;
assign n_1295 =  n_1293 &  n_1294;
assign n_1296 =  n_1291 &  n_1295;
assign n_1297 =  n_1248 &  n_1296;
assign n_1298 =  n_1290 &  n_1297;
assign n_1299 =  i_104 &  n_1054;
assign n_1300 = ~x_291 &  n_1154;
assign n_1301 = ~i_88 & ~n_1300;
assign n_1302 =  n_1251 &  n_1301;
assign n_1303 =  n_1302 &  n_1160;
assign n_1304 = ~n_1299 & ~n_1303;
assign n_1305 =  n_1143 & ~n_1304;
assign n_1306 =  n_1053 &  n_1168;
assign n_1307 =  n_1138 &  n_1306;
assign n_1308 =  x_287 &  n_1050;
assign n_1309 =  i_88 &  n_1156;
assign n_1310 = ~n_1308 & ~n_1309;
assign n_1311 = ~i_19 &  x_294;
assign n_1312 = ~n_1310 &  n_1311;
assign n_1313 = ~n_1307 & ~n_1312;
assign n_1314 = ~n_1305 &  n_1313;
assign n_1315 = ~n_1298 &  n_1314;
assign n_1316 = ~n_1272 &  n_1315;
assign n_1317 = ~n_1268 &  n_1316;
assign n_1318 =  n_1073 & ~n_1317;
assign n_1319 = ~i_130 &  n_1206;
assign n_1320 =  n_1319 &  n_1205;
assign n_1321 =  x_289 &  n_1077;
assign n_1322 = ~n_1320 & ~n_1321;
assign n_1323 = ~n_1318 &  n_1322;
assign n_1324 =  x_289 & ~n_1323;
assign n_1325 = ~x_289 &  n_1323;
assign n_1326 = ~n_1324 & ~n_1325;
assign n_1327 = ~i_126 &  n_1219;
assign n_1328 = ~x_294 & ~x_295;
assign n_1329 = ~n_1051 &  n_1328;
assign n_1330 =  n_1275 &  n_1329;
assign n_1331 =  n_1327 &  n_1330;
assign n_1332 = ~i_108 &  n_1173;
assign n_1333 =  n_1188 &  n_1332;
assign n_1334 =  n_1145 &  n_1333;
assign n_1335 =  n_1331 &  n_1334;
assign n_1336 =  n_1053 &  n_1220;
assign n_1337 = ~x_295 &  n_1273;
assign n_1338 =  n_1193 &  n_1278;
assign n_1339 =  n_1337 &  n_1338;
assign n_1340 =  n_1336 &  n_1339;
assign n_1341 = ~n_1335 & ~n_1340;
assign n_1342 =  x_286 &  n_1186;
assign n_1343 = ~n_1341 &  n_1342;
assign n_1344 =  x_294 &  n_1138;
assign n_1345 =  x_292 &  n_1328;
assign n_1346 =  n_1175 &  n_1345;
assign n_1347 =  n_1053 &  n_1160;
assign n_1348 = ~n_1346 & ~n_1347;
assign n_1349 =  n_1259 & ~n_1348;
assign n_1350 = ~n_1344 & ~n_1349;
assign n_1351 =  n_1337 & ~n_1350;
assign n_1352 =  x_291 & ~x_294;
assign n_1353 =  n_1130 &  n_1352;
assign n_1354 =  n_1051 &  n_1353;
assign n_1355 = ~i_84 &  n_1243;
assign n_1356 =  n_1158 &  n_1355;
assign n_1357 = ~n_1354 & ~n_1356;
assign n_1358 =  n_1345 & ~n_1357;
assign n_1359 =  n_1153 &  n_1331;
assign n_1360 = ~n_1358 & ~n_1359;
assign n_1361 = ~n_1351 &  n_1360;
assign n_1362 = ~n_1343 &  n_1361;
assign n_1363 =  n_1073 & ~n_1362;
assign n_1364 =  x_288 &  n_1077;
assign n_1365 = ~i_131 &  i_133;
assign n_1366 =  n_1108 &  n_1365;
assign n_1367 = ~i_134 &  n_1087;
assign n_1368 = ~i_130 &  n_1367;
assign n_1369 =  n_1366 &  n_1368;
assign n_1370 = ~n_1364 & ~n_1369;
assign n_1371 = ~n_1363 &  n_1370;
assign n_1372 =  x_288 & ~n_1371;
assign n_1373 = ~x_288 &  n_1371;
assign n_1374 = ~n_1372 & ~n_1373;
assign n_1375 =  n_1217 &  n_1126;
assign n_1376 = ~n_1055 &  n_1281;
assign n_1377 =  n_1236 &  n_1376;
assign n_1378 =  n_1375 &  n_1377;
assign n_1379 =  n_1153 &  n_1378;
assign n_1380 =  n_1336 &  n_1379;
assign n_1381 = ~i_103 & ~x_291;
assign n_1382 =  n_1173 &  n_1381;
assign n_1383 =  n_1053 &  n_1382;
assign n_1384 =  n_1236 &  n_1189;
assign n_1385 =  n_1383 &  n_1384;
assign n_1386 =  n_1291 &  n_1138;
assign n_1387 =  n_1053 &  n_1175;
assign n_1388 = ~n_1386 & ~n_1387;
assign n_1389 = ~i_113 &  x_286;
assign n_1390 = ~x_289 &  n_1389;
assign n_1391 =  n_1043 &  n_1390;
assign n_1392 = ~n_1388 &  n_1391;
assign n_1393 = ~n_1385 & ~n_1392;
assign n_1394 = ~i_105 &  x_295;
assign n_1395 =  n_1148 &  n_1394;
assign n_1396 =  n_1218 &  n_1395;
assign n_1397 = ~n_1393 &  n_1396;
assign n_1398 = ~n_1380 & ~n_1397;
assign n_1399 =  n_1293 & ~n_1398;
assign n_1400 = ~n_1399 & ~n_1354;
assign n_1401 = ~n_1400 &  n_1277;
assign n_1402 =  n_1258 &  n_1160;
assign n_1403 = ~n_1328 &  n_1158;
assign n_1404 = ~n_1402 & ~n_1403;
assign n_1405 =  x_295 &  n_1292;
assign n_1406 =  n_1222 &  n_1405;
assign n_1407 =  n_1273 &  n_1406;
assign n_1408 =  n_1053 &  n_1148;
assign n_1409 =  n_1407 &  n_1408;
assign n_1410 =  n_1375 &  n_1409;
assign n_1411 = ~n_1404 &  n_1410;
assign n_1412 =  n_1327 &  n_1411;
assign n_1413 = ~i_76 & ~x_294;
assign n_1414 =  n_1243 &  n_1413;
assign n_1415 =  n_1193 &  n_1414;
assign n_1416 =  n_1290 &  n_1415;
assign n_1417 = ~n_1412 & ~n_1416;
assign n_1418 = ~n_1401 &  n_1417;
assign n_1419 =  n_1073 & ~n_1418;
assign n_1420 =  x_287 &  n_1077;
assign n_1421 =  i_130 &  n_1367;
assign n_1422 =  n_1366 &  n_1421;
assign n_1423 = ~n_1420 & ~n_1422;
assign n_1424 = ~n_1419 &  n_1423;
assign n_1425 =  x_287 & ~n_1424;
assign n_1426 = ~x_287 &  n_1424;
assign n_1427 = ~n_1425 & ~n_1426;
assign n_1428 =  n_1172 &  n_1267;
assign n_1429 =  n_1044 &  n_1271;
assign n_1430 =  i_18 &  n_1249;
assign n_1431 = ~n_1118 &  n_1430;
assign n_1432 =  n_1155 &  n_1431;
assign n_1433 =  x_287 &  n_1193;
assign n_1434 =  i_96 &  n_1054;
assign n_1435 =  i_69 &  n_1051;
assign n_1436 = ~n_1434 & ~n_1435;
assign n_1437 = ~n_1433 &  n_1436;
assign n_1438 = ~n_1432 &  n_1437;
assign n_1439 =  x_294 & ~n_1438;
assign n_1440 = ~i_96 &  n_1188;
assign n_1441 =  n_1151 &  n_1440;
assign n_1442 =  n_1302 &  n_1441;
assign n_1443 = ~n_1442 &  n_1073;
assign n_1444 = ~n_1439 &  n_1443;
assign n_1445 = ~n_1429 &  n_1444;
assign n_1446 = ~n_1428 &  n_1445;
assign n_1447 =  x_286 &  n_1077;
assign n_1448 = ~i_133 &  n_1204;
assign n_1449 =  n_1319 &  n_1448;
assign n_1450 =  x_242 & ~n_1449;
assign n_1451 = ~n_1447 & ~n_1450;
assign n_1452 = ~n_1446 &  n_1451;
assign n_1453 =  x_286 & ~n_1452;
assign n_1454 = ~x_286 &  n_1452;
assign n_1455 = ~n_1453 & ~n_1454;
assign n_1456 =  i_129 &  x_242;
assign n_1457 =  n_1011 &  n_1105;
assign n_1458 = ~x_285 & ~n_1457;
assign n_1459 =  x_285 &  n_1457;
assign n_1460 = ~x_242 & ~n_1459;
assign n_1461 = ~n_1458 &  n_1460;
assign n_1462 = ~n_1456 & ~n_1461;
assign n_1463 =  x_285 & ~n_1462;
assign n_1464 = ~x_285 &  n_1462;
assign n_1465 = ~n_1463 & ~n_1464;
assign n_1466 =  x_284 &  n_967;
assign n_1467 = ~x_284 & ~n_967;
assign n_1468 = ~n_1466 & ~n_1467;
assign n_1469 =  x_283 &  x_307;
assign n_1470 = ~x_283 & ~x_307;
assign n_1471 = ~n_1469 & ~n_1470;
assign n_1472 =  x_275 &  x_276;
assign n_1473 = ~x_274 &  n_1472;
assign n_1474 = ~x_275 & ~x_276;
assign n_1475 =  x_274 &  n_1474;
assign n_1476 =  i_99 & ~x_278;
assign n_1477 =  i_102 &  x_280;
assign n_1478 = ~n_1476 & ~n_1477;
assign n_1479 =  i_57 &  i_98;
assign n_1480 =  i_97 &  x_277;
assign n_1481 = ~n_1479 & ~n_1480;
assign n_1482 =  n_1478 &  n_1481;
assign n_1483 =  i_103 &  x_281;
assign n_1484 =  i_58 &  i_101;
assign n_1485 = ~n_1483 & ~n_1484;
assign n_1486 =  i_100 &  x_279;
assign n_1487 =  i_56 &  i_96;
assign n_1488 = ~n_1486 & ~n_1487;
assign n_1489 =  n_1485 &  n_1488;
assign n_1490 =  n_1482 &  n_1489;
assign n_1491 =  n_1475 & ~n_1490;
assign n_1492 =  x_275 & ~x_276;
assign n_1493 =  x_274 &  n_1492;
assign n_1494 =  i_119 &  x_281;
assign n_1495 =  i_56 &  i_112;
assign n_1496 = ~n_1494 & ~n_1495;
assign n_1497 =  i_58 &  i_117;
assign n_1498 =  i_113 &  x_277;
assign n_1499 = ~n_1497 & ~n_1498;
assign n_1500 =  n_1496 &  n_1499;
assign n_1501 = ~x_275 &  x_276;
assign n_1502 =  x_274 &  n_1501;
assign n_1503 =  i_115 & ~x_278;
assign n_1504 =  i_118 &  x_280;
assign n_1505 = ~n_1503 & ~n_1504;
assign n_1506 =  i_116 &  x_279;
assign n_1507 =  i_57 &  i_114;
assign n_1508 = ~n_1506 & ~n_1507;
assign n_1509 =  n_1505 &  n_1508;
assign n_1510 =  n_1502 &  n_1509;
assign n_1511 =  n_1500 &  n_1510;
assign n_1512 =  i_57 &  i_122;
assign n_1513 =  i_123 & ~x_278;
assign n_1514 = ~n_1512 & ~n_1513;
assign n_1515 =  i_124 &  x_279;
assign n_1516 =  i_58 &  i_125;
assign n_1517 = ~n_1515 & ~n_1516;
assign n_1518 =  n_1514 &  n_1517;
assign n_1519 =  i_126 &  x_280;
assign n_1520 =  i_56 &  i_120;
assign n_1521 = ~n_1519 & ~n_1520;
assign n_1522 =  i_127 &  x_281;
assign n_1523 =  i_121 &  x_277;
assign n_1524 = ~n_1522 & ~n_1523;
assign n_1525 =  n_1521 &  n_1524;
assign n_1526 = ~n_1502 &  n_1525;
assign n_1527 =  n_1518 &  n_1526;
assign n_1528 = ~n_1511 & ~n_1527;
assign n_1529 = ~n_1493 & ~n_1528;
assign n_1530 =  i_58 &  i_109;
assign n_1531 =  i_110 &  x_280;
assign n_1532 = ~n_1530 & ~n_1531;
assign n_1533 =  i_111 &  x_281;
assign n_1534 =  i_107 & ~x_278;
assign n_1535 = ~n_1533 & ~n_1534;
assign n_1536 =  n_1532 &  n_1535;
assign n_1537 =  i_57 &  i_106;
assign n_1538 =  i_105 &  x_277;
assign n_1539 = ~n_1537 & ~n_1538;
assign n_1540 =  i_56 &  i_104;
assign n_1541 =  i_108 &  x_279;
assign n_1542 = ~n_1540 & ~n_1541;
assign n_1543 =  n_1539 &  n_1542;
assign n_1544 =  n_1493 &  n_1543;
assign n_1545 =  n_1536 &  n_1544;
assign n_1546 = ~n_1475 & ~n_1545;
assign n_1547 = ~n_1529 &  n_1546;
assign n_1548 = ~n_1491 & ~n_1547;
assign n_1549 = ~n_1473 & ~n_1548;
assign n_1550 = ~x_274 &  n_1501;
assign n_1551 =  i_58 &  i_93;
assign n_1552 =  i_91 & ~x_278;
assign n_1553 = ~n_1551 & ~n_1552;
assign n_1554 =  i_94 &  x_280;
assign n_1555 =  i_95 &  x_281;
assign n_1556 = ~n_1554 & ~n_1555;
assign n_1557 =  n_1553 &  n_1556;
assign n_1558 =  i_89 &  x_277;
assign n_1559 =  i_57 &  i_90;
assign n_1560 = ~n_1558 & ~n_1559;
assign n_1561 =  i_56 &  i_88;
assign n_1562 =  i_92 &  x_279;
assign n_1563 = ~n_1561 & ~n_1562;
assign n_1564 =  n_1560 &  n_1563;
assign n_1565 =  n_1557 &  n_1564;
assign n_1566 =  n_1473 & ~n_1565;
assign n_1567 = ~n_1550 & ~n_1566;
assign n_1568 = ~n_1549 &  n_1567;
assign n_1569 = ~x_274 &  n_1492;
assign n_1570 =  i_84 &  x_279;
assign n_1571 =  i_87 &  x_281;
assign n_1572 = ~n_1570 & ~n_1571;
assign n_1573 =  i_57 &  i_82;
assign n_1574 =  i_86 &  x_280;
assign n_1575 = ~n_1573 & ~n_1574;
assign n_1576 =  n_1572 &  n_1575;
assign n_1577 =  i_81 &  x_277;
assign n_1578 =  i_58 &  i_85;
assign n_1579 = ~n_1577 & ~n_1578;
assign n_1580 =  i_83 & ~x_278;
assign n_1581 =  i_56 &  i_80;
assign n_1582 = ~n_1580 & ~n_1581;
assign n_1583 =  n_1579 &  n_1582;
assign n_1584 =  n_1550 &  n_1583;
assign n_1585 =  n_1576 &  n_1584;
assign n_1586 = ~n_1569 & ~n_1585;
assign n_1587 = ~n_1568 &  n_1586;
assign n_1588 = ~x_274 &  n_1474;
assign n_1589 =  i_58 &  x_290;
assign n_1590 = ~x_278 &  x_289;
assign n_1591 = ~n_1589 & ~n_1590;
assign n_1592 =  i_78 &  x_280;
assign n_1593 =  i_79 &  x_281;
assign n_1594 = ~n_1592 & ~n_1593;
assign n_1595 =  n_1591 &  n_1594;
assign n_1596 =  i_56 &  x_287;
assign n_1597 =  i_57 &  x_288;
assign n_1598 = ~n_1596 & ~n_1597;
assign n_1599 =  i_77 &  x_279;
assign n_1600 =  i_76 &  x_277;
assign n_1601 = ~n_1599 & ~n_1600;
assign n_1602 =  n_1598 &  n_1601;
assign n_1603 =  n_1595 &  n_1602;
assign n_1604 =  n_1569 & ~n_1603;
assign n_1605 = ~n_1588 & ~n_1604;
assign n_1606 = ~n_1587 &  n_1605;
assign n_1607 =  i_57 &  i_71;
assign n_1608 =  i_75 &  x_281;
assign n_1609 = ~n_1607 & ~n_1608;
assign n_1610 =  i_58 &  i_73;
assign n_1611 =  i_74 &  x_280;
assign n_1612 = ~n_1610 & ~n_1611;
assign n_1613 =  n_1609 &  n_1612;
assign n_1614 =  i_72 &  x_279;
assign n_1615 = ~x_278 & ~x_286;
assign n_1616 = ~n_1614 & ~n_1615;
assign n_1617 =  i_56 &  i_69;
assign n_1618 =  i_70 &  x_277;
assign n_1619 = ~n_1617 & ~n_1618;
assign n_1620 =  n_1616 &  n_1619;
assign n_1621 =  n_1588 &  n_1620;
assign n_1622 =  n_1613 &  n_1621;
assign n_1623 = ~n_1017 & ~n_1622;
assign n_1624 = ~n_1606 &  n_1623;
assign n_1625 = ~x_270 &  n_1;
assign n_1626 = ~x_262 & ~n_1625;
assign n_1627 = ~x_270 & ~x_341;
assign n_1628 = ~x_228 & ~n_1627;
assign n_1629 = ~x_232 & ~n_1628;
assign n_1630 =  n_1042 & ~n_1626;
assign n_1631 =  n_1629 & ~n_1630;
assign n_1632 = ~n_1626 &  n_1631;
assign n_1633 = ~n_1624 &  n_1632;
assign n_1634 =  x_274 &  n_1472;
assign n_1635 =  i_60 &  n_1634;
assign n_1636 =  x_282 &  n_1635;
assign n_1637 = ~x_282 & ~n_1635;
assign n_1638 = ~n_1636 & ~n_1637;
assign n_1639 =  n_1633 &  n_1638;
assign n_1640 = ~i_28 &  n_1628;
assign n_1641 = ~x_232 & ~n_1640;
assign n_1642 = ~i_208 & ~n_1641;
assign n_1643 =  i_35 &  i_36;
assign n_1644 = ~n_1010 &  n_1643;
assign n_1645 =  x_236 &  n_1010;
assign n_1646 =  x_237 &  n_1645;
assign n_1647 = ~n_1644 & ~n_1646;
assign n_1648 =  x_238 &  n_1010;
assign n_1649 =  i_34 & ~n_1010;
assign n_1650 = ~n_1648 & ~n_1649;
assign n_1651 = ~n_1647 & ~n_1650;
assign n_1652 =  x_239 &  n_1010;
assign n_1653 =  i_33 & ~n_1010;
assign n_1654 = ~n_1652 & ~n_1653;
assign n_1655 =  n_1651 & ~n_1654;
assign n_1656 =  i_32 & ~n_1010;
assign n_1657 =  x_240 &  n_1010;
assign n_1658 = ~n_1656 & ~n_1657;
assign n_1659 =  n_1655 & ~n_1658;
assign n_1660 = ~n_1655 &  n_1658;
assign n_1661 = ~n_1659 & ~n_1660;
assign n_1662 =  n_1630 & ~n_1661;
assign n_1663 = ~x_282 & ~n_1630;
assign n_1664 = ~n_1662 & ~n_1663;
assign n_1665 =  n_1629 & ~n_1664;
assign n_1666 = ~n_1642 & ~n_1665;
assign n_1667 = ~n_1633 &  n_1666;
assign n_1668 = ~n_1639 & ~n_1667;
assign n_1669 =  x_282 & ~n_1668;
assign n_1670 = ~x_282 &  n_1668;
assign n_1671 = ~n_1669 & ~n_1670;
assign n_1672 =  n_1629 &  n_1630;
assign n_1673 =  x_281 & ~n_1010;
assign n_1674 = ~x_241 &  n_1010;
assign n_1675 = ~n_1651 &  n_1654;
assign n_1676 = ~n_1655 & ~n_1675;
assign n_1677 =  n_1674 &  n_1676;
assign n_1678 = ~n_1658 &  n_1677;
assign n_1679 = ~n_1673 & ~n_1678;
assign n_1680 =  n_1672 & ~n_1679;
assign n_1681 =  x_281 &  n_1631;
assign n_1682 =  i_208 & ~i_209;
assign n_1683 =  i_211 &  n_1682;
assign n_1684 = ~i_29 & ~x_232;
assign n_1685 =  i_28 & ~i_30;
assign n_1686 =  n_1684 &  n_1685;
assign n_1687 = ~n_1683 & ~n_1686;
assign n_1688 = ~n_1629 & ~n_1687;
assign n_1689 = ~n_1681 & ~n_1688;
assign n_1690 = ~n_1680 &  n_1689;
assign n_1691 = ~n_1633 & ~n_1690;
assign n_1692 =  i_59 &  n_1636;
assign n_1693 = ~i_59 & ~n_1636;
assign n_1694 = ~n_1692 & ~n_1693;
assign n_1695 =  n_1633 & ~n_1694;
assign n_1696 = ~i_60 & ~n_1634;
assign n_1697 = ~n_1635 & ~n_1696;
assign n_1698 =  x_282 &  n_1697;
assign n_1699 =  n_1695 &  n_1698;
assign n_1700 = ~n_1691 & ~n_1699;
assign n_1701 =  x_281 & ~n_1700;
assign n_1702 = ~x_281 &  n_1700;
assign n_1703 = ~n_1701 & ~n_1702;
assign n_1704 =  x_280 & ~n_1010;
assign n_1705 = ~x_240 &  n_1677;
assign n_1706 = ~n_1704 & ~n_1705;
assign n_1707 =  n_1672 & ~n_1706;
assign n_1708 =  x_280 &  n_1631;
assign n_1709 =  i_211 &  i_212;
assign n_1710 =  i_209 &  n_1709;
assign n_1711 =  x_232 & ~n_1710;
assign n_1712 =  n_1709 &  n_1711;
assign n_1713 = ~i_28 &  i_30;
assign n_1714 = ~i_29 &  n_1713;
assign n_1715 = ~i_28 &  n_1684;
assign n_1716 = ~n_1714 &  n_1715;
assign n_1717 = ~n_1712 & ~n_1716;
assign n_1718 = ~n_1629 & ~n_1717;
assign n_1719 = ~n_1708 & ~n_1718;
assign n_1720 = ~n_1707 &  n_1719;
assign n_1721 = ~n_1633 & ~n_1720;
assign n_1722 =  n_1637 & ~n_1696;
assign n_1723 =  n_1695 &  n_1722;
assign n_1724 = ~n_1721 & ~n_1723;
assign n_1725 =  x_280 & ~n_1724;
assign n_1726 = ~x_280 &  n_1724;
assign n_1727 = ~n_1725 & ~n_1726;
assign n_1728 = ~x_278 & ~n_1630;
assign n_1729 = ~i_37 & ~n_1010;
assign n_1730 = ~n_1729 & ~n_1674;
assign n_1731 =  n_1730 &  n_1659;
assign n_1732 = ~n_1730 & ~n_1659;
assign n_1733 = ~n_1731 & ~n_1732;
assign n_1734 = ~n_1733 & ~n_1676;
assign n_1735 =  n_1662 &  n_1734;
assign n_1736 = ~n_1728 & ~n_1735;
assign n_1737 =  n_1629 & ~n_1736;
assign n_1738 = ~x_232 & ~n_1714;
assign n_1739 = ~n_1629 & ~n_1738;
assign n_1740 = ~n_1711 &  n_1739;
assign n_1741 = ~n_1737 & ~n_1740;
assign n_1742 = ~n_1633 & ~n_1741;
assign n_1743 = ~n_1638 & ~n_1697;
assign n_1744 =  n_1695 &  n_1743;
assign n_1745 = ~n_1742 & ~n_1744;
assign n_1746 =  x_278 &  n_1745;
assign n_1747 = ~x_278 & ~n_1745;
assign n_1748 = ~n_1746 & ~n_1747;
assign n_1749 =  x_277 & ~n_1010;
assign n_1750 =  n_1010 & ~n_1676;
assign n_1751 =  n_1733 &  n_1750;
assign n_1752 =  n_1661 &  n_1751;
assign n_1753 = ~n_1749 & ~n_1752;
assign n_1754 =  n_1672 & ~n_1753;
assign n_1755 =  x_277 &  n_1631;
assign n_1756 =  i_208 &  i_209;
assign n_1757 = ~i_211 &  n_1756;
assign n_1758 =  i_29 & ~x_232;
assign n_1759 =  i_28 &  i_30;
assign n_1760 =  n_1758 &  n_1759;
assign n_1761 = ~n_1757 & ~n_1760;
assign n_1762 = ~n_1629 & ~n_1761;
assign n_1763 = ~n_1755 & ~n_1762;
assign n_1764 = ~n_1754 &  n_1763;
assign n_1765 = ~n_1633 & ~n_1764;
assign n_1766 =  n_1694 & ~n_1697;
assign n_1767 =  n_1639 &  n_1766;
assign n_1768 = ~n_1765 & ~n_1767;
assign n_1769 =  x_277 & ~n_1768;
assign n_1770 = ~x_277 &  n_1768;
assign n_1771 = ~n_1769 & ~n_1770;
assign n_1772 = ~i_54 & ~n_1629;
assign n_1773 = ~x_236 & ~x_237;
assign n_1774 =  n_1630 & ~n_1773;
assign n_1775 =  n_1647 &  n_1774;
assign n_1776 =  x_276 & ~n_1630;
assign n_1777 =  n_1629 & ~n_1776;
assign n_1778 = ~n_1775 &  n_1777;
assign n_1779 = ~n_1772 & ~n_1778;
assign n_1780 = ~n_1633 & ~n_1779;
assign n_1781 = ~n_1492 & ~n_1501;
assign n_1782 =  n_1633 &  n_1781;
assign n_1783 = ~n_1780 & ~n_1782;
assign n_1784 =  x_276 &  n_1783;
assign n_1785 = ~x_276 & ~n_1783;
assign n_1786 = ~n_1784 & ~n_1785;
assign n_1787 = ~i_53 & ~n_1629;
assign n_1788 =  n_1630 & ~n_1645;
assign n_1789 =  x_275 & ~n_1630;
assign n_1790 =  n_1629 & ~n_1789;
assign n_1791 = ~n_1788 &  n_1790;
assign n_1792 = ~n_1787 & ~n_1791;
assign n_1793 = ~n_1633 &  n_1792;
assign n_1794 = ~x_275 &  n_1633;
assign n_1795 = ~n_1793 & ~n_1794;
assign n_1796 =  x_275 & ~n_1795;
assign n_1797 = ~x_275 &  n_1795;
assign n_1798 = ~n_1796 & ~n_1797;
assign n_1799 =  x_307 &  x_348;
assign n_1800 = ~x_425 & ~n_839;
assign n_1801 = ~n_223 &  n_1800;
assign n_1802 = ~i_155 &  x_214;
assign n_1803 =  n_839 & ~n_1802;
assign n_1804 =  x_424 &  n_223;
assign n_1805 = ~n_1803 & ~n_1804;
assign n_1806 = ~n_1801 &  n_1805;
assign n_1807 = ~x_307 & ~n_1806;
assign n_1808 = ~n_1799 & ~n_1807;
assign n_1809 =  x_425 &  n_1808;
assign n_1810 = ~x_425 & ~n_1808;
assign n_1811 = ~n_1809 & ~n_1810;
assign n_1812 = ~x_424 & ~n_839;
assign n_1813 = ~n_1803 & ~n_1812;
assign n_1814 = ~x_307 & ~n_1813;
assign n_1815 =  x_307 &  x_344;
assign n_1816 = ~n_1814 & ~n_1815;
assign n_1817 =  x_424 &  n_1816;
assign n_1818 = ~x_424 & ~n_1816;
assign n_1819 = ~n_1817 & ~n_1818;
assign n_1820 =  x_307 & ~x_345;
assign n_1821 = ~x_304 & ~n_8;
assign n_1822 =  n_20 &  n_1821;
assign n_1823 = ~x_423 &  n_1822;
assign n_1824 =  x_423 & ~n_1822;
assign n_1825 = ~n_1823 & ~n_1824;
assign n_1826 = ~n_839 & ~n_1825;
assign n_1827 = ~n_1820 & ~n_1826;
assign n_1828 =  x_423 & ~n_1827;
assign n_1829 = ~x_423 &  n_1827;
assign n_1830 = ~n_1828 & ~n_1829;
assign n_1831 =  x_307 & ~x_323;
assign n_1832 =  x_422 &  n_1823;
assign n_1833 = ~x_422 & ~n_1823;
assign n_1834 = ~n_839 & ~n_1833;
assign n_1835 = ~n_1832 &  n_1834;
assign n_1836 = ~n_1831 & ~n_1835;
assign n_1837 =  x_422 & ~n_1836;
assign n_1838 = ~x_422 &  n_1836;
assign n_1839 = ~n_1837 & ~n_1838;
assign n_1840 =  x_307 &  x_347;
assign n_1841 =  x_421 & ~n_213;
assign n_1842 = ~i_162 &  x_214;
assign n_1843 =  n_838 & ~n_1842;
assign n_1844 = ~n_1841 & ~n_1843;
assign n_1845 = ~n_8 & ~n_1844;
assign n_1846 = ~x_421 & ~n_1821;
assign n_1847 = ~n_1845 & ~n_1846;
assign n_1848 = ~x_307 & ~n_1847;
assign n_1849 = ~n_1840 & ~n_1848;
assign n_1850 =  x_421 &  n_1849;
assign n_1851 = ~x_421 & ~n_1849;
assign n_1852 = ~n_1850 & ~n_1851;
assign n_1853 = ~n_213 &  n_35;
assign n_1854 = ~i_159 &  x_214;
assign n_1855 =  n_838 & ~n_1854;
assign n_1856 = ~n_8 & ~n_1855;
assign n_1857 = ~n_1853 &  n_1856;
assign n_1858 = ~n_8 & ~n_1857;
assign n_1859 =  x_420 & ~n_1858;
assign n_1860 = ~x_304 &  n_1857;
assign n_1861 = ~n_1859 & ~n_1860;
assign n_1862 = ~x_307 & ~n_1861;
assign n_1863 =  x_307 & ~x_346;
assign n_1864 = ~n_1862 & ~n_1863;
assign n_1865 =  x_420 & ~n_1864;
assign n_1866 = ~x_420 &  n_1864;
assign n_1867 = ~n_1865 & ~n_1866;
assign n_1868 =  x_419 & ~n_831;
assign n_1869 = ~x_419 &  n_831;
assign n_1870 = ~n_1868 & ~n_1869;
assign n_1871 =  x_418 &  n_959;
assign n_1872 = ~x_418 & ~n_959;
assign n_1873 = ~n_1871 & ~n_1872;
assign n_1874 =  x_417 &  n_3;
assign n_1875 = ~x_417 & ~n_3;
assign n_1876 = ~n_1874 & ~n_1875;
assign n_1877 = ~x_228 &  n_5;
assign n_1878 =  n_1877 & ~n_98;
assign n_1879 =  x_416 & ~n_1878;
assign n_1880 = ~x_416 &  n_1878;
assign n_1881 = ~n_1879 & ~n_1880;
assign n_1882 = ~x_228 & ~n_812;
assign n_1883 =  n_6 &  n_1882;
assign n_1884 =  n_733 &  n_1883;
assign n_1885 = ~x_305 & ~x_311;
assign n_1886 = ~n_3 &  n_1885;
assign n_1887 =  x_415 &  n_1886;
assign n_1888 =  i_169 &  x_311;
assign n_1889 =  n_213 & ~n_1888;
assign n_1890 = ~n_1887 &  n_1889;
assign n_1891 =  n_239 & ~n_1890;
assign n_1892 = ~n_1884 & ~n_1891;
assign n_1893 =  x_415 & ~n_1892;
assign n_1894 = ~x_415 &  n_1892;
assign n_1895 = ~n_1893 & ~n_1894;
assign n_1896 =  x_352 &  n_283;
assign n_1897 = ~n_361 &  n_1896;
assign n_1898 =  x_414 &  n_1897;
assign n_1899 = ~x_414 & ~n_1897;
assign n_1900 = ~n_1898 & ~n_1899;
assign n_1901 =  x_354 &  n_283;
assign n_1902 = ~n_337 &  n_1901;
assign n_1903 =  x_413 &  n_1902;
assign n_1904 = ~x_413 & ~n_1902;
assign n_1905 = ~n_1903 & ~n_1904;
assign n_1906 =  x_353 &  n_283;
assign n_1907 = ~n_349 &  n_1906;
assign n_1908 =  x_412 &  n_1907;
assign n_1909 = ~x_412 & ~n_1907;
assign n_1910 = ~n_1908 & ~n_1909;
assign n_1911 =  x_358 &  n_283;
assign n_1912 = ~n_289 &  n_1911;
assign n_1913 =  x_411 &  n_1912;
assign n_1914 = ~x_411 & ~n_1912;
assign n_1915 = ~n_1913 & ~n_1914;
assign n_1916 =  x_357 &  n_283;
assign n_1917 = ~n_301 &  n_1916;
assign n_1918 =  x_410 &  n_1917;
assign n_1919 = ~x_410 & ~n_1917;
assign n_1920 = ~n_1918 & ~n_1919;
assign n_1921 =  x_356 &  n_283;
assign n_1922 = ~n_313 &  n_1921;
assign n_1923 =  x_409 &  n_1922;
assign n_1924 = ~x_409 & ~n_1922;
assign n_1925 = ~n_1923 & ~n_1924;
assign n_1926 =  x_355 &  n_283;
assign n_1927 = ~n_325 &  n_1926;
assign n_1928 =  x_408 &  n_1927;
assign n_1929 = ~x_408 & ~n_1927;
assign n_1930 = ~n_1928 & ~n_1929;
assign n_1931 =  x_407 &  n_8;
assign n_1932 = ~n_9 & ~n_1931;
assign n_1933 = ~x_228 & ~n_1932;
assign n_1934 =  x_407 &  n_1933;
assign n_1935 = ~x_407 & ~n_1933;
assign n_1936 = ~n_1934 & ~n_1935;
assign n_1937 =  x_406 & ~n_1;
assign n_1938 =  x_310 &  n_4;
assign n_1939 =  i_154 &  n_1938;
assign n_1940 = ~n_1937 & ~n_1939;
assign n_1941 =  n_119 & ~n_1940;
assign n_1942 =  x_406 &  n_1941;
assign n_1943 = ~x_406 & ~n_1941;
assign n_1944 = ~n_1942 & ~n_1943;
assign n_1945 = ~x_232 &  x_405;
assign n_1946 = ~x_227 & ~n_1945;
assign n_1947 = ~x_337 & ~n_1946;
assign n_1948 =  x_405 &  n_1947;
assign n_1949 = ~x_405 & ~n_1947;
assign n_1950 = ~n_1948 & ~n_1949;
assign n_1951 = ~n_8 &  n_725;
assign n_1952 =  x_391 &  n_1951;
assign n_1953 = ~i_186 & ~x_390;
assign n_1954 =  x_411 & ~n_1953;
assign n_1955 = ~x_358 & ~n_1954;
assign n_1956 = ~n_290 &  n_1955;
assign n_1957 = ~n_1952 &  n_1956;
assign n_1958 =  x_404 &  n_1957;
assign n_1959 = ~x_404 & ~n_1957;
assign n_1960 = ~n_1958 & ~n_1959;
assign n_1961 = ~i_187 & ~x_387;
assign n_1962 =  x_408 & ~n_1961;
assign n_1963 = ~x_355 & ~n_1962;
assign n_1964 = ~n_326 &  n_1963;
assign n_1965 = ~n_1952 &  n_1964;
assign n_1966 =  x_403 &  n_1965;
assign n_1967 = ~x_403 & ~n_1965;
assign n_1968 = ~n_1966 & ~n_1967;
assign n_1969 =  x_305 & ~n_834;
assign n_1970 =  x_402 &  n_1969;
assign n_1971 = ~x_402 & ~n_1969;
assign n_1972 = ~n_1970 & ~n_1971;
assign n_1973 =  x_401 &  n_1886;
assign n_1974 =  i_192 &  x_311;
assign n_1975 = ~n_1973 & ~n_1974;
assign n_1976 =  n_239 & ~n_1975;
assign n_1977 =  n_390 &  n_1883;
assign n_1978 = ~n_1976 & ~n_1977;
assign n_1979 =  x_401 & ~n_1978;
assign n_1980 = ~x_401 &  n_1978;
assign n_1981 = ~n_1979 & ~n_1980;
assign n_1982 =  x_349 &  n_1938;
assign n_1983 =  i_181 & ~x_394;
assign n_1984 = ~i_181 & ~x_398;
assign n_1985 = ~i_183 & ~n_1984;
assign n_1986 = ~n_1983 &  n_1985;
assign n_1987 =  i_181 & ~x_392;
assign n_1988 = ~i_181 & ~x_399;
assign n_1989 =  i_183 & ~n_1988;
assign n_1990 = ~n_1987 &  n_1989;
assign n_1991 =  i_182 & ~n_1990;
assign n_1992 = ~n_1986 &  n_1991;
assign n_1993 =  i_181 & ~x_393;
assign n_1994 = ~i_181 & ~x_397;
assign n_1995 =  i_183 & ~n_1994;
assign n_1996 = ~n_1993 &  n_1995;
assign n_1997 =  i_181 & ~x_396;
assign n_1998 = ~i_181 & ~x_395;
assign n_1999 = ~i_183 & ~n_1998;
assign n_2000 = ~n_1997 &  n_1999;
assign n_2001 = ~i_182 & ~n_2000;
assign n_2002 = ~n_1996 &  n_2001;
assign n_2003 =  i_154 & ~n_2002;
assign n_2004 = ~n_1992 &  n_2003;
assign n_2005 =  x_399 &  n_867;
assign n_2006 =  x_396 &  n_880;
assign n_2007 = ~n_2005 & ~n_2006;
assign n_2008 =  x_394 &  n_871;
assign n_2009 =  x_397 &  n_885;
assign n_2010 = ~n_2008 & ~n_2009;
assign n_2011 =  n_2007 &  n_2010;
assign n_2012 =  x_392 &  n_873;
assign n_2013 =  x_393 &  n_864;
assign n_2014 = ~n_2012 & ~n_2013;
assign n_2015 =  x_395 &  n_883;
assign n_2016 =  x_398 &  n_877;
assign n_2017 = ~n_2015 & ~n_2016;
assign n_2018 =  n_2014 &  n_2017;
assign n_2019 =  n_2011 &  n_2018;
assign n_2020 = ~n_2004 &  n_2019;
assign n_2021 =  n_1982 & ~n_2020;
assign n_2022 = ~i_180 &  n_873;
assign n_2023 = ~x_404 &  n_867;
assign n_2024 = ~n_2022 & ~n_2023;
assign n_2025 = ~i_197 &  n_864;
assign n_2026 = ~i_196 &  n_883;
assign n_2027 = ~n_2025 & ~n_2026;
assign n_2028 =  n_2024 &  n_2027;
assign n_2029 = ~i_195 &  n_871;
assign n_2030 = ~i_194 &  n_877;
assign n_2031 = ~n_2029 & ~n_2030;
assign n_2032 = ~x_403 &  n_880;
assign n_2033 = ~i_193 &  n_885;
assign n_2034 = ~n_2032 & ~n_2033;
assign n_2035 =  n_2031 &  n_2034;
assign n_2036 =  n_2028 &  n_2035;
assign n_2037 =  n_921 & ~n_2036;
assign n_2038 = ~x_305 & ~x_310;
assign n_2039 = ~x_406 & ~x_407;
assign n_2040 =  n_2038 &  n_2039;
assign n_2041 =  i_15 & ~x_262;
assign n_2042 = ~n_2040 &  n_2041;
assign n_2043 =  x_258 & ~n_438;
assign n_2044 = ~x_337 &  n_1945;
assign n_2045 = ~x_265 & ~x_299;
assign n_2046 = ~n_2044 &  n_2045;
assign n_2047 = ~n_2043 &  n_2046;
assign n_2048 = ~n_2042 &  n_2047;
assign n_2049 = ~n_2037 &  n_2048;
assign n_2050 = ~n_2021 &  n_2049;
assign n_2051 =  x_400 & ~n_2050;
assign n_2052 = ~x_400 &  n_2050;
assign n_2053 = ~n_2051 & ~n_2052;
assign n_2054 =  n_1877 &  n_97;
assign n_2055 = ~x_242 &  x_250;
assign n_2056 =  n_104 &  n_2055;
assign n_2057 = ~n_5 &  n_2056;
assign n_2058 = ~n_2054 & ~n_2057;
assign n_2059 =  x_271 & ~n_2058;
assign n_2060 = ~x_271 &  n_2058;
assign n_2061 = ~n_2059 & ~n_2060;
assign n_2062 =  x_270 &  n_958;
assign n_2063 = ~x_270 & ~n_958;
assign n_2064 = ~n_2062 & ~n_2063;
assign n_2065 =  x_269 & ~n_1;
assign n_2066 = ~n_2065 & ~n_921;
assign n_2067 =  n_119 & ~n_2066;
assign n_2068 =  x_269 &  n_2067;
assign n_2069 = ~x_269 & ~n_2067;
assign n_2070 = ~n_2068 & ~n_2069;
assign n_2071 = ~x_400 & ~x_415;
assign n_2072 = ~i_68 & ~x_269;
assign n_2073 =  x_400 &  n_2072;
assign n_2074 = ~n_2071 & ~n_2073;
assign n_2075 =  x_268 &  n_2074;
assign n_2076 = ~x_268 & ~n_2074;
assign n_2077 = ~n_2075 & ~n_2076;
assign n_2078 =  x_267 &  n_440;
assign n_2079 = ~x_267 & ~n_440;
assign n_2080 = ~n_2078 & ~n_2079;
assign n_2081 =  x_266 & ~n_998;
assign n_2082 =  x_349 &  n_889;
assign n_2083 = ~x_349 & ~x_383;
assign n_2084 =  n_998 & ~n_2083;
assign n_2085 = ~n_2082 &  n_2084;
assign n_2086 = ~n_2081 & ~n_2085;
assign n_2087 =  x_266 & ~n_2086;
assign n_2088 = ~x_266 &  n_2086;
assign n_2089 = ~n_2087 & ~n_2088;
assign n_2090 =  x_265 &  n_2043;
assign n_2091 = ~x_265 & ~n_2043;
assign n_2092 = ~n_2090 & ~n_2091;
assign n_2093 =  x_264 &  x_400;
assign n_2094 = ~x_283 & ~x_303;
assign n_2095 =  n_1982 &  n_2094;
assign n_2096 = ~n_2093 & ~n_2095;
assign n_2097 =  n_119 & ~n_2096;
assign n_2098 =  x_264 &  n_2097;
assign n_2099 = ~x_264 & ~n_2097;
assign n_2100 = ~n_2098 & ~n_2099;
assign n_2101 =  x_263 & ~n_1;
assign n_2102 = ~x_263 &  n_1;
assign n_2103 = ~n_2101 & ~n_2102;
assign n_2104 =  x_262 & ~n_119;
assign n_2105 = ~x_262 &  n_119;
assign n_2106 = ~n_2104 & ~n_2105;
assign n_2107 =  x_261 &  x_342;
assign n_2108 = ~x_261 & ~x_342;
assign n_2109 = ~n_2107 & ~n_2108;
assign n_2110 =  x_260 &  x_340;
assign n_2111 = ~x_260 & ~x_340;
assign n_2112 = ~n_2110 & ~n_2111;
assign n_2113 =  x_259 &  x_339;
assign n_2114 = ~x_259 & ~x_339;
assign n_2115 = ~n_2113 & ~n_2114;
assign n_2116 =  x_258 &  x_337;
assign n_2117 = ~x_258 & ~x_337;
assign n_2118 = ~n_2116 & ~n_2117;
assign n_2119 =  x_257 &  x_336;
assign n_2120 = ~n_495 & ~n_2119;
assign n_2121 =  x_256 &  x_334;
assign n_2122 = ~x_256 & ~x_334;
assign n_2123 = ~n_2121 & ~n_2122;
assign n_2124 =  x_255 &  x_333;
assign n_2125 = ~x_255 & ~x_333;
assign n_2126 = ~n_2124 & ~n_2125;
assign n_2127 =  x_254 &  x_332;
assign n_2128 = ~x_254 & ~x_332;
assign n_2129 = ~n_2127 & ~n_2128;
assign n_2130 =  x_253 &  x_331;
assign n_2131 = ~x_253 & ~x_331;
assign n_2132 = ~n_2130 & ~n_2131;
assign n_2133 =  x_252 &  x_330;
assign n_2134 = ~x_252 & ~x_330;
assign n_2135 = ~n_2133 & ~n_2134;
assign n_2136 =  x_251 &  x_329;
assign n_2137 = ~x_251 & ~x_329;
assign n_2138 = ~n_2136 & ~n_2137;
assign n_2139 =  x_250 &  x_328;
assign n_2140 = ~x_250 & ~x_328;
assign n_2141 = ~n_2139 & ~n_2140;
assign n_2142 = ~x_228 &  x_242;
assign n_2143 =  n_95 &  n_2142;
assign n_2144 =  x_249 &  n_2143;
assign n_2145 = ~x_249 & ~n_2143;
assign n_2146 = ~n_2144 & ~n_2145;
assign n_2147 =  x_248 &  x_321;
assign n_2148 = ~x_248 & ~x_321;
assign n_2149 = ~n_2147 & ~n_2148;
assign n_2150 =  x_247 &  x_320;
assign n_2151 = ~x_247 & ~x_320;
assign n_2152 = ~n_2150 & ~n_2151;
assign n_2153 =  x_246 &  x_305;
assign n_2154 = ~x_246 & ~x_305;
assign n_2155 = ~n_2153 & ~n_2154;
assign n_2156 =  x_245 &  n_1042;
assign n_2157 = ~x_245 & ~n_1042;
assign n_2158 = ~n_2156 & ~n_2157;
assign n_2159 =  x_244 &  x_262;
assign n_2160 = ~x_244 & ~x_262;
assign n_2161 = ~n_2159 & ~n_2160;
assign n_2162 =  x_243 &  x_259;
assign n_2163 = ~n_442 & ~n_2162;
assign n_2164 =  x_242 &  x_257;
assign n_2165 = ~x_242 & ~x_257;
assign n_2166 = ~n_2164 & ~n_2165;
assign n_2167 =  x_241 &  x_256;
assign n_2168 = ~x_241 & ~x_256;
assign n_2169 = ~n_2167 & ~n_2168;
assign n_2170 =  x_240 &  x_255;
assign n_2171 = ~x_240 & ~x_255;
assign n_2172 = ~n_2170 & ~n_2171;
assign n_2173 =  x_239 &  x_254;
assign n_2174 = ~x_239 & ~x_254;
assign n_2175 = ~n_2173 & ~n_2174;
assign n_2176 =  x_238 &  x_253;
assign n_2177 = ~x_238 & ~x_253;
assign n_2178 = ~n_2176 & ~n_2177;
assign n_2179 =  x_237 &  x_252;
assign n_2180 = ~x_237 & ~x_252;
assign n_2181 = ~n_2179 & ~n_2180;
assign n_2182 =  x_236 &  x_251;
assign n_2183 = ~x_236 & ~x_251;
assign n_2184 = ~n_2182 & ~n_2183;
assign n_2185 =  x_225 &  x_235;
assign n_2186 = ~x_225 & ~x_235;
assign n_2187 = ~n_2185 & ~n_2186;
assign n_2188 =  x_234 &  x_248;
assign n_2189 = ~x_234 & ~x_248;
assign n_2190 = ~n_2188 & ~n_2189;
assign n_2191 =  x_233 &  x_247;
assign n_2192 = ~x_233 & ~x_247;
assign n_2193 = ~n_2191 & ~n_2192;
assign n_2194 =  x_230 &  x_232;
assign n_2195 = ~x_230 & ~x_232;
assign n_2196 = ~n_2194 & ~n_2195;
assign n_2197 =  x_229 &  x_231;
assign n_2198 = ~x_229 & ~x_231;
assign n_2199 = ~n_2197 & ~n_2198;
assign n_2200 =  x_230 &  x_231;
assign n_2201 = ~n_445 & ~n_2200;
assign n_2202 =  x_229 &  x_243;
assign n_2203 = ~x_229 & ~x_243;
assign n_2204 = ~n_2202 & ~n_2203;
assign n_2205 =  x_228 &  x_232;
assign n_2206 = ~n_119 & ~n_2205;
assign n_2207 =  x_227 &  x_228;
assign n_2208 = ~x_227 & ~x_228;
assign n_2209 = ~n_2207 & ~n_2208;
assign n_2210 =  x_226 &  x_235;
assign n_2211 = ~n_1009 & ~n_2210;
assign n_2212 =  x_225 &  x_242;
assign n_2213 = ~n_494 & ~n_2212;
assign n_2214 =  x_224 &  x_234;
assign n_2215 = ~x_224 & ~x_234;
assign n_2216 = ~n_2214 & ~n_2215;
assign n_2217 =  x_223 &  x_224;
assign n_2218 = ~x_223 & ~x_224;
assign n_2219 = ~n_2217 & ~n_2218;
assign n_2220 =  x_222 &  x_223;
assign n_2221 = ~x_222 & ~x_223;
assign n_2222 = ~n_2220 & ~n_2221;
assign n_2223 =  x_221 &  x_222;
assign n_2224 = ~x_221 & ~x_222;
assign n_2225 = ~n_2223 & ~n_2224;
assign n_2226 =  x_220 &  x_233;
assign n_2227 = ~x_220 & ~x_233;
assign n_2228 = ~n_2226 & ~n_2227;
assign n_2229 =  x_219 &  x_220;
assign n_2230 = ~x_219 & ~x_220;
assign n_2231 = ~n_2229 & ~n_2230;
assign n_2232 =  x_218 &  x_219;
assign n_2233 = ~x_218 & ~x_219;
assign n_2234 = ~n_2232 & ~n_2233;
assign n_2235 =  x_216 &  x_217;
assign n_2236 = ~x_216 & ~x_217;
assign n_2237 = ~n_2235 & ~n_2236;
assign n_2238 =  x_215 &  x_216;
assign n_2239 = ~x_215 & ~x_216;
assign n_2240 = ~n_2238 & ~n_2239;
assign n_2241 =  i_5 &  x_215;
assign n_2242 = ~i_5 & ~x_215;
assign n_2243 = ~n_2241 & ~n_2242;
assign n_2244 = ~i_52 & ~n_1629;
assign n_2245 =  n_1647 &  n_1650;
assign n_2246 =  n_1630 & ~n_1651;
assign n_2247 = ~n_2245 &  n_2246;
assign n_2248 =  x_274 & ~n_1630;
assign n_2249 =  n_1629 & ~n_2248;
assign n_2250 = ~n_2247 &  n_2249;
assign n_2251 = ~n_2244 & ~n_2250;
assign n_2252 = ~n_1633 & ~n_2251;
assign n_2253 =  x_274 & ~n_1472;
assign n_2254 = ~n_1473 & ~n_2253;
assign n_2255 =  n_1633 &  n_2254;
assign n_2256 = ~n_2252 & ~n_2255;
assign n_2257 =  x_274 &  n_2256;
assign n_2258 = ~x_274 & ~n_2256;
assign n_2259 = ~n_2257 & ~n_2258;
assign n_2260 =  i_51 & ~n_1629;
assign n_2261 =  i_31 &  n_1010;
assign n_2262 =  i_38 & ~n_1010;
assign n_2263 = ~n_2261 & ~n_2262;
assign n_2264 =  n_1731 &  n_2263;
assign n_2265 = ~n_1731 & ~n_2263;
assign n_2266 =  n_1630 & ~n_2265;
assign n_2267 = ~n_2264 &  n_2266;
assign n_2268 = ~x_273 & ~n_1630;
assign n_2269 =  n_1629 & ~n_2268;
assign n_2270 = ~n_2267 &  n_2269;
assign n_2271 = ~n_2260 & ~n_2270;
assign n_2272 = ~n_1633 &  n_2271;
assign n_2273 =  x_273 & ~n_1692;
assign n_2274 = ~x_273 &  n_1692;
assign n_2275 = ~n_2273 & ~n_2274;
assign n_2276 =  n_1633 &  n_2275;
assign n_2277 = ~n_2272 & ~n_2276;
assign n_2278 =  x_273 &  n_2277;
assign n_2279 = ~x_273 & ~n_2277;
assign n_2280 = ~n_2278 & ~n_2279;
assign n_2281 =  i_55 &  x_249;
assign n_2282 =  x_272 & ~x_301;
assign n_2283 =  n_102 &  n_2282;
assign n_2284 = ~n_2281 &  n_2283;
assign n_2285 =  n_1626 &  n_2284;
assign n_2286 = ~n_1626 & ~n_1038;
assign n_2287 = ~n_1624 &  n_2286;
assign n_2288 = ~n_2285 & ~n_2287;
assign n_2289 =  x_272 & ~n_2288;
assign n_2290 = ~x_272 &  n_2288;
assign n_2291 = ~n_2289 & ~n_2290;
assign n_2292 =  x_279 & ~n_1010;
assign n_2293 = ~n_1661 &  n_1751;
assign n_2294 = ~n_2292 & ~n_2293;
assign n_2295 =  n_1672 & ~n_2294;
assign n_2296 =  x_279 &  n_1631;
assign n_2297 =  n_1758 &  n_1713;
assign n_2298 =  i_209 &  i_210;
assign n_2299 =  i_212 &  n_2298;
assign n_2300 = ~n_2297 & ~n_2299;
assign n_2301 = ~n_1629 & ~n_2300;
assign n_2302 = ~n_2296 & ~n_2301;
assign n_2303 = ~n_2295 &  n_2302;
assign n_2304 = ~n_1633 & ~n_2303;
assign n_2305 = ~n_1638 &  n_1766;
assign n_2306 =  n_1633 &  n_2305;
assign n_2307 = ~n_2304 & ~n_2306;
assign n_2308 =  x_279 & ~n_2307;
assign n_2309 = ~x_279 &  n_2307;
assign n_2310 = ~n_2308 & ~n_2309;
assign n_2311 =  n_285 &  n_1952;
assign n_2312 =  n_284 &  n_1951;
assign n_2313 =  x_358 &  x_399;
assign n_2314 = ~n_1951 &  n_2313;
assign n_2315 = ~n_2312 & ~n_2314;
assign n_2316 = ~n_2311 &  n_2315;
assign n_2317 =  x_399 & ~n_2316;
assign n_2318 = ~x_399 &  n_2316;
assign n_2319 = ~n_2317 & ~n_2318;
assign n_2320 =  n_297 &  n_1952;
assign n_2321 =  n_296 &  n_1951;
assign n_2322 =  x_357 &  x_398;
assign n_2323 = ~n_1951 &  n_2322;
assign n_2324 = ~n_2321 & ~n_2323;
assign n_2325 = ~n_2320 &  n_2324;
assign n_2326 =  x_398 & ~n_2325;
assign n_2327 = ~x_398 &  n_2325;
assign n_2328 = ~n_2326 & ~n_2327;
assign n_2329 =  n_309 &  n_1952;
assign n_2330 =  n_308 &  n_1951;
assign n_2331 =  x_356 &  x_397;
assign n_2332 = ~n_1951 &  n_2331;
assign n_2333 = ~n_2330 & ~n_2332;
assign n_2334 = ~n_2329 &  n_2333;
assign n_2335 =  x_397 & ~n_2334;
assign n_2336 = ~x_397 &  n_2334;
assign n_2337 = ~n_2335 & ~n_2336;
assign n_2338 =  n_321 &  n_1952;
assign n_2339 =  n_320 &  n_1951;
assign n_2340 =  x_355 &  x_396;
assign n_2341 = ~n_1951 &  n_2340;
assign n_2342 = ~n_2339 & ~n_2341;
assign n_2343 = ~n_2338 &  n_2342;
assign n_2344 =  x_396 & ~n_2343;
assign n_2345 = ~x_396 &  n_2343;
assign n_2346 = ~n_2344 & ~n_2345;
assign n_2347 =  n_333 &  n_1952;
assign n_2348 =  n_332 &  n_1951;
assign n_2349 =  x_354 &  x_395;
assign n_2350 = ~n_1951 &  n_2349;
assign n_2351 = ~n_2348 & ~n_2350;
assign n_2352 = ~n_2347 &  n_2351;
assign n_2353 =  x_395 & ~n_2352;
assign n_2354 = ~x_395 &  n_2352;
assign n_2355 = ~n_2353 & ~n_2354;
assign n_2356 =  n_345 &  n_1952;
assign n_2357 =  n_344 &  n_1951;
assign n_2358 =  x_353 &  x_394;
assign n_2359 = ~n_1951 &  n_2358;
assign n_2360 = ~n_2357 & ~n_2359;
assign n_2361 = ~n_2356 &  n_2360;
assign n_2362 =  x_394 & ~n_2361;
assign n_2363 = ~x_394 &  n_2361;
assign n_2364 = ~n_2362 & ~n_2363;
assign n_2365 =  n_357 &  n_1952;
assign n_2366 =  n_356 &  n_1951;
assign n_2367 =  x_352 &  x_393;
assign n_2368 = ~n_1951 &  n_2367;
assign n_2369 = ~n_2366 & ~n_2368;
assign n_2370 = ~n_2365 &  n_2369;
assign n_2371 =  x_393 & ~n_2370;
assign n_2372 = ~x_393 &  n_2370;
assign n_2373 = ~n_2371 & ~n_2372;
assign n_2374 =  n_371 &  n_1952;
assign n_2375 =  n_369 &  n_1951;
assign n_2376 = ~i_184 & ~x_383;
assign n_2377 =  x_351 & ~n_2376;
assign n_2378 = ~n_1951 &  n_2377;
assign n_2379 = ~n_2375 & ~n_2378;
assign n_2380 = ~n_2374 &  n_2379;
assign n_2381 =  x_392 & ~n_2380;
assign n_2382 = ~x_392 &  n_2380;
assign n_2383 = ~n_2381 & ~n_2382;
assign n_2384 =  x_391 &  n_8;
assign n_2385 = ~x_364 & ~n_2384;
assign n_2386 =  x_391 & ~n_2385;
assign n_2387 = ~x_391 &  n_2385;
assign n_2388 = ~n_2386 & ~n_2387;
assign n_2389 =  x_390 & ~n_290;
assign n_2390 = ~n_2389 & ~n_2312;
assign n_2391 =  x_390 & ~n_2390;
assign n_2392 = ~x_390 &  n_2390;
assign n_2393 = ~n_2391 & ~n_2392;
assign n_2394 =  x_389 & ~n_302;
assign n_2395 = ~n_2394 & ~n_2321;
assign n_2396 =  x_389 & ~n_2395;
assign n_2397 = ~x_389 &  n_2395;
assign n_2398 = ~n_2396 & ~n_2397;
assign n_2399 =  x_388 & ~n_314;
assign n_2400 = ~n_2399 & ~n_2330;
assign n_2401 =  x_388 & ~n_2400;
assign n_2402 = ~x_388 &  n_2400;
assign n_2403 = ~n_2401 & ~n_2402;
assign n_2404 =  x_387 & ~n_326;
assign n_2405 = ~n_2404 & ~n_2339;
assign n_2406 =  x_387 & ~n_2405;
assign n_2407 = ~x_387 &  n_2405;
assign n_2408 = ~n_2406 & ~n_2407;
assign n_2409 =  x_386 & ~n_338;
assign n_2410 = ~n_2409 & ~n_2348;
assign n_2411 =  x_386 & ~n_2410;
assign n_2412 = ~x_386 &  n_2410;
assign n_2413 = ~n_2411 & ~n_2412;
assign n_2414 =  x_385 & ~n_350;
assign n_2415 = ~n_2414 & ~n_2357;
assign n_2416 =  x_385 & ~n_2415;
assign n_2417 = ~x_385 &  n_2415;
assign n_2418 = ~n_2416 & ~n_2417;
assign n_2419 =  x_384 & ~n_362;
assign n_2420 = ~n_2419 & ~n_2366;
assign n_2421 =  x_384 & ~n_2420;
assign n_2422 = ~x_384 &  n_2420;
assign n_2423 = ~n_2421 & ~n_2422;
assign n_2424 =  x_383 & ~n_377;
assign n_2425 = ~n_2424 & ~n_2375;
assign n_2426 =  x_383 & ~n_2425;
assign n_2427 = ~x_383 &  n_2425;
assign n_2428 = ~n_2426 & ~n_2427;
assign n_2429 =  i_13 & ~x_325;
assign n_2430 =  i_167 &  x_325;
assign n_2431 = ~n_2429 & ~n_2430;
assign n_2432 =  n_4 &  n_2431;
assign n_2433 =  x_214 & ~x_382;
assign n_2434 = ~n_4 &  n_2433;
assign n_2435 = ~n_2432 & ~n_2434;
assign n_2436 =  x_382 &  n_2435;
assign n_2437 = ~x_382 & ~n_2435;
assign n_2438 = ~n_2436 & ~n_2437;
assign n_2439 =  i_12 & ~x_325;
assign n_2440 =  i_166 &  x_325;
assign n_2441 = ~n_2439 & ~n_2440;
assign n_2442 =  n_4 &  n_2441;
assign n_2443 =  x_214 & ~x_381;
assign n_2444 = ~n_4 &  n_2443;
assign n_2445 = ~n_2442 & ~n_2444;
assign n_2446 =  x_381 &  n_2445;
assign n_2447 = ~x_381 & ~n_2445;
assign n_2448 = ~n_2446 & ~n_2447;
assign n_2449 =  i_14 & ~x_325;
assign n_2450 =  i_168 &  x_325;
assign n_2451 = ~n_2449 & ~n_2450;
assign n_2452 =  n_4 &  n_2451;
assign n_2453 =  x_214 & ~x_380;
assign n_2454 = ~n_4 &  n_2453;
assign n_2455 = ~n_2452 & ~n_2454;
assign n_2456 =  x_380 &  n_2455;
assign n_2457 = ~x_380 & ~n_2455;
assign n_2458 = ~n_2456 & ~n_2457;
assign n_2459 = ~n_232 &  n_233;
assign n_2460 =  n_18 &  n_29;
assign n_2461 =  n_2459 & ~n_2460;
assign n_2462 = ~x_311 &  n_49;
assign n_2463 =  n_29 &  n_2462;
assign n_2464 =  n_2461 & ~n_2463;
assign n_2465 =  n_18 &  n_23;
assign n_2466 =  n_48 &  n_45;
assign n_2467 = ~n_2465 & ~n_2466;
assign n_2468 =  n_2464 &  n_2467;
assign n_2469 = ~n_368 &  n_11;
assign n_2470 = ~n_6 & ~n_2469;
assign n_2471 = ~n_2468 &  n_2470;
assign n_2472 =  x_379 & ~n_2471;
assign n_2473 = ~x_379 &  n_2471;
assign n_2474 = ~n_2472 & ~n_2473;
assign n_2475 =  n_5 & ~n_372;
assign n_2476 = ~i_9 & ~x_325;
assign n_2477 = ~i_157 &  x_325;
assign n_2478 = ~n_2476 & ~n_2477;
assign n_2479 = ~n_5 &  n_2478;
assign n_2480 = ~i_10 & ~x_325;
assign n_2481 = ~i_161 &  x_325;
assign n_2482 = ~n_2480 & ~n_2481;
assign n_2483 = ~i_11 & ~x_325;
assign n_2484 = ~i_164 &  x_325;
assign n_2485 = ~n_2483 & ~n_2484;
assign n_2486 =  n_2482 &  n_2485;
assign n_2487 =  n_2479 &  n_2486;
assign n_2488 = ~n_2475 & ~n_2487;
assign n_2489 =  x_378 & ~n_2488;
assign n_2490 = ~x_378 &  n_2488;
assign n_2491 = ~n_2489 & ~n_2490;
assign n_2492 =  x_377 &  n_12;
assign n_2493 =  n_2464 &  n_2465;
assign n_2494 = ~n_2492 & ~n_2493;
assign n_2495 =  x_377 & ~n_2494;
assign n_2496 = ~x_377 &  n_2494;
assign n_2497 = ~n_2495 & ~n_2496;
assign n_2498 =  x_376 &  n_12;
assign n_2499 = ~i_204 &  i_205;
assign n_2500 =  n_80 &  n_2499;
assign n_2501 =  n_250 &  n_2500;
assign n_2502 = ~n_249 & ~n_86;
assign n_2503 =  n_252 &  n_2502;
assign n_2504 = ~n_2501 &  n_2503;
assign n_2505 = ~i_204 & ~i_205;
assign n_2506 = ~i_207 &  n_2505;
assign n_2507 =  n_250 &  n_2506;
assign n_2508 =  n_2504 &  n_2507;
assign n_2509 = ~n_2498 & ~n_2508;
assign n_2510 =  x_376 & ~n_2509;
assign n_2511 = ~x_376 &  n_2509;
assign n_2512 = ~n_2510 & ~n_2511;
assign n_2513 =  x_375 &  n_5;
assign n_2514 = ~n_2478 &  n_2486;
assign n_2515 = ~n_5 &  n_2514;
assign n_2516 = ~n_2513 & ~n_2515;
assign n_2517 =  x_375 & ~n_2516;
assign n_2518 = ~x_375 &  n_2516;
assign n_2519 = ~n_2517 & ~n_2518;
assign n_2520 =  x_374 &  n_12;
assign n_2521 =  n_2461 &  n_2463;
assign n_2522 = ~n_2520 & ~n_2521;
assign n_2523 =  x_374 & ~n_2522;
assign n_2524 = ~x_374 &  n_2522;
assign n_2525 = ~n_2523 & ~n_2524;
assign n_2526 =  x_373 &  n_12;
assign n_2527 =  n_84 &  n_2500;
assign n_2528 =  n_2504 &  n_2527;
assign n_2529 = ~n_2526 & ~n_2528;
assign n_2530 =  x_373 & ~n_2529;
assign n_2531 = ~x_373 &  n_2529;
assign n_2532 = ~n_2530 & ~n_2531;
assign n_2533 =  x_372 &  n_5;
assign n_2534 =  n_2482 & ~n_2485;
assign n_2535 =  n_2479 &  n_2534;
assign n_2536 = ~n_2533 & ~n_2535;
assign n_2537 =  x_372 & ~n_2536;
assign n_2538 = ~x_372 &  n_2536;
assign n_2539 = ~n_2537 & ~n_2538;
assign n_2540 =  x_371 &  n_12;
assign n_2541 =  n_19 &  n_52;
assign n_2542 = ~n_2540 & ~n_2541;
assign n_2543 =  x_371 & ~n_2542;
assign n_2544 = ~x_371 &  n_2542;
assign n_2545 = ~n_2543 & ~n_2544;
assign n_2546 =  x_369 &  n_12;
assign n_2547 =  n_2501 &  n_2503;
assign n_2548 = ~n_2546 & ~n_2547;
assign n_2549 =  x_369 & ~n_2548;
assign n_2550 = ~x_369 &  n_2548;
assign n_2551 = ~n_2549 & ~n_2550;
assign n_2552 =  x_370 &  n_12;
assign n_2553 =  n_2459 &  n_2460;
assign n_2554 = ~n_2552 & ~n_2553;
assign n_2555 =  x_370 & ~n_2554;
assign n_2556 = ~x_370 &  n_2554;
assign n_2557 = ~n_2555 & ~n_2556;
assign n_2558 = ~n_2551 & ~n_2557;
assign n_2559 = ~n_2545 &  n_2558;
assign n_2560 = ~n_2539 &  n_2559;
assign n_2561 = ~n_2532 &  n_2560;
assign n_2562 = ~n_2525 &  n_2561;
assign n_2563 = ~n_2519 &  n_2562;
assign n_2564 = ~n_2512 &  n_2563;
assign n_2565 = ~n_2497 &  n_2564;
assign n_2566 = ~n_2491 &  n_2565;
assign n_2567 = ~n_2474 &  n_2566;
assign n_2568 = ~n_2458 &  n_2567;
assign n_2569 = ~n_2448 &  n_2568;
assign n_2570 = ~n_2438 &  n_2569;
assign n_2571 = ~n_2428 &  n_2570;
assign n_2572 = ~n_2423 &  n_2571;
assign n_2573 = ~n_2418 &  n_2572;
assign n_2574 = ~n_2413 &  n_2573;
assign n_2575 = ~n_2408 &  n_2574;
assign n_2576 = ~n_2403 &  n_2575;
assign n_2577 = ~n_2398 &  n_2576;
assign n_2578 = ~n_2393 &  n_2577;
assign n_2579 = ~n_2388 &  n_2578;
assign n_2580 = ~n_2383 &  n_2579;
assign n_2581 = ~n_2373 &  n_2580;
assign n_2582 = ~n_2364 &  n_2581;
assign n_2583 = ~n_2355 &  n_2582;
assign n_2584 = ~n_2346 &  n_2583;
assign n_2585 = ~n_2337 &  n_2584;
assign n_2586 = ~n_2328 &  n_2585;
assign n_2587 = ~n_2319 &  n_2586;
assign n_2588 =  x_214 &  n_2587;
assign n_2589 = ~n_2310 &  n_2588;
assign n_2590 = ~n_2291 &  n_2589;
assign n_2591 = ~n_2280 &  n_2590;
assign n_2592 = ~n_2259 &  n_2591;
assign n_2593 = ~n_2243 &  n_2592;
assign n_2594 = ~n_2240 &  n_2593;
assign n_2595 = ~n_2237 &  n_2594;
assign n_2596 = ~n_2234 &  n_2595;
assign n_2597 = ~n_2231 &  n_2596;
assign n_2598 = ~n_2228 &  n_2597;
assign n_2599 = ~n_2225 &  n_2598;
assign n_2600 = ~n_2222 &  n_2599;
assign n_2601 = ~n_2219 &  n_2600;
assign n_2602 = ~n_2216 &  n_2601;
assign n_2603 = ~n_2213 &  n_2602;
assign n_2604 = ~n_2211 &  n_2603;
assign n_2605 = ~n_2209 &  n_2604;
assign n_2606 = ~n_2206 &  n_2605;
assign n_2607 = ~n_2204 &  n_2606;
assign n_2608 = ~n_2201 &  n_2607;
assign n_2609 = ~n_2199 &  n_2608;
assign n_2610 = ~n_2196 &  n_2609;
assign n_2611 = ~n_2193 &  n_2610;
assign n_2612 = ~n_2190 &  n_2611;
assign n_2613 = ~n_2187 &  n_2612;
assign n_2614 = ~n_2184 &  n_2613;
assign n_2615 = ~n_2181 &  n_2614;
assign n_2616 = ~n_2178 &  n_2615;
assign n_2617 = ~n_2175 &  n_2616;
assign n_2618 = ~n_2172 &  n_2617;
assign n_2619 = ~n_2169 &  n_2618;
assign n_2620 = ~n_2166 &  n_2619;
assign n_2621 = ~n_2163 &  n_2620;
assign n_2622 = ~n_2161 &  n_2621;
assign n_2623 = ~n_2158 &  n_2622;
assign n_2624 = ~n_2155 &  n_2623;
assign n_2625 = ~n_2152 &  n_2624;
assign n_2626 = ~n_2149 &  n_2625;
assign n_2627 = ~n_2146 &  n_2626;
assign n_2628 = ~n_2141 &  n_2627;
assign n_2629 = ~n_2138 &  n_2628;
assign n_2630 = ~n_2135 &  n_2629;
assign n_2631 = ~n_2132 &  n_2630;
assign n_2632 = ~n_2129 &  n_2631;
assign n_2633 = ~n_2126 &  n_2632;
assign n_2634 = ~n_2123 &  n_2633;
assign n_2635 = ~n_2120 &  n_2634;
assign n_2636 = ~n_2118 &  n_2635;
assign n_2637 = ~n_2115 &  n_2636;
assign n_2638 = ~n_2112 &  n_2637;
assign n_2639 = ~n_2109 &  n_2638;
assign n_2640 = ~n_2106 &  n_2639;
assign n_2641 = ~n_2103 &  n_2640;
assign n_2642 = ~n_2100 &  n_2641;
assign n_2643 = ~n_2092 &  n_2642;
assign n_2644 = ~n_2089 &  n_2643;
assign n_2645 = ~n_2080 &  n_2644;
assign n_2646 = ~n_2077 &  n_2645;
assign n_2647 = ~n_2070 &  n_2646;
assign n_2648 = ~n_2064 &  n_2647;
assign n_2649 = ~n_2061 &  n_2648;
assign n_2650 = ~n_2053 &  n_2649;
assign n_2651 = ~n_1981 &  n_2650;
assign n_2652 = ~n_1972 &  n_2651;
assign n_2653 = ~n_1968 &  n_2652;
assign n_2654 = ~n_1960 &  n_2653;
assign n_2655 = ~n_1950 &  n_2654;
assign n_2656 = ~n_1944 &  n_2655;
assign n_2657 = ~n_1936 &  n_2656;
assign n_2658 = ~n_1930 &  n_2657;
assign n_2659 = ~n_1925 &  n_2658;
assign n_2660 = ~n_1920 &  n_2659;
assign n_2661 = ~n_1915 &  n_2660;
assign n_2662 = ~n_1910 &  n_2661;
assign n_2663 = ~n_1905 &  n_2662;
assign n_2664 = ~n_1900 &  n_2663;
assign n_2665 = ~n_1895 &  n_2664;
assign n_2666 = ~n_1881 &  n_2665;
assign n_2667 = ~n_1876 &  n_2666;
assign n_2668 = ~n_1873 &  n_2667;
assign n_2669 = ~n_1870 &  n_2668;
assign n_2670 = ~n_1867 &  n_2669;
assign n_2671 = ~n_1852 &  n_2670;
assign n_2672 = ~n_1839 &  n_2671;
assign n_2673 = ~n_1830 &  n_2672;
assign n_2674 = ~n_1819 &  n_2673;
assign n_2675 = ~n_1811 &  n_2674;
assign n_2676 = ~n_1798 &  n_2675;
assign n_2677 = ~n_1786 &  n_2676;
assign n_2678 = ~n_1771 &  n_2677;
assign n_2679 = ~n_1748 &  n_2678;
assign n_2680 = ~n_1727 &  n_2679;
assign n_2681 = ~n_1703 &  n_2680;
assign n_2682 = ~n_1671 &  n_2681;
assign n_2683 = ~n_1471 &  n_2682;
assign n_2684 = ~n_1468 &  n_2683;
assign n_2685 = ~n_1465 &  n_2684;
assign n_2686 = ~n_1455 &  n_2685;
assign n_2687 = ~n_1427 &  n_2686;
assign n_2688 = ~n_1374 &  n_2687;
assign n_2689 = ~n_1326 &  n_2688;
assign n_2690 = ~n_1213 &  n_2689;
assign n_2691 = ~n_1124 &  n_2690;
assign n_2692 = ~n_1114 &  n_2691;
assign n_2693 = ~n_1103 &  n_2692;
assign n_2694 = ~n_1093 &  n_2693;
assign n_2695 = ~n_1083 &  n_2694;
assign n_2696 = ~n_1049 &  n_2695;
assign n_2697 = ~n_1008 &  n_2696;
assign n_2698 = ~n_1004 &  n_2697;
assign n_2699 = ~n_996 &  n_2698;
assign n_2700 = ~n_973 &  n_2699;
assign n_2701 = ~n_965 &  n_2700;
assign n_2702 = ~n_927 &  n_2701;
assign n_2703 = ~n_862 &  n_2702;
assign n_2704 = ~n_857 &  n_2703;
assign n_2705 = ~n_854 &  n_2704;
assign n_2706 = ~n_836 &  n_2705;
assign n_2707 = ~n_833 &  n_2706;
assign n_2708 = ~n_828 &  n_2707;
assign n_2709 = ~n_825 &  n_2708;
assign n_2710 = ~n_819 &  n_2709;
assign n_2711 = ~n_809 &  n_2710;
assign n_2712 = ~n_803 &  n_2711;
assign n_2713 = ~n_796 &  n_2712;
assign n_2714 = ~n_790 &  n_2713;
assign n_2715 = ~n_784 &  n_2714;
assign n_2716 = ~n_778 &  n_2715;
assign n_2717 = ~n_774 &  n_2716;
assign n_2718 = ~n_770 &  n_2717;
assign n_2719 = ~n_766 &  n_2718;
assign n_2720 = ~n_762 &  n_2719;
assign n_2721 = ~n_759 &  n_2720;
assign n_2722 = ~n_752 &  n_2721;
assign n_2723 = ~n_745 &  n_2722;
assign n_2724 = ~n_739 &  n_2723;
assign n_2725 = ~n_732 &  n_2724;
assign n_2726 = ~n_724 &  n_2725;
assign n_2727 = ~n_720 &  n_2726;
assign n_2728 = ~n_716 &  n_2727;
assign n_2729 = ~n_713 &  n_2728;
assign n_2730 = ~n_703 &  n_2729;
assign n_2731 = ~n_682 &  n_2730;
assign n_2732 = ~n_650 &  n_2731;
assign n_2733 = ~n_606 &  n_2732;
assign n_2734 = ~n_561 &  n_2733;
assign n_2735 = ~n_503 &  n_2734;
assign n_2736 = ~n_500 &  n_2735;
assign n_2737 = ~n_468 &  n_2736;
assign n_2738 = ~n_465 &  n_2737;
assign n_2739 = ~n_462 &  n_2738;
assign n_2740 = ~n_452 &  n_2739;
assign n_2741 = ~n_436 &  n_2740;
assign n_2742 = ~n_432 &  n_2741;
assign n_2743 = ~n_429 &  n_2742;
assign n_2744 = ~n_423 &  n_2743;
assign n_2745 = ~n_418 &  n_2744;
assign n_2746 = ~n_412 &  n_2745;
assign n_2747 = ~n_406 &  n_2746;
assign n_2748 = ~n_400 &  n_2747;
assign n_2749 = ~n_394 &  n_2748;
assign n_2750 = ~n_386 &  n_2749;
assign n_2751 = ~n_381 &  n_2750;
assign n_2752 = ~n_366 &  n_2751;
assign n_2753 = ~n_354 &  n_2752;
assign n_2754 = ~n_342 &  n_2753;
assign n_2755 = ~n_330 &  n_2754;
assign n_2756 = ~n_318 &  n_2755;
assign n_2757 = ~n_306 &  n_2756;
assign n_2758 = ~n_294 &  n_2757;
assign n_2759 = ~n_281 &  n_2758;
assign n_2760 = ~n_271 &  n_2759;
assign n_2761 = ~n_257 &  n_2760;
assign n_2762 = ~n_246 &  n_2761;
assign n_2763 = ~n_238 &  n_2762;
assign n_2764 = ~n_230 &  n_2763;
assign n_2765 = ~n_118 &  n_2764;
assign n_2766 = ~n_91 &  n_2765;
assign n_2767 = ~n_67 &  n_2766;
assign n_2768 = ~n_61 &  n_2767;
assign o_1 = ~n_2768;
endmodule

