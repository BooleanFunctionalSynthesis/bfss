// Verilog file written by procedure writeCombinationalCircuitInVerilog
//Skolem functions to be generated for i_ variables
module pdtpmsmiim_all_bit_differing_from_cycle ( i_1, i_2, i_3, i_4, i_5, i_6, i_7, i_8, i_9, i_10, i_11, i_12, i_13, i_14, i_15, i_16, i_17, i_18, i_19, i_20, i_21, i_22, i_23, i_24, i_25, i_26, i_27, i_28, i_29, i_30, i_31, i_32, i_33, i_34, i_35, i_36, i_37, i_38, i_39, i_40, i_41, x_42, x_43, x_44, x_45, x_46, x_47, x_48, x_49, x_50, x_51, x_52, x_53, x_54, x_55, x_56, x_57, x_58, x_59, x_60, x_61, x_62, x_63, x_64, x_65, x_66, x_67, x_68, x_69, x_70, x_71, x_72, x_73, x_74, x_75, x_76, x_77, x_78, x_79, x_80, x_81, x_82, x_83, x_84, x_85, x_86, x_87, x_88, x_89, x_90, x_91, x_92, x_93, x_94, x_95, x_96, x_97, x_98, x_99, x_100, x_101, x_102, x_103, x_104, x_105, x_106, x_107, x_108, x_109, x_110, x_111, x_112, x_113, x_114, x_115, x_116, x_117, x_118, x_119, x_120, x_121, x_122, x_123, x_124, x_125, x_126, x_127, x_128, x_129, x_130, x_131, x_132, x_133, x_134, x_135, x_136, x_137, x_138, x_139, x_140, x_141, x_142, x_143, x_144, x_145, x_146, x_147, x_148, x_149, x_150, x_151, x_152, x_153, x_154, x_155, x_156, x_157, x_158, x_159, x_160, x_161, x_162, x_163, x_164, x_165, x_166, x_167, x_168, x_169, x_170, x_171, x_172, x_173, x_174, x_175, x_176, x_177, x_178, x_179, x_180, x_181, x_182, x_183, x_184, x_185, x_186, x_187, x_188, x_189, x_190, x_191, x_192, x_193, x_194, x_195, x_196, x_197, x_198, x_199, x_200, x_201, x_202, x_203, x_204, x_205, x_206, x_207, x_208, x_209, x_210, x_211, x_212, x_213, x_214, x_215, x_216, x_217, x_218, x_219, x_220, x_221, x_222, x_223, x_224, x_225, x_226, x_227, x_228, x_229, x_230, x_231, x_232, x_233, x_234, x_235, x_236, x_237, x_238, x_239, x_240, x_241, x_242, x_243, x_244, x_245, x_246, x_247, x_248, x_249, x_250, x_251, x_252, x_253, x_254, x_255, x_256, x_257, x_258, x_259, x_260, x_261, x_262, x_263, x_264, x_265, x_266, x_267, x_268, x_269, x_270, x_271, x_272, x_273, x_274, x_275, x_276, x_277, x_278, x_279, x_280, x_281, x_282, x_283, x_284, x_285, x_286, x_287, x_288, x_289, x_290, x_291, x_292, x_293, x_294, x_295, x_296, x_297, x_298, x_299, x_300, x_301, x_302, x_303, x_304, x_305, x_306, x_307, x_308, x_309, x_310, x_311, x_312, x_313, x_314, x_315, x_316, x_317, x_318, x_319, x_320, x_321, x_322, x_323, x_324, x_325, x_326, x_327, x_328, x_329, x_330, x_331, x_332, x_333, x_334, x_335, x_336, x_337, x_338, x_339, x_340, x_341, x_342, x_343, x_344, x_345, x_346, x_347, x_348, x_349, x_350, x_351, x_352, x_353, x_354, x_355, x_356, x_357, x_358, x_359, x_360, x_361, x_362, x_363, x_364, x_365, x_366, x_367, x_368, x_369, x_370, x_371, x_372, x_373, x_374, x_375, x_376, x_377, x_378, x_379, x_380, x_381, x_382, x_383, x_384, x_385, x_386, x_387, x_388, x_389, x_390, x_391, x_392, x_393, x_394, x_395, x_396, x_397, x_398, x_399, x_400, x_401, x_402, x_403, x_404, x_405, x_406, x_407, x_408, x_409, x_410, x_411, x_412, x_413, x_414, x_415, x_416, x_417, x_418, x_419, x_420, x_421, x_422, x_423, x_424, x_425, x_426, x_427, x_428, x_429, x_430, x_431, x_432, x_433, x_434, x_435, x_436, x_437, x_438, x_439, x_440, x_441, x_442, x_443, x_444, x_445, x_446, x_447, x_448, x_449, x_450, x_451, x_452, x_453, x_454, x_455, x_456, x_457, x_458, x_459, o_1 );
input i_1;
input i_2;
input i_3;
input i_4;
input i_5;
input i_6;
input i_7;
input i_8;
input i_9;
input i_10;
input i_11;
input i_12;
input i_13;
input i_14;
input i_15;
input i_16;
input i_17;
input i_18;
input i_19;
input i_20;
input i_21;
input i_22;
input i_23;
input i_24;
input i_25;
input i_26;
input i_27;
input i_28;
input i_29;
input i_30;
input i_31;
input i_32;
input i_33;
input i_34;
input i_35;
input i_36;
input i_37;
input i_38;
input i_39;
input i_40;
input i_41;
input x_42;
input x_43;
input x_44;
input x_45;
input x_46;
input x_47;
input x_48;
input x_49;
input x_50;
input x_51;
input x_52;
input x_53;
input x_54;
input x_55;
input x_56;
input x_57;
input x_58;
input x_59;
input x_60;
input x_61;
input x_62;
input x_63;
input x_64;
input x_65;
input x_66;
input x_67;
input x_68;
input x_69;
input x_70;
input x_71;
input x_72;
input x_73;
input x_74;
input x_75;
input x_76;
input x_77;
input x_78;
input x_79;
input x_80;
input x_81;
input x_82;
input x_83;
input x_84;
input x_85;
input x_86;
input x_87;
input x_88;
input x_89;
input x_90;
input x_91;
input x_92;
input x_93;
input x_94;
input x_95;
input x_96;
input x_97;
input x_98;
input x_99;
input x_100;
input x_101;
input x_102;
input x_103;
input x_104;
input x_105;
input x_106;
input x_107;
input x_108;
input x_109;
input x_110;
input x_111;
input x_112;
input x_113;
input x_114;
input x_115;
input x_116;
input x_117;
input x_118;
input x_119;
input x_120;
input x_121;
input x_122;
input x_123;
input x_124;
input x_125;
input x_126;
input x_127;
input x_128;
input x_129;
input x_130;
input x_131;
input x_132;
input x_133;
input x_134;
input x_135;
input x_136;
input x_137;
input x_138;
input x_139;
input x_140;
input x_141;
input x_142;
input x_143;
input x_144;
input x_145;
input x_146;
input x_147;
input x_148;
input x_149;
input x_150;
input x_151;
input x_152;
input x_153;
input x_154;
input x_155;
input x_156;
input x_157;
input x_158;
input x_159;
input x_160;
input x_161;
input x_162;
input x_163;
input x_164;
input x_165;
input x_166;
input x_167;
input x_168;
input x_169;
input x_170;
input x_171;
input x_172;
input x_173;
input x_174;
input x_175;
input x_176;
input x_177;
input x_178;
input x_179;
input x_180;
input x_181;
input x_182;
input x_183;
input x_184;
input x_185;
input x_186;
input x_187;
input x_188;
input x_189;
input x_190;
input x_191;
input x_192;
input x_193;
input x_194;
input x_195;
input x_196;
input x_197;
input x_198;
input x_199;
input x_200;
input x_201;
input x_202;
input x_203;
input x_204;
input x_205;
input x_206;
input x_207;
input x_208;
input x_209;
input x_210;
input x_211;
input x_212;
input x_213;
input x_214;
input x_215;
input x_216;
input x_217;
input x_218;
input x_219;
input x_220;
input x_221;
input x_222;
input x_223;
input x_224;
input x_225;
input x_226;
input x_227;
input x_228;
input x_229;
input x_230;
input x_231;
input x_232;
input x_233;
input x_234;
input x_235;
input x_236;
input x_237;
input x_238;
input x_239;
input x_240;
input x_241;
input x_242;
input x_243;
input x_244;
input x_245;
input x_246;
input x_247;
input x_248;
input x_249;
input x_250;
input x_251;
input x_252;
input x_253;
input x_254;
input x_255;
input x_256;
input x_257;
input x_258;
input x_259;
input x_260;
input x_261;
input x_262;
input x_263;
input x_264;
input x_265;
input x_266;
input x_267;
input x_268;
input x_269;
input x_270;
input x_271;
input x_272;
input x_273;
input x_274;
input x_275;
input x_276;
input x_277;
input x_278;
input x_279;
input x_280;
input x_281;
input x_282;
input x_283;
input x_284;
input x_285;
input x_286;
input x_287;
input x_288;
input x_289;
input x_290;
input x_291;
input x_292;
input x_293;
input x_294;
input x_295;
input x_296;
input x_297;
input x_298;
input x_299;
input x_300;
input x_301;
input x_302;
input x_303;
input x_304;
input x_305;
input x_306;
input x_307;
input x_308;
input x_309;
input x_310;
input x_311;
input x_312;
input x_313;
input x_314;
input x_315;
input x_316;
input x_317;
input x_318;
input x_319;
input x_320;
input x_321;
input x_322;
input x_323;
input x_324;
input x_325;
input x_326;
input x_327;
input x_328;
input x_329;
input x_330;
input x_331;
input x_332;
input x_333;
input x_334;
input x_335;
input x_336;
input x_337;
input x_338;
input x_339;
input x_340;
input x_341;
input x_342;
input x_343;
input x_344;
input x_345;
input x_346;
input x_347;
input x_348;
input x_349;
input x_350;
input x_351;
input x_352;
input x_353;
input x_354;
input x_355;
input x_356;
input x_357;
input x_358;
input x_359;
input x_360;
input x_361;
input x_362;
input x_363;
input x_364;
input x_365;
input x_366;
input x_367;
input x_368;
input x_369;
input x_370;
input x_371;
input x_372;
input x_373;
input x_374;
input x_375;
input x_376;
input x_377;
input x_378;
input x_379;
input x_380;
input x_381;
input x_382;
input x_383;
input x_384;
input x_385;
input x_386;
input x_387;
input x_388;
input x_389;
input x_390;
input x_391;
input x_392;
input x_393;
input x_394;
input x_395;
input x_396;
input x_397;
input x_398;
input x_399;
input x_400;
input x_401;
input x_402;
input x_403;
input x_404;
input x_405;
input x_406;
input x_407;
input x_408;
input x_409;
input x_410;
input x_411;
input x_412;
input x_413;
input x_414;
input x_415;
input x_416;
input x_417;
input x_418;
input x_419;
input x_420;
input x_421;
input x_422;
input x_423;
input x_424;
input x_425;
input x_426;
input x_427;
input x_428;
input x_429;
input x_430;
input x_431;
input x_432;
input x_433;
input x_434;
input x_435;
input x_436;
input x_437;
input x_438;
input x_439;
input x_440;
input x_441;
input x_442;
input x_443;
input x_444;
input x_445;
input x_446;
input x_447;
input x_448;
input x_449;
input x_450;
input x_451;
input x_452;
input x_453;
input x_454;
input x_455;
input x_456;
input x_457;
input x_458;
input x_459;
output o_1;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_12;
wire n_13;
wire n_14;
wire n_15;
wire n_16;
wire n_17;
wire n_18;
wire n_19;
wire n_20;
wire n_21;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_27;
wire n_28;
wire n_29;
wire n_30;
wire n_31;
wire n_32;
wire n_33;
wire n_34;
wire n_35;
wire n_36;
wire n_37;
wire n_38;
wire n_39;
wire n_40;
wire n_41;
wire n_42;
wire n_43;
wire n_44;
wire n_45;
wire n_46;
wire n_47;
wire n_48;
wire n_49;
wire n_50;
wire n_51;
wire n_52;
wire n_53;
wire n_54;
wire n_55;
wire n_56;
wire n_57;
wire n_58;
wire n_59;
wire n_60;
wire n_61;
wire n_62;
wire n_63;
wire n_64;
wire n_65;
wire n_66;
wire n_67;
wire n_68;
wire n_69;
wire n_70;
wire n_71;
wire n_72;
wire n_73;
wire n_74;
wire n_75;
wire n_76;
wire n_77;
wire n_78;
wire n_79;
wire n_80;
wire n_81;
wire n_82;
wire n_83;
wire n_84;
wire n_85;
wire n_86;
wire n_87;
wire n_88;
wire n_89;
wire n_90;
wire n_91;
wire n_92;
wire n_93;
wire n_94;
wire n_95;
wire n_96;
wire n_97;
wire n_98;
wire n_99;
wire n_100;
wire n_101;
wire n_102;
wire n_103;
wire n_104;
wire n_105;
wire n_106;
wire n_107;
wire n_108;
wire n_109;
wire n_110;
wire n_111;
wire n_112;
wire n_113;
wire n_114;
wire n_115;
wire n_116;
wire n_117;
wire n_118;
wire n_119;
wire n_120;
wire n_121;
wire n_122;
wire n_123;
wire n_124;
wire n_125;
wire n_126;
wire n_127;
wire n_128;
wire n_129;
wire n_130;
wire n_131;
wire n_132;
wire n_133;
wire n_134;
wire n_135;
wire n_136;
wire n_137;
wire n_138;
wire n_139;
wire n_140;
wire n_141;
wire n_142;
wire n_143;
wire n_144;
wire n_145;
wire n_146;
wire n_147;
wire n_148;
wire n_149;
wire n_150;
wire n_151;
wire n_152;
wire n_153;
wire n_154;
wire n_155;
wire n_156;
wire n_157;
wire n_158;
wire n_159;
wire n_160;
wire n_161;
wire n_162;
wire n_163;
wire n_164;
wire n_165;
wire n_166;
wire n_167;
wire n_168;
wire n_169;
wire n_170;
wire n_171;
wire n_172;
wire n_173;
wire n_174;
wire n_175;
wire n_176;
wire n_177;
wire n_178;
wire n_179;
wire n_180;
wire n_181;
wire n_182;
wire n_183;
wire n_184;
wire n_185;
wire n_186;
wire n_187;
wire n_188;
wire n_189;
wire n_190;
wire n_191;
wire n_192;
wire n_193;
wire n_194;
wire n_195;
wire n_196;
wire n_197;
wire n_198;
wire n_199;
wire n_200;
wire n_201;
wire n_202;
wire n_203;
wire n_204;
wire n_205;
wire n_206;
wire n_207;
wire n_208;
wire n_209;
wire n_210;
wire n_211;
wire n_212;
wire n_213;
wire n_214;
wire n_215;
wire n_216;
wire n_217;
wire n_218;
wire n_219;
wire n_220;
wire n_221;
wire n_222;
wire n_223;
wire n_224;
wire n_225;
wire n_226;
wire n_227;
wire n_228;
wire n_229;
wire n_230;
wire n_231;
wire n_232;
wire n_233;
wire n_234;
wire n_235;
wire n_236;
wire n_237;
wire n_238;
wire n_239;
wire n_240;
wire n_241;
wire n_242;
wire n_243;
wire n_244;
wire n_245;
wire n_246;
wire n_247;
wire n_248;
wire n_249;
wire n_250;
wire n_251;
wire n_252;
wire n_253;
wire n_254;
wire n_255;
wire n_256;
wire n_257;
wire n_258;
wire n_259;
wire n_260;
wire n_261;
wire n_262;
wire n_263;
wire n_264;
wire n_265;
wire n_266;
wire n_267;
wire n_268;
wire n_269;
wire n_270;
wire n_271;
wire n_272;
wire n_273;
wire n_274;
wire n_275;
wire n_276;
wire n_277;
wire n_278;
wire n_279;
wire n_280;
wire n_281;
wire n_282;
wire n_283;
wire n_284;
wire n_285;
wire n_286;
wire n_287;
wire n_288;
wire n_289;
wire n_290;
wire n_291;
wire n_292;
wire n_293;
wire n_294;
wire n_295;
wire n_296;
wire n_297;
wire n_298;
wire n_299;
wire n_300;
wire n_301;
wire n_302;
wire n_303;
wire n_304;
wire n_305;
wire n_306;
wire n_307;
wire n_308;
wire n_309;
wire n_310;
wire n_311;
wire n_312;
wire n_313;
wire n_314;
wire n_315;
wire n_316;
wire n_317;
wire n_318;
wire n_319;
wire n_320;
wire n_321;
wire n_322;
wire n_323;
wire n_324;
wire n_325;
wire n_326;
wire n_327;
wire n_328;
wire n_329;
wire n_330;
wire n_331;
wire n_332;
wire n_333;
wire n_334;
wire n_335;
wire n_336;
wire n_337;
wire n_338;
wire n_339;
wire n_340;
wire n_341;
wire n_342;
wire n_343;
wire n_344;
wire n_345;
wire n_346;
wire n_347;
wire n_348;
wire n_349;
wire n_350;
wire n_351;
wire n_352;
wire n_353;
wire n_354;
wire n_355;
wire n_356;
wire n_357;
wire n_358;
wire n_359;
wire n_360;
wire n_361;
wire n_362;
wire n_363;
wire n_364;
wire n_365;
wire n_366;
wire n_367;
wire n_368;
wire n_369;
wire n_370;
wire n_371;
wire n_372;
wire n_373;
wire n_374;
wire n_375;
wire n_376;
wire n_377;
wire n_378;
wire n_379;
wire n_380;
wire n_381;
wire n_382;
wire n_383;
wire n_384;
wire n_385;
wire n_386;
wire n_387;
wire n_388;
wire n_389;
wire n_390;
wire n_391;
wire n_392;
wire n_393;
wire n_394;
wire n_395;
wire n_396;
wire n_397;
wire n_398;
wire n_399;
wire n_400;
wire n_401;
wire n_402;
wire n_403;
wire n_404;
wire n_405;
wire n_406;
wire n_407;
wire n_408;
wire n_409;
wire n_410;
wire n_411;
wire n_412;
wire n_413;
wire n_414;
wire n_415;
wire n_416;
wire n_417;
wire n_418;
wire n_419;
wire n_420;
wire n_421;
wire n_422;
wire n_423;
wire n_424;
wire n_425;
wire n_426;
wire n_427;
wire n_428;
wire n_429;
wire n_430;
wire n_431;
wire n_432;
wire n_433;
wire n_434;
wire n_435;
wire n_436;
wire n_437;
wire n_438;
wire n_439;
wire n_440;
wire n_441;
wire n_442;
wire n_443;
wire n_444;
wire n_445;
wire n_446;
wire n_447;
wire n_448;
wire n_449;
wire n_450;
wire n_451;
wire n_452;
wire n_453;
wire n_454;
wire n_455;
wire n_456;
wire n_457;
wire n_458;
wire n_459;
wire n_460;
wire n_461;
wire n_462;
wire n_463;
wire n_464;
wire n_465;
wire n_466;
wire n_467;
wire n_468;
wire n_469;
wire n_470;
wire n_471;
wire n_472;
wire n_473;
wire n_474;
wire n_475;
wire n_476;
wire n_477;
wire n_478;
wire n_479;
wire n_480;
wire n_481;
wire n_482;
wire n_483;
wire n_484;
wire n_485;
wire n_486;
wire n_487;
wire n_488;
wire n_489;
wire n_490;
wire n_491;
wire n_492;
wire n_493;
wire n_494;
wire n_495;
wire n_496;
wire n_497;
wire n_498;
wire n_499;
wire n_500;
wire n_501;
wire n_502;
wire n_503;
wire n_504;
wire n_505;
wire n_506;
wire n_507;
wire n_508;
wire n_509;
wire n_510;
wire n_511;
wire n_512;
wire n_513;
wire n_514;
wire n_515;
wire n_516;
wire n_517;
wire n_518;
wire n_519;
wire n_520;
wire n_521;
wire n_522;
wire n_523;
wire n_524;
wire n_525;
wire n_526;
wire n_527;
wire n_528;
wire n_529;
wire n_530;
wire n_531;
wire n_532;
wire n_533;
wire n_534;
wire n_535;
wire n_536;
wire n_537;
wire n_538;
wire n_539;
wire n_540;
wire n_541;
wire n_542;
wire n_543;
wire n_544;
wire n_545;
wire n_546;
wire n_547;
wire n_548;
wire n_549;
wire n_550;
wire n_551;
wire n_552;
wire n_553;
wire n_554;
wire n_555;
wire n_556;
wire n_557;
wire n_558;
wire n_559;
wire n_560;
wire n_561;
wire n_562;
wire n_563;
wire n_564;
wire n_565;
wire n_566;
wire n_567;
wire n_568;
wire n_569;
wire n_570;
wire n_571;
wire n_572;
wire n_573;
wire n_574;
wire n_575;
wire n_576;
wire n_577;
wire n_578;
wire n_579;
wire n_580;
wire n_581;
wire n_582;
wire n_583;
wire n_584;
wire n_585;
wire n_586;
wire n_587;
wire n_588;
wire n_589;
wire n_590;
wire n_591;
wire n_592;
wire n_593;
wire n_594;
wire n_595;
wire n_596;
wire n_597;
wire n_598;
wire n_599;
wire n_600;
wire n_601;
wire n_602;
wire n_603;
wire n_604;
wire n_605;
wire n_606;
wire n_607;
wire n_608;
wire n_609;
wire n_610;
wire n_611;
wire n_612;
wire n_613;
wire n_614;
wire n_615;
wire n_616;
wire n_617;
wire n_618;
wire n_619;
wire n_620;
wire n_621;
wire n_622;
wire n_623;
wire n_624;
wire n_625;
wire n_626;
wire n_627;
wire n_628;
wire n_629;
wire n_630;
wire n_631;
wire n_632;
wire n_633;
wire n_634;
wire n_635;
wire n_636;
wire n_637;
wire n_638;
wire n_639;
wire n_640;
wire n_641;
wire n_642;
wire n_643;
wire n_644;
wire n_645;
wire n_646;
wire n_647;
wire n_648;
wire n_649;
wire n_650;
wire n_651;
wire n_652;
wire n_653;
wire n_654;
wire n_655;
wire n_656;
wire n_657;
wire n_658;
wire n_659;
wire n_660;
wire n_661;
wire n_662;
wire n_663;
wire n_664;
wire n_665;
wire n_666;
wire n_667;
wire n_668;
wire n_669;
wire n_670;
wire n_671;
wire n_672;
wire n_673;
wire n_674;
wire n_675;
wire n_676;
wire n_677;
wire n_678;
wire n_679;
wire n_680;
wire n_681;
wire n_682;
wire n_683;
wire n_684;
wire n_685;
wire n_686;
wire n_687;
wire n_688;
wire n_689;
wire n_690;
wire n_691;
wire n_692;
wire n_693;
wire n_694;
wire n_695;
wire n_696;
wire n_697;
wire n_698;
wire n_699;
wire n_700;
wire n_701;
wire n_702;
wire n_703;
wire n_704;
wire n_705;
wire n_706;
wire n_707;
wire n_708;
wire n_709;
wire n_710;
wire n_711;
wire n_712;
wire n_713;
wire n_714;
wire n_715;
wire n_716;
wire n_717;
wire n_718;
wire n_719;
wire n_720;
wire n_721;
wire n_722;
wire n_723;
wire n_724;
wire n_725;
wire n_726;
wire n_727;
wire n_728;
wire n_729;
wire n_730;
wire n_731;
wire n_732;
wire n_733;
wire n_734;
wire n_735;
wire n_736;
wire n_737;
wire n_738;
wire n_739;
wire n_740;
wire n_741;
wire n_742;
wire n_743;
wire n_744;
wire n_745;
wire n_746;
wire n_747;
wire n_748;
wire n_749;
wire n_750;
wire n_751;
wire n_752;
wire n_753;
wire n_754;
wire n_755;
wire n_756;
wire n_757;
wire n_758;
wire n_759;
wire n_760;
wire n_761;
wire n_762;
wire n_763;
wire n_764;
wire n_765;
wire n_766;
wire n_767;
wire n_768;
wire n_769;
wire n_770;
wire n_771;
wire n_772;
wire n_773;
wire n_774;
wire n_775;
wire n_776;
wire n_777;
wire n_778;
wire n_779;
wire n_780;
wire n_781;
wire n_782;
wire n_783;
wire n_784;
wire n_785;
wire n_786;
wire n_787;
wire n_788;
wire n_789;
wire n_790;
wire n_791;
wire n_792;
wire n_793;
wire n_794;
wire n_795;
wire n_796;
wire n_797;
wire n_798;
wire n_799;
wire n_800;
wire n_801;
wire n_802;
wire n_803;
wire n_804;
wire n_805;
wire n_806;
wire n_807;
wire n_808;
wire n_809;
wire n_810;
wire n_811;
wire n_812;
wire n_813;
wire n_814;
wire n_815;
wire n_816;
wire n_817;
wire n_818;
wire n_819;
wire n_820;
wire n_821;
wire n_822;
wire n_823;
wire n_824;
wire n_825;
wire n_826;
wire n_827;
wire n_828;
wire n_829;
wire n_830;
wire n_831;
wire n_832;
wire n_833;
wire n_834;
wire n_835;
wire n_836;
wire n_837;
wire n_838;
wire n_839;
wire n_840;
wire n_841;
wire n_842;
wire n_843;
wire n_844;
wire n_845;
wire n_846;
wire n_847;
wire n_848;
wire n_849;
wire n_850;
wire n_851;
wire n_852;
wire n_853;
wire n_854;
wire n_855;
wire n_856;
wire n_857;
wire n_858;
wire n_859;
wire n_860;
wire n_861;
wire n_862;
wire n_863;
wire n_864;
wire n_865;
wire n_866;
wire n_867;
wire n_868;
wire n_869;
wire n_870;
wire n_871;
wire n_872;
wire n_873;
wire n_874;
wire n_875;
wire n_876;
wire n_877;
wire n_878;
wire n_879;
wire n_880;
wire n_881;
wire n_882;
wire n_883;
wire n_884;
wire n_885;
wire n_886;
wire n_887;
wire n_888;
wire n_889;
wire n_890;
wire n_891;
wire n_892;
wire n_893;
wire n_894;
wire n_895;
wire n_896;
wire n_897;
wire n_898;
wire n_899;
wire n_900;
wire n_901;
wire n_902;
wire n_903;
wire n_904;
wire n_905;
wire n_906;
wire n_907;
wire n_908;
wire n_909;
wire n_910;
wire n_911;
wire n_912;
wire n_913;
wire n_914;
wire n_915;
wire n_916;
wire n_917;
wire n_918;
wire n_919;
wire n_920;
wire n_921;
wire n_922;
wire n_923;
wire n_924;
wire n_925;
wire n_926;
wire n_927;
wire n_928;
wire n_929;
wire n_930;
wire n_931;
wire n_932;
wire n_933;
wire n_934;
wire n_935;
wire n_936;
wire n_937;
wire n_938;
wire n_939;
wire n_940;
wire n_941;
wire n_942;
wire n_943;
wire n_944;
wire n_945;
wire n_946;
wire n_947;
wire n_948;
wire n_949;
wire n_950;
wire n_951;
wire n_952;
wire n_953;
wire n_954;
wire n_955;
wire n_956;
wire n_957;
wire n_958;
wire n_959;
wire n_960;
wire n_961;
wire n_962;
wire n_963;
wire n_964;
wire n_965;
wire n_966;
wire n_967;
wire n_968;
wire n_969;
wire n_970;
wire n_971;
wire n_972;
wire n_973;
wire n_974;
wire n_975;
wire n_976;
wire n_977;
wire n_978;
wire n_979;
wire n_980;
wire n_981;
wire n_982;
wire n_983;
wire n_984;
wire n_985;
wire n_986;
wire n_987;
wire n_988;
wire n_989;
wire n_990;
wire n_991;
wire n_992;
wire n_993;
wire n_994;
wire n_995;
wire n_996;
wire n_997;
wire n_998;
wire n_999;
wire n_1000;
wire n_1001;
wire n_1002;
wire n_1003;
wire n_1004;
wire n_1005;
wire n_1006;
wire n_1007;
wire n_1008;
wire n_1009;
wire n_1010;
wire n_1011;
wire n_1012;
wire n_1013;
wire n_1014;
wire n_1015;
wire n_1016;
wire n_1017;
wire n_1018;
wire n_1019;
wire n_1020;
wire n_1021;
wire n_1022;
wire n_1023;
wire n_1024;
wire n_1025;
wire n_1026;
wire n_1027;
wire n_1028;
wire n_1029;
wire n_1030;
wire n_1031;
wire n_1032;
wire n_1033;
wire n_1034;
wire n_1035;
wire n_1036;
wire n_1037;
wire n_1038;
wire n_1039;
wire n_1040;
wire n_1041;
wire n_1042;
wire n_1043;
wire n_1044;
wire n_1045;
wire n_1046;
wire n_1047;
wire n_1048;
wire n_1049;
wire n_1050;
wire n_1051;
wire n_1052;
wire n_1053;
wire n_1054;
wire n_1055;
wire n_1056;
wire n_1057;
wire n_1058;
wire n_1059;
wire n_1060;
wire n_1061;
wire n_1062;
wire n_1063;
wire n_1064;
wire n_1065;
wire n_1066;
wire n_1067;
wire n_1068;
wire n_1069;
wire n_1070;
wire n_1071;
wire n_1072;
wire n_1073;
wire n_1074;
wire n_1075;
wire n_1076;
wire n_1077;
wire n_1078;
wire n_1079;
wire n_1080;
wire n_1081;
wire n_1082;
wire n_1083;
wire n_1084;
wire n_1085;
wire n_1086;
wire n_1087;
wire n_1088;
wire n_1089;
wire n_1090;
wire n_1091;
wire n_1092;
wire n_1093;
wire n_1094;
wire n_1095;
wire n_1096;
wire n_1097;
wire n_1098;
wire n_1099;
wire n_1100;
wire n_1101;
wire n_1102;
wire n_1103;
wire n_1104;
wire n_1105;
wire n_1106;
wire n_1107;
wire n_1108;
wire n_1109;
wire n_1110;
wire n_1111;
wire n_1112;
wire n_1113;
wire n_1114;
wire n_1115;
wire n_1116;
wire n_1117;
wire n_1118;
wire n_1119;
wire n_1120;
wire n_1121;
wire n_1122;
wire n_1123;
wire n_1124;
wire n_1125;
wire n_1126;
wire n_1127;
wire n_1128;
wire n_1129;
wire n_1130;
wire n_1131;
wire n_1132;
wire n_1133;
wire n_1134;
wire n_1135;
wire n_1136;
wire n_1137;
wire n_1138;
wire n_1139;
wire n_1140;
wire n_1141;
wire n_1142;
wire n_1143;
wire n_1144;
wire n_1145;
wire n_1146;
wire n_1147;
wire n_1148;
wire n_1149;
wire n_1150;
wire n_1151;
wire n_1152;
wire n_1153;
wire n_1154;
wire n_1155;
wire n_1156;
wire n_1157;
wire n_1158;
wire n_1159;
wire n_1160;
wire n_1161;
wire n_1162;
wire n_1163;
wire n_1164;
wire n_1165;
wire n_1166;
wire n_1167;
wire n_1168;
wire n_1169;
wire n_1170;
wire n_1171;
wire n_1172;
wire n_1173;
wire n_1174;
wire n_1175;
wire n_1176;
wire n_1177;
wire n_1178;
wire n_1179;
wire n_1180;
wire n_1181;
wire n_1182;
wire n_1183;
wire n_1184;
wire n_1185;
wire n_1186;
wire n_1187;
wire n_1188;
wire n_1189;
wire n_1190;
wire n_1191;
wire n_1192;
wire n_1193;
wire n_1194;
wire n_1195;
wire n_1196;
wire n_1197;
wire n_1198;
wire n_1199;
wire n_1200;
wire n_1201;
wire n_1202;
wire n_1203;
wire n_1204;
wire n_1205;
wire n_1206;
wire n_1207;
wire n_1208;
wire n_1209;
wire n_1210;
wire n_1211;
wire n_1212;
wire n_1213;
wire n_1214;
wire n_1215;
wire n_1216;
wire n_1217;
wire n_1218;
wire n_1219;
wire n_1220;
wire n_1221;
wire n_1222;
wire n_1223;
wire n_1224;
wire n_1225;
wire n_1226;
wire n_1227;
wire n_1228;
wire n_1229;
wire n_1230;
wire n_1231;
wire n_1232;
wire n_1233;
wire n_1234;
wire n_1235;
wire n_1236;
wire n_1237;
wire n_1238;
wire n_1239;
wire n_1240;
wire n_1241;
wire n_1242;
wire n_1243;
wire n_1244;
wire n_1245;
wire n_1246;
wire n_1247;
wire n_1248;
wire n_1249;
wire n_1250;
wire n_1251;
wire n_1252;
wire n_1253;
wire n_1254;
wire n_1255;
wire n_1256;
wire n_1257;
wire n_1258;
wire n_1259;
wire n_1260;
wire n_1261;
wire n_1262;
wire n_1263;
wire n_1264;
wire n_1265;
wire n_1266;
wire n_1267;
wire n_1268;
wire n_1269;
wire n_1270;
wire n_1271;
wire n_1272;
wire n_1273;
wire n_1274;
wire n_1275;
wire n_1276;
wire n_1277;
wire n_1278;
wire n_1279;
wire n_1280;
wire n_1281;
wire n_1282;
wire n_1283;
wire n_1284;
wire n_1285;
wire n_1286;
wire n_1287;
wire n_1288;
wire n_1289;
wire n_1290;
wire n_1291;
wire n_1292;
wire n_1293;
wire n_1294;
wire n_1295;
wire n_1296;
wire n_1297;
wire n_1298;
wire n_1299;
wire n_1300;
wire n_1301;
wire n_1302;
wire n_1303;
wire n_1304;
wire n_1305;
wire n_1306;
wire n_1307;
wire n_1308;
wire n_1309;
wire n_1310;
wire n_1311;
wire n_1312;
wire n_1313;
wire n_1314;
wire n_1315;
wire n_1316;
wire n_1317;
wire n_1318;
wire n_1319;
wire n_1320;
wire n_1321;
wire n_1322;
wire n_1323;
wire n_1324;
wire n_1325;
wire n_1326;
wire n_1327;
wire n_1328;
wire n_1329;
wire n_1330;
wire n_1331;
wire n_1332;
wire n_1333;
wire n_1334;
wire n_1335;
wire n_1336;
wire n_1337;
wire n_1338;
wire n_1339;
wire n_1340;
wire n_1341;
wire n_1342;
wire n_1343;
wire n_1344;
wire n_1345;
wire n_1346;
wire n_1347;
wire n_1348;
wire n_1349;
wire n_1350;
wire n_1351;
wire n_1352;
wire n_1353;
wire n_1354;
wire n_1355;
wire n_1356;
wire n_1357;
wire n_1358;
wire n_1359;
wire n_1360;
wire n_1361;
wire n_1362;
wire n_1363;
wire n_1364;
wire n_1365;
wire n_1366;
wire n_1367;
wire n_1368;
wire n_1369;
wire n_1370;
wire n_1371;
wire n_1372;
wire n_1373;
wire n_1374;
wire n_1375;
wire n_1376;
wire n_1377;
wire n_1378;
wire n_1379;
wire n_1380;
wire n_1381;
wire n_1382;
wire n_1383;
wire n_1384;
wire n_1385;
wire n_1386;
wire n_1387;
wire n_1388;
wire n_1389;
wire n_1390;
wire n_1391;
wire n_1392;
wire n_1393;
wire n_1394;
wire n_1395;
wire n_1396;
wire n_1397;
wire n_1398;
wire n_1399;
wire n_1400;
wire n_1401;
wire n_1402;
wire n_1403;
wire n_1404;
wire n_1405;
wire n_1406;
wire n_1407;
wire n_1408;
wire n_1409;
wire n_1410;
wire n_1411;
wire n_1412;
wire n_1413;
wire n_1414;
wire n_1415;
wire n_1416;
wire n_1417;
wire n_1418;
wire n_1419;
wire n_1420;
wire n_1421;
wire n_1422;
wire n_1423;
wire n_1424;
wire n_1425;
wire n_1426;
wire n_1427;
wire n_1428;
wire n_1429;
wire n_1430;
wire n_1431;
wire n_1432;
wire n_1433;
wire n_1434;
wire n_1435;
wire n_1436;
wire n_1437;
wire n_1438;
wire n_1439;
wire n_1440;
wire n_1441;
wire n_1442;
wire n_1443;
wire n_1444;
wire n_1445;
wire n_1446;
wire n_1447;
wire n_1448;
wire n_1449;
wire n_1450;
wire n_1451;
wire n_1452;
wire n_1453;
wire n_1454;
wire n_1455;
wire n_1456;
wire n_1457;
wire n_1458;
wire n_1459;
wire n_1460;
wire n_1461;
wire n_1462;
wire n_1463;
wire n_1464;
wire n_1465;
wire n_1466;
wire n_1467;
wire n_1468;
wire n_1469;
wire n_1470;
wire n_1471;
wire n_1472;
wire n_1473;
wire n_1474;
wire n_1475;
wire n_1476;
wire n_1477;
wire n_1478;
wire n_1479;
wire n_1480;
assign n_1 = ~x_191 & ~x_249;
assign n_2 =  x_182 & ~n_1;
assign n_3 =  x_128 &  n_2;
assign n_4 = ~x_182 &  x_191;
assign n_5 =  x_46 &  n_4;
assign n_6 = ~x_182 & ~x_191;
assign n_7 = ~n_1 & ~n_6;
assign n_8 =  x_104 & ~n_7;
assign n_9 = ~n_5 & ~n_8;
assign n_10 = ~n_3 &  n_9;
assign n_11 =  x_104 & ~n_10;
assign n_12 = ~x_104 &  n_10;
assign n_13 = ~n_11 & ~n_12;
assign n_14 = ~i_2 &  i_16;
assign n_15 =  x_103 &  n_14;
assign n_16 = ~x_103 & ~n_14;
assign n_17 = ~n_15 & ~n_16;
assign n_18 = ~x_157 & ~x_211;
assign n_19 = ~x_209 &  n_18;
assign n_20 = ~x_154 &  n_19;
assign n_21 = ~x_90 &  n_20;
assign n_22 = ~x_53 &  n_21;
assign n_23 = ~x_98 &  n_22;
assign n_24 = ~i_2 &  x_102;
assign n_25 = ~n_23 &  n_24;
assign n_26 =  x_102 &  n_25;
assign n_27 = ~x_102 & ~n_25;
assign n_28 = ~n_26 & ~n_27;
assign n_29 = ~x_102 &  n_23;
assign n_30 = ~x_45 &  n_29;
assign n_31 = ~x_76 &  n_30;
assign n_32 = ~i_2 & ~n_31;
assign n_33 = ~x_100 & ~n_30;
assign n_34 =  n_32 & ~n_33;
assign n_35 =  x_100 &  n_34;
assign n_36 = ~x_100 & ~n_34;
assign n_37 = ~n_35 & ~n_36;
assign n_38 = ~x_59 & ~x_170;
assign n_39 =  x_191 & ~n_38;
assign n_40 = ~x_248 & ~n_39;
assign n_41 = ~n_6 & ~n_40;
assign n_42 =  x_78 & ~n_41;
assign n_43 =  x_79 &  x_182;
assign n_44 =  x_99 &  n_4;
assign n_45 = ~n_43 & ~n_44;
assign n_46 = ~n_40 & ~n_45;
assign n_47 = ~n_42 & ~n_46;
assign n_48 =  x_196 &  n_2;
assign n_49 =  x_205 & ~n_7;
assign n_50 =  x_237 &  n_4;
assign n_51 = ~n_49 & ~n_50;
assign n_52 = ~n_48 &  n_51;
assign n_53 =  x_61 &  n_2;
assign n_54 =  x_185 &  n_4;
assign n_55 =  x_215 & ~n_7;
assign n_56 = ~n_54 & ~n_55;
assign n_57 = ~n_53 &  n_56;
assign n_58 = ~x_119 &  n_4;
assign n_59 =  x_172 &  x_182;
assign n_60 = ~x_123 & ~x_191;
assign n_61 = ~n_59 &  n_60;
assign n_62 = ~x_172 & ~x_191;
assign n_63 =  x_182 & ~x_194;
assign n_64 = ~n_62 &  n_63;
assign n_65 = ~n_61 & ~n_64;
assign n_66 = ~n_58 &  n_65;
assign n_67 =  n_57 &  n_66;
assign n_68 =  n_52 &  n_67;
assign n_69 =  n_47 &  n_68;
assign n_70 =  x_188 &  n_2;
assign n_71 =  x_58 & ~n_7;
assign n_72 =  x_108 &  n_4;
assign n_73 = ~n_71 & ~n_72;
assign n_74 = ~n_70 &  n_73;
assign n_75 =  x_60 &  n_2;
assign n_76 =  x_161 &  n_4;
assign n_77 =  x_227 & ~n_7;
assign n_78 = ~n_76 & ~n_77;
assign n_79 = ~n_75 &  n_78;
assign n_80 = ~n_74 &  n_79;
assign n_81 =  x_48 &  n_2;
assign n_82 =  x_43 & ~n_7;
assign n_83 =  x_176 &  n_4;
assign n_84 = ~n_82 & ~n_83;
assign n_85 = ~n_81 &  n_84;
assign n_86 =  n_85 & ~n_10;
assign n_87 = ~n_80 & ~n_86;
assign n_88 = ~n_69 &  n_87;
assign n_89 = ~x_94 & ~x_191;
assign n_90 =  x_182 & ~n_89;
assign n_91 =  x_54 &  n_90;
assign n_92 =  x_93 &  n_4;
assign n_93 = ~n_6 & ~n_89;
assign n_94 =  x_62 & ~n_93;
assign n_95 = ~n_92 & ~n_94;
assign n_96 = ~n_91 &  n_95;
assign n_97 =  x_193 &  n_90;
assign n_98 =  x_178 & ~n_93;
assign n_99 =  x_179 &  n_4;
assign n_100 = ~n_98 & ~n_99;
assign n_101 = ~n_97 &  n_100;
assign n_102 =  x_158 &  n_90;
assign n_103 =  x_84 & ~n_93;
assign n_104 =  x_51 &  n_4;
assign n_105 = ~n_103 & ~n_104;
assign n_106 = ~n_102 &  n_105;
assign n_107 =  x_228 &  n_90;
assign n_108 =  x_143 & ~n_93;
assign n_109 =  x_189 &  n_4;
assign n_110 = ~n_108 & ~n_109;
assign n_111 = ~n_107 &  n_110;
assign n_112 =  x_124 &  n_90;
assign n_113 =  x_112 & ~n_93;
assign n_114 =  x_233 &  n_4;
assign n_115 = ~n_113 & ~n_114;
assign n_116 = ~n_112 &  n_115;
assign n_117 =  x_206 &  n_90;
assign n_118 =  x_234 & ~n_93;
assign n_119 =  x_165 &  n_4;
assign n_120 = ~n_118 & ~n_119;
assign n_121 = ~n_117 &  n_120;
assign n_122 = ~n_116 & ~n_121;
assign n_123 = ~n_111 &  n_122;
assign n_124 = ~n_106 &  n_123;
assign n_125 = ~n_101 &  n_124;
assign n_126 = ~n_96 &  n_125;
assign n_127 = ~n_47 & ~n_126;
assign n_128 =  n_88 & ~n_127;
assign n_129 =  x_99 & ~n_128;
assign n_130 = ~x_99 &  n_128;
assign n_131 = ~n_129 & ~n_130;
assign n_132 = ~i_5 & ~i_7;
assign n_133 = ~i_8 & ~i_9;
assign n_134 = ~i_10 & ~i_11;
assign n_135 =  n_133 &  n_134;
assign n_136 =  n_132 &  n_135;
assign n_137 = ~i_6 & ~n_136;
assign n_138 = ~i_5 &  n_137;
assign n_139 = ~i_7 &  n_138;
assign n_140 = ~i_11 &  n_139;
assign n_141 = ~i_9 &  n_140;
assign n_142 = ~i_10 &  n_141;
assign n_143 =  n_29 & ~n_142;
assign n_144 =  i_8 &  n_143;
assign n_145 =  x_102 &  n_23;
assign n_146 =  x_98 & ~n_22;
assign n_147 = ~n_145 & ~n_146;
assign n_148 = ~n_144 &  n_147;
assign n_149 = ~i_2 & ~n_148;
assign n_150 =  x_98 &  n_149;
assign n_151 = ~x_98 & ~n_149;
assign n_152 = ~n_150 & ~n_151;
assign n_153 =  x_97 &  n_137;
assign n_154 = ~x_97 & ~n_137;
assign n_155 = ~n_153 & ~n_154;
assign n_156 =  x_182 &  x_222;
assign n_157 = ~x_97 &  x_235;
assign n_158 = ~x_207 & ~x_235;
assign n_159 = ~x_182 & ~n_158;
assign n_160 = ~n_157 &  n_159;
assign n_161 = ~n_156 & ~n_160;
assign n_162 =  x_183 & ~n_161;
assign n_163 =  x_95 & ~x_183;
assign n_164 = ~n_162 & ~n_163;
assign n_165 =  x_95 & ~n_164;
assign n_166 = ~x_95 &  n_164;
assign n_167 = ~n_165 & ~n_166;
assign n_168 =  i_2 &  x_94;
assign n_169 = ~i_2 & ~x_94;
assign n_170 = ~n_168 & ~n_169;
assign n_171 =  n_111 &  n_96;
assign n_172 =  n_101 &  n_171;
assign n_173 =  n_116 &  n_121;
assign n_174 =  i_4 &  n_106;
assign n_175 =  n_173 &  n_174;
assign n_176 =  n_172 &  n_175;
assign n_177 =  n_96 & ~n_125;
assign n_178 = ~n_126 & ~n_177;
assign n_179 = ~n_176 & ~n_178;
assign n_180 = ~n_57 & ~n_179;
assign n_181 =  x_93 &  n_180;
assign n_182 = ~x_93 & ~n_180;
assign n_183 = ~n_181 & ~n_182;
assign n_184 = ~i_2 & ~x_88;
assign n_185 = ~x_63 &  x_244;
assign n_186 = ~x_92 & ~n_185;
assign n_187 =  n_184 & ~n_186;
assign n_188 =  x_92 &  n_187;
assign n_189 = ~x_92 & ~n_187;
assign n_190 = ~n_188 & ~n_189;
assign n_191 = ~i_2 &  x_213;
assign n_192 =  x_91 &  n_191;
assign n_193 = ~x_91 & ~n_191;
assign n_194 = ~n_192 & ~n_193;
assign n_195 =  i_9 & ~n_140;
assign n_196 =  n_29 & ~n_141;
assign n_197 = ~n_195 &  n_196;
assign n_198 =  x_90 & ~n_20;
assign n_199 = ~n_21 & ~n_198;
assign n_200 = ~i_2 & ~n_199;
assign n_201 = ~n_197 &  n_200;
assign n_202 =  x_90 &  n_201;
assign n_203 = ~x_90 & ~n_201;
assign n_204 = ~n_202 & ~n_203;
assign n_205 = ~x_89 & ~n_30;
assign n_206 = ~x_92 &  n_30;
assign n_207 = ~i_2 & ~n_206;
assign n_208 = ~n_205 &  n_207;
assign n_209 =  x_89 &  n_208;
assign n_210 = ~x_89 & ~n_208;
assign n_211 = ~n_209 & ~n_210;
assign n_212 = ~i_2 & ~x_100;
assign n_213 =  x_132 &  n_212;
assign n_214 =  x_88 &  n_213;
assign n_215 = ~x_88 & ~n_213;
assign n_216 = ~n_214 & ~n_215;
assign n_217 = ~x_177 &  x_213;
assign n_218 = ~x_87 & ~x_213;
assign n_219 = ~i_2 & ~n_218;
assign n_220 = ~n_217 &  n_219;
assign n_221 =  x_87 &  n_220;
assign n_222 = ~x_87 & ~n_220;
assign n_223 = ~n_221 & ~n_222;
assign n_224 = ~x_183 &  x_232;
assign n_225 = ~x_117 & ~x_221;
assign n_226 =  x_117 &  x_221;
assign n_227 =  x_238 & ~n_226;
assign n_228 = ~n_225 & ~n_227;
assign n_229 = ~x_147 & ~n_228;
assign n_230 =  x_147 &  n_228;
assign n_231 = ~n_229 & ~n_230;
assign n_232 = ~x_239 & ~n_231;
assign n_233 =  x_239 & ~n_230;
assign n_234 = ~n_229 &  n_233;
assign n_235 =  x_235 & ~n_234;
assign n_236 = ~n_232 &  n_235;
assign n_237 =  x_85 & ~x_235;
assign n_238 = ~x_182 & ~n_237;
assign n_239 = ~n_236 &  n_238;
assign n_240 = ~x_136 &  x_182;
assign n_241 =  x_183 & ~n_240;
assign n_242 = ~n_239 &  n_241;
assign n_243 = ~n_224 & ~n_242;
assign n_244 =  x_182 &  x_184;
assign n_245 = ~x_219 &  x_235;
assign n_246 = ~x_173 & ~x_235;
assign n_247 = ~x_182 & ~n_246;
assign n_248 = ~n_245 &  n_247;
assign n_249 = ~n_244 & ~n_248;
assign n_250 =  x_183 & ~n_249;
assign n_251 = ~x_183 &  x_199;
assign n_252 = ~n_250 & ~n_251;
assign n_253 =  n_164 &  n_252;
assign n_254 =  x_182 &  x_243;
assign n_255 = ~x_140 &  x_235;
assign n_256 = ~x_52 & ~x_235;
assign n_257 = ~x_182 & ~n_256;
assign n_258 = ~n_255 &  n_257;
assign n_259 = ~n_254 & ~n_258;
assign n_260 =  x_183 & ~n_259;
assign n_261 =  x_80 & ~x_183;
assign n_262 = ~n_260 & ~n_261;
assign n_263 =  n_253 &  n_262;
assign n_264 =  x_175 & ~x_183;
assign n_265 = ~n_225 & ~n_226;
assign n_266 = ~x_238 & ~n_265;
assign n_267 = ~n_225 &  n_227;
assign n_268 =  x_235 & ~n_267;
assign n_269 = ~n_266 &  n_268;
assign n_270 =  x_201 & ~x_235;
assign n_271 = ~x_182 & ~n_270;
assign n_272 = ~n_269 &  n_271;
assign n_273 = ~x_44 &  x_182;
assign n_274 =  x_183 & ~n_273;
assign n_275 = ~n_272 &  n_274;
assign n_276 = ~n_264 & ~n_275;
assign n_277 =  n_263 &  n_276;
assign n_278 =  n_243 &  n_277;
assign n_279 = ~n_243 & ~n_277;
assign n_280 = ~n_278 & ~n_279;
assign n_281 =  x_85 & ~n_280;
assign n_282 = ~x_85 &  n_280;
assign n_283 = ~n_281 & ~n_282;
assign n_284 =  x_84 & ~n_106;
assign n_285 = ~x_84 &  n_106;
assign n_286 = ~n_284 & ~n_285;
assign n_287 = ~i_2 & ~n_30;
assign n_288 =  x_83 &  n_287;
assign n_289 = ~i_2 &  n_30;
assign n_290 = ~x_77 & ~x_129;
assign n_291 = ~x_75 &  n_290;
assign n_292 = ~x_226 &  n_291;
assign n_293 =  i_4 & ~x_171;
assign n_294 =  n_292 &  n_293;
assign n_295 = ~x_180 &  n_294;
assign n_296 = ~x_171 &  x_180;
assign n_297 = ~i_4 &  n_296;
assign n_298 =  n_292 &  n_297;
assign n_299 = ~n_295 & ~n_298;
assign n_300 =  x_76 & ~n_299;
assign n_301 =  x_76 &  x_226;
assign n_302 =  n_296 &  n_301;
assign n_303 =  n_291 &  n_302;
assign n_304 =  x_76 &  x_162;
assign n_305 =  x_171 &  x_180;
assign n_306 =  n_304 &  n_305;
assign n_307 =  n_291 &  n_306;
assign n_308 = ~n_303 & ~n_307;
assign n_309 = ~n_300 &  n_308;
assign n_310 =  x_231 &  n_309;
assign n_311 =  x_192 &  n_300;
assign n_312 =  n_292 &  n_306;
assign n_313 =  i_29 &  n_312;
assign n_314 =  i_22 &  n_303;
assign n_315 =  x_226 &  n_307;
assign n_316 =  i_30 &  n_315;
assign n_317 = ~n_314 & ~n_316;
assign n_318 = ~n_313 &  n_317;
assign n_319 = ~n_311 &  n_318;
assign n_320 = ~n_310 &  n_319;
assign n_321 =  n_289 & ~n_320;
assign n_322 = ~n_288 & ~n_321;
assign n_323 =  x_83 & ~n_322;
assign n_324 = ~x_83 &  n_322;
assign n_325 = ~n_323 & ~n_324;
assign n_326 =  x_82 & ~n_47;
assign n_327 = ~x_82 &  n_47;
assign n_328 = ~n_326 & ~n_327;
assign n_329 = ~x_81 & ~n_30;
assign n_330 = ~n_329 &  n_32;
assign n_331 =  x_81 &  n_330;
assign n_332 = ~x_81 & ~n_330;
assign n_333 = ~n_331 & ~n_332;
assign n_334 =  x_80 & ~n_262;
assign n_335 = ~x_80 &  n_262;
assign n_336 = ~n_334 & ~n_335;
assign n_337 =  x_78 & ~n_47;
assign n_338 = ~x_78 &  n_47;
assign n_339 = ~n_337 & ~n_338;
assign n_340 = ~i_2 &  x_81;
assign n_341 =  n_30 &  n_340;
assign n_342 = ~x_77 & ~n_341;
assign n_343 =  x_77 & ~n_287;
assign n_344 = ~n_342 & ~n_343;
assign n_345 =  x_77 &  n_344;
assign n_346 = ~x_77 & ~n_344;
assign n_347 = ~n_345 & ~n_346;
assign n_348 =  x_64 & ~x_76;
assign n_349 = ~x_81 & ~x_100;
assign n_350 =  n_348 &  n_349;
assign n_351 = ~x_66 &  x_241;
assign n_352 =  x_89 & ~x_110;
assign n_353 = ~n_351 & ~n_352;
assign n_354 = ~n_350 &  n_353;
assign n_355 =  n_289 & ~n_354;
assign n_356 =  x_77 &  x_129;
assign n_357 =  x_75 &  n_356;
assign n_358 =  x_226 &  n_357;
assign n_359 =  n_305 &  n_358;
assign n_360 =  n_354 & ~n_359;
assign n_361 =  n_30 & ~n_360;
assign n_362 = ~i_2 &  x_76;
assign n_363 = ~n_361 &  n_362;
assign n_364 = ~n_355 & ~n_363;
assign n_365 =  x_76 & ~n_364;
assign n_366 = ~x_76 &  n_364;
assign n_367 = ~n_365 & ~n_366;
assign n_368 =  x_75 &  n_287;
assign n_369 = ~x_75 & ~n_356;
assign n_370 = ~n_369 & ~n_357;
assign n_371 =  n_341 &  n_370;
assign n_372 = ~n_368 & ~n_371;
assign n_373 =  x_75 & ~n_372;
assign n_374 = ~x_75 &  n_372;
assign n_375 = ~n_373 & ~n_374;
assign n_376 =  x_50 & ~x_183;
assign n_377 = ~n_229 & ~n_233;
assign n_378 = ~x_181 & ~n_377;
assign n_379 =  x_181 &  n_377;
assign n_380 =  x_69 & ~n_379;
assign n_381 = ~n_378 & ~n_380;
assign n_382 =  x_96 &  n_381;
assign n_383 = ~x_96 & ~n_381;
assign n_384 = ~n_382 & ~n_383;
assign n_385 =  x_202 &  n_384;
assign n_386 = ~x_202 & ~n_384;
assign n_387 =  x_235 & ~n_386;
assign n_388 = ~n_385 &  n_387;
assign n_389 =  x_74 & ~x_235;
assign n_390 = ~x_182 & ~n_389;
assign n_391 = ~n_388 &  n_390;
assign n_392 = ~x_86 &  x_182;
assign n_393 =  x_183 & ~n_392;
assign n_394 = ~n_391 &  n_393;
assign n_395 = ~n_376 & ~n_394;
assign n_396 =  x_135 & ~x_183;
assign n_397 = ~n_378 & ~n_379;
assign n_398 = ~x_69 & ~n_397;
assign n_399 = ~n_378 &  n_380;
assign n_400 =  x_235 & ~n_399;
assign n_401 = ~n_398 &  n_400;
assign n_402 =  x_190 & ~x_235;
assign n_403 = ~x_182 & ~n_402;
assign n_404 = ~n_401 &  n_403;
assign n_405 = ~x_111 &  x_182;
assign n_406 =  x_183 & ~n_405;
assign n_407 = ~n_404 &  n_406;
assign n_408 = ~n_396 & ~n_407;
assign n_409 =  n_408 &  n_278;
assign n_410 =  n_395 &  n_409;
assign n_411 = ~n_395 & ~n_409;
assign n_412 = ~n_410 & ~n_411;
assign n_413 =  x_74 & ~n_412;
assign n_414 = ~x_74 &  n_412;
assign n_415 = ~n_413 & ~n_414;
assign n_416 = ~i_2 & ~x_217;
assign n_417 =  x_121 & ~x_159;
assign n_418 = ~x_73 & ~n_417;
assign n_419 =  n_416 & ~n_418;
assign n_420 =  x_73 &  n_419;
assign n_421 = ~x_73 & ~n_419;
assign n_422 = ~n_420 & ~n_421;
assign n_423 =  x_72 &  n_287;
assign n_424 =  x_125 &  n_309;
assign n_425 =  x_76 & ~x_162;
assign n_426 =  n_425 & ~n_299;
assign n_427 =  i_20 &  n_315;
assign n_428 =  i_21 &  n_303;
assign n_429 =  i_19 &  n_312;
assign n_430 = ~n_428 & ~n_429;
assign n_431 = ~n_427 &  n_430;
assign n_432 = ~n_426 &  n_431;
assign n_433 = ~n_424 &  n_432;
assign n_434 =  n_289 & ~n_433;
assign n_435 = ~n_423 & ~n_434;
assign n_436 =  x_72 & ~n_435;
assign n_437 = ~x_72 &  n_435;
assign n_438 = ~n_436 & ~n_437;
assign n_439 =  x_213 & ~x_231;
assign n_440 = ~x_71 & ~x_213;
assign n_441 = ~i_2 & ~n_440;
assign n_442 = ~n_439 &  n_441;
assign n_443 =  x_71 &  n_442;
assign n_444 = ~x_71 & ~n_442;
assign n_445 = ~n_443 & ~n_444;
assign n_446 =  x_138 &  n_303;
assign n_447 =  i_1 &  x_64;
assign n_448 =  n_30 &  n_447;
assign n_449 =  n_446 &  n_448;
assign n_450 =  x_70 &  n_449;
assign n_451 =  x_220 &  n_450;
assign n_452 =  x_127 &  n_451;
assign n_453 =  x_192 &  n_452;
assign n_454 =  i_1 & ~i_2;
assign n_455 = ~n_453 &  n_454;
assign n_456 = ~x_70 & ~n_449;
assign n_457 = ~n_450 & ~n_456;
assign n_458 =  n_455 &  n_457;
assign n_459 =  i_3 & ~n_455;
assign n_460 = ~n_458 & ~n_459;
assign n_461 =  x_70 & ~n_460;
assign n_462 = ~x_70 &  n_460;
assign n_463 = ~n_461 & ~n_462;
assign n_464 =  i_10 &  x_69;
assign n_465 = ~i_10 & ~x_69;
assign n_466 = ~n_464 & ~n_465;
assign n_467 = ~x_149 & ~x_191;
assign n_468 =  x_182 & ~n_467;
assign n_469 =  x_126 &  n_468;
assign n_470 = ~n_6 & ~n_467;
assign n_471 =  x_142 & ~n_470;
assign n_472 =  x_82 &  n_4;
assign n_473 = ~n_471 & ~n_472;
assign n_474 = ~n_469 &  n_473;
assign n_475 = ~i_2 & ~n_474;
assign n_476 =  x_68 &  n_475;
assign n_477 = ~x_68 & ~n_475;
assign n_478 = ~n_476 & ~n_477;
assign n_479 = ~i_2 &  i_18;
assign n_480 =  x_67 &  n_479;
assign n_481 = ~x_67 & ~n_479;
assign n_482 = ~n_480 & ~n_481;
assign n_483 =  x_66 &  n_287;
assign n_484 =  x_141 &  n_289;
assign n_485 = ~n_483 & ~n_484;
assign n_486 =  x_66 & ~n_485;
assign n_487 = ~x_66 &  n_485;
assign n_488 = ~n_486 & ~n_487;
assign n_489 =  x_210 & ~x_213;
assign n_490 = ~x_83 &  n_489;
assign n_491 = ~x_65 & ~n_489;
assign n_492 = ~i_2 & ~n_491;
assign n_493 = ~n_490 &  n_492;
assign n_494 =  x_65 &  n_493;
assign n_495 = ~x_65 & ~n_493;
assign n_496 = ~n_494 & ~n_495;
assign n_497 =  x_64 &  n_287;
assign n_498 = ~i_2 &  i_12;
assign n_499 =  n_30 &  n_498;
assign n_500 = ~n_497 & ~n_499;
assign n_501 =  x_64 & ~n_500;
assign n_502 = ~x_64 &  n_500;
assign n_503 = ~n_501 & ~n_502;
assign n_504 =  x_63 &  n_14;
assign n_505 = ~x_63 & ~n_14;
assign n_506 = ~n_504 & ~n_505;
assign n_507 =  x_62 & ~n_96;
assign n_508 = ~x_62 &  n_96;
assign n_509 = ~n_507 & ~n_508;
assign n_510 =  x_59 & ~n_88;
assign n_511 = ~x_59 &  n_88;
assign n_512 = ~n_510 & ~n_511;
assign n_513 =  x_58 & ~n_74;
assign n_514 = ~x_58 &  n_74;
assign n_515 = ~n_513 & ~n_514;
assign n_516 = ~x_180 & ~n_294;
assign n_517 =  n_304 & ~n_516;
assign n_518 =  x_75 &  x_129;
assign n_519 =  x_226 &  n_518;
assign n_520 =  n_296 & ~n_519;
assign n_521 = ~n_295 & ~n_520;
assign n_522 =  n_425 & ~n_521;
assign n_523 = ~n_517 & ~n_522;
assign n_524 =  x_76 & ~x_180;
assign n_525 =  n_523 & ~n_524;
assign n_526 =  n_289 & ~n_525;
assign n_527 =  x_57 &  n_287;
assign n_528 = ~n_526 & ~n_527;
assign n_529 =  x_57 & ~n_528;
assign n_530 = ~x_57 &  n_528;
assign n_531 = ~n_529 & ~n_530;
assign n_532 =  i_2 &  x_56;
assign n_533 = ~i_2 & ~x_56;
assign n_534 = ~n_532 & ~n_533;
assign n_535 =  x_55 &  x_73;
assign n_536 = ~x_55 & ~x_73;
assign n_537 = ~n_535 & ~n_536;
assign n_538 =  i_10 & ~n_141;
assign n_539 = ~n_538 &  n_143;
assign n_540 =  x_53 & ~n_21;
assign n_541 = ~n_22 & ~n_540;
assign n_542 = ~i_2 & ~n_541;
assign n_543 = ~n_539 &  n_542;
assign n_544 =  x_53 &  n_543;
assign n_545 = ~x_53 & ~n_543;
assign n_546 = ~n_544 & ~n_545;
assign n_547 = ~n_253 & ~n_262;
assign n_548 = ~n_263 & ~n_547;
assign n_549 =  x_52 & ~n_548;
assign n_550 = ~x_52 &  n_548;
assign n_551 = ~n_549 & ~n_550;
assign n_552 = ~n_57 & ~n_176;
assign n_553 =  n_106 & ~n_123;
assign n_554 = ~n_124 & ~n_553;
assign n_555 =  n_552 &  n_554;
assign n_556 =  x_51 &  n_555;
assign n_557 = ~x_51 & ~n_555;
assign n_558 = ~n_556 & ~n_557;
assign n_559 =  x_50 & ~n_395;
assign n_560 = ~x_50 &  n_395;
assign n_561 = ~n_559 & ~n_560;
assign n_562 = ~x_114 &  n_489;
assign n_563 = ~x_49 & ~n_489;
assign n_564 = ~i_2 & ~n_563;
assign n_565 = ~n_562 &  n_564;
assign n_566 =  x_49 &  n_565;
assign n_567 = ~x_49 & ~n_565;
assign n_568 = ~n_566 & ~n_567;
assign n_569 =  x_46 &  x_73;
assign n_570 = ~x_46 & ~x_73;
assign n_571 = ~n_569 & ~n_570;
assign n_572 =  x_145 &  n_29;
assign n_573 =  x_45 &  n_572;
assign n_574 = ~x_45 & ~n_572;
assign n_575 = ~i_2 & ~n_574;
assign n_576 = ~n_573 &  n_575;
assign n_577 =  x_45 &  n_576;
assign n_578 = ~x_45 & ~n_576;
assign n_579 = ~n_577 & ~n_578;
assign n_580 =  x_43 & ~n_85;
assign n_581 = ~x_43 &  n_85;
assign n_582 = ~n_580 & ~n_581;
assign n_583 =  x_42 &  n_287;
assign n_584 =  n_289 & ~n_523;
assign n_585 = ~n_583 & ~n_584;
assign n_586 =  x_42 & ~n_585;
assign n_587 = ~x_42 &  n_585;
assign n_588 = ~n_586 & ~n_587;
assign n_589 =  x_168 &  x_250;
assign n_590 = ~x_168 & ~x_250;
assign n_591 = ~n_589 & ~n_590;
assign n_592 =  i_2 &  x_249;
assign n_593 = ~i_2 & ~x_249;
assign n_594 = ~n_592 & ~n_593;
assign n_595 =  i_2 &  x_248;
assign n_596 = ~i_2 & ~x_248;
assign n_597 = ~n_595 & ~n_596;
assign n_598 =  x_213 & ~x_225;
assign n_599 = ~x_213 & ~x_247;
assign n_600 = ~i_2 & ~n_599;
assign n_601 = ~n_598 &  n_600;
assign n_602 =  x_247 &  n_601;
assign n_603 = ~x_247 & ~n_601;
assign n_604 = ~n_602 & ~n_603;
assign n_605 =  x_246 &  n_287;
assign n_606 =  n_425 &  n_305;
assign n_607 =  n_358 &  n_606;
assign n_608 =  n_289 &  n_607;
assign n_609 = ~n_605 & ~n_608;
assign n_610 =  x_246 & ~n_609;
assign n_611 = ~x_246 &  n_609;
assign n_612 = ~n_610 & ~n_611;
assign n_613 =  x_245 &  n_479;
assign n_614 = ~x_245 & ~n_479;
assign n_615 = ~n_613 & ~n_614;
assign n_616 =  x_244 &  n_14;
assign n_617 = ~x_244 & ~n_14;
assign n_618 = ~n_616 & ~n_617;
assign n_619 = ~x_242 & ~n_30;
assign n_620 =  n_32 & ~n_619;
assign n_621 =  x_242 &  n_620;
assign n_622 = ~x_242 & ~n_620;
assign n_623 = ~n_621 & ~n_622;
assign n_624 =  x_241 &  n_287;
assign n_625 = ~n_484 & ~n_624;
assign n_626 =  x_241 & ~n_625;
assign n_627 = ~x_241 &  n_625;
assign n_628 = ~n_626 & ~n_627;
assign n_629 =  x_240 &  n_176;
assign n_630 = ~x_240 & ~n_176;
assign n_631 = ~n_629 & ~n_630;
assign n_632 =  i_9 &  x_239;
assign n_633 = ~i_9 & ~x_239;
assign n_634 = ~n_632 & ~n_633;
assign n_635 =  i_11 &  x_238;
assign n_636 = ~i_11 & ~x_238;
assign n_637 = ~n_635 & ~n_636;
assign n_638 =  x_237 & ~n_47;
assign n_639 = ~x_237 &  n_47;
assign n_640 = ~n_638 & ~n_639;
assign n_641 =  x_166 & ~x_183;
assign n_642 = ~x_47 & ~x_160;
assign n_643 =  x_47 &  x_160;
assign n_644 = ~n_642 & ~n_643;
assign n_645 =  x_202 & ~n_382;
assign n_646 = ~n_383 & ~n_645;
assign n_647 =  n_644 &  n_646;
assign n_648 = ~n_644 & ~n_646;
assign n_649 =  x_235 & ~n_648;
assign n_650 = ~n_647 &  n_649;
assign n_651 =  x_169 & ~x_235;
assign n_652 = ~x_182 & ~n_651;
assign n_653 = ~n_650 &  n_652;
assign n_654 = ~x_130 &  x_182;
assign n_655 =  x_183 & ~n_654;
assign n_656 = ~n_653 &  n_655;
assign n_657 = ~n_641 & ~n_656;
assign n_658 =  n_410 &  n_657;
assign n_659 =  x_235 &  n_658;
assign n_660 = ~x_235 & ~n_658;
assign n_661 = ~n_659 & ~n_660;
assign n_662 =  x_234 & ~n_121;
assign n_663 = ~x_234 &  n_121;
assign n_664 = ~n_662 & ~n_663;
assign n_665 = ~n_57 &  n_116;
assign n_666 =  x_233 &  n_665;
assign n_667 = ~x_233 & ~n_665;
assign n_668 = ~n_666 & ~n_667;
assign n_669 =  x_232 & ~n_243;
assign n_670 = ~x_232 &  n_243;
assign n_671 = ~n_669 & ~n_670;
assign n_672 =  x_231 &  n_287;
assign n_673 =  x_105 &  n_309;
assign n_674 =  x_127 &  n_300;
assign n_675 =  i_31 &  n_312;
assign n_676 =  i_23 &  n_303;
assign n_677 =  i_32 &  n_315;
assign n_678 = ~n_676 & ~n_677;
assign n_679 = ~n_675 &  n_678;
assign n_680 = ~n_674 &  n_679;
assign n_681 = ~n_673 &  n_680;
assign n_682 =  n_289 & ~n_681;
assign n_683 = ~n_672 & ~n_682;
assign n_684 =  x_231 & ~n_683;
assign n_685 = ~x_231 &  n_683;
assign n_686 = ~n_684 & ~n_685;
assign n_687 = ~x_105 &  n_489;
assign n_688 = ~x_230 & ~n_489;
assign n_689 = ~i_2 & ~n_688;
assign n_690 = ~n_687 &  n_689;
assign n_691 =  x_230 &  n_690;
assign n_692 = ~x_230 & ~n_690;
assign n_693 = ~n_691 & ~n_692;
assign n_694 = ~i_2 &  x_57;
assign n_695 =  x_229 &  n_694;
assign n_696 = ~x_229 & ~n_694;
assign n_697 = ~n_695 & ~n_696;
assign n_698 =  x_227 & ~n_79;
assign n_699 = ~x_227 &  n_79;
assign n_700 = ~n_698 & ~n_699;
assign n_701 =  x_226 &  n_287;
assign n_702 = ~x_226 & ~n_357;
assign n_703 = ~n_358 & ~n_702;
assign n_704 =  n_341 &  n_703;
assign n_705 = ~n_701 & ~n_704;
assign n_706 =  x_226 & ~n_705;
assign n_707 = ~x_226 &  n_705;
assign n_708 = ~n_706 & ~n_707;
assign n_709 =  x_225 &  n_287;
assign n_710 = ~i_14 & ~x_226;
assign n_711 = ~i_13 &  x_226;
assign n_712 = ~n_710 & ~n_711;
assign n_713 =  n_307 & ~n_712;
assign n_714 = ~x_72 & ~n_307;
assign n_715 = ~n_303 & ~n_714;
assign n_716 = ~n_713 &  n_715;
assign n_717 =  i_15 &  n_303;
assign n_718 = ~n_716 & ~n_717;
assign n_719 = ~n_300 &  n_718;
assign n_720 =  n_289 & ~n_719;
assign n_721 = ~n_709 & ~n_720;
assign n_722 =  x_225 & ~n_721;
assign n_723 = ~x_225 &  n_721;
assign n_724 = ~n_722 & ~n_723;
assign n_725 =  x_88 &  x_156;
assign n_726 = ~x_88 & ~x_156;
assign n_727 = ~n_725 & ~n_726;
assign n_728 =  x_186 &  n_4;
assign n_729 =  x_182 &  x_187;
assign n_730 = ~n_728 & ~n_729;
assign n_731 =  x_59 & ~x_115;
assign n_732 = ~x_248 &  n_731;
assign n_733 = ~n_40 & ~n_732;
assign n_734 = ~n_730 &  n_733;
assign n_735 = ~n_6 &  n_733;
assign n_736 =  x_155 & ~n_735;
assign n_737 = ~n_734 & ~n_736;
assign n_738 =  x_155 & ~n_737;
assign n_739 = ~x_155 &  n_737;
assign n_740 = ~n_738 & ~n_739;
assign n_741 =  i_11 & ~n_139;
assign n_742 =  n_29 & ~n_140;
assign n_743 = ~n_741 &  n_742;
assign n_744 =  x_154 & ~n_19;
assign n_745 = ~n_20 & ~n_744;
assign n_746 = ~i_2 & ~n_745;
assign n_747 = ~n_743 &  n_746;
assign n_748 =  x_154 &  n_747;
assign n_749 = ~x_154 & ~n_747;
assign n_750 = ~n_748 & ~n_749;
assign n_751 =  x_42 & ~x_114;
assign n_752 = ~i_2 & ~n_751;
assign n_753 =  x_153 &  n_752;
assign n_754 = ~x_153 & ~n_752;
assign n_755 = ~n_753 & ~n_754;
assign n_756 =  x_152 &  n_498;
assign n_757 = ~x_152 & ~n_498;
assign n_758 = ~n_756 & ~n_757;
assign n_759 = ~x_72 &  n_489;
assign n_760 = ~x_151 & ~n_489;
assign n_761 = ~i_2 & ~n_760;
assign n_762 = ~n_759 &  n_761;
assign n_763 =  x_151 &  n_762;
assign n_764 = ~x_151 & ~n_762;
assign n_765 = ~n_763 & ~n_764;
assign n_766 = ~x_231 &  n_489;
assign n_767 = ~x_150 & ~n_489;
assign n_768 = ~i_2 & ~n_767;
assign n_769 = ~n_766 &  n_768;
assign n_770 =  x_150 &  n_769;
assign n_771 = ~x_150 & ~n_769;
assign n_772 = ~n_770 & ~n_771;
assign n_773 =  i_2 &  x_149;
assign n_774 = ~i_2 & ~x_149;
assign n_775 = ~n_773 & ~n_774;
assign n_776 =  x_148 &  n_694;
assign n_777 = ~x_148 & ~n_694;
assign n_778 = ~n_776 & ~n_777;
assign n_779 =  x_146 &  n_57;
assign n_780 = ~x_146 & ~n_57;
assign n_781 = ~n_779 & ~n_780;
assign n_782 = ~i_2 &  x_242;
assign n_783 =  x_145 &  n_782;
assign n_784 = ~x_145 & ~n_782;
assign n_785 = ~n_783 & ~n_784;
assign n_786 = ~x_105 &  x_213;
assign n_787 = ~x_144 & ~x_213;
assign n_788 = ~i_2 & ~n_787;
assign n_789 = ~n_786 &  n_788;
assign n_790 =  x_144 &  n_789;
assign n_791 = ~x_144 & ~n_789;
assign n_792 = ~n_790 & ~n_791;
assign n_793 =  x_143 & ~n_111;
assign n_794 = ~x_143 &  n_111;
assign n_795 = ~n_793 & ~n_794;
assign n_796 =  x_142 & ~n_474;
assign n_797 = ~x_142 &  n_474;
assign n_798 = ~n_796 & ~n_797;
assign n_799 = ~x_224 &  x_245;
assign n_800 = ~x_141 & ~n_799;
assign n_801 =  n_184 & ~n_800;
assign n_802 =  x_141 &  n_801;
assign n_803 = ~x_141 & ~n_801;
assign n_804 = ~n_802 & ~n_803;
assign n_805 = ~i_5 & ~i_6;
assign n_806 =  i_7 & ~n_805;
assign n_807 = ~n_139 & ~n_806;
assign n_808 =  x_140 & ~n_807;
assign n_809 = ~x_140 &  n_807;
assign n_810 = ~n_808 & ~n_809;
assign n_811 =  x_139 &  x_141;
assign n_812 = ~x_139 & ~x_141;
assign n_813 = ~n_811 & ~n_812;
assign n_814 =  i_38 & ~n_455;
assign n_815 =  n_303 &  n_448;
assign n_816 = ~x_138 & ~n_815;
assign n_817 = ~n_449 & ~n_816;
assign n_818 =  n_455 &  n_817;
assign n_819 = ~n_814 & ~n_818;
assign n_820 =  x_138 & ~n_819;
assign n_821 = ~x_138 &  n_819;
assign n_822 = ~n_820 & ~n_821;
assign n_823 =  x_68 &  n_658;
assign n_824 =  x_137 &  n_823;
assign n_825 = ~x_137 & ~n_823;
assign n_826 = ~n_824 & ~n_825;
assign n_827 =  x_135 & ~n_408;
assign n_828 = ~x_135 &  n_408;
assign n_829 = ~n_827 & ~n_828;
assign n_830 =  x_134 &  n_14;
assign n_831 = ~x_134 & ~n_14;
assign n_832 = ~n_830 & ~n_831;
assign n_833 = ~x_132 & ~n_30;
assign n_834 =  n_32 & ~n_833;
assign n_835 =  x_132 &  n_834;
assign n_836 = ~x_132 & ~n_834;
assign n_837 = ~n_835 & ~n_836;
assign n_838 = ~n_111 & ~n_106;
assign n_839 = ~n_121 &  n_838;
assign n_840 =  n_101 & ~n_839;
assign n_841 = ~n_96 &  n_737;
assign n_842 = ~n_840 &  n_841;
assign n_843 = ~n_47 & ~n_842;
assign n_844 =  x_131 &  n_843;
assign n_845 = ~x_131 & ~n_843;
assign n_846 = ~n_844 & ~n_845;
assign n_847 =  x_129 &  n_287;
assign n_848 =  x_81 & ~n_290;
assign n_849 = ~n_356 &  n_848;
assign n_850 =  n_289 &  n_849;
assign n_851 = ~n_847 & ~n_850;
assign n_852 =  x_129 & ~n_851;
assign n_853 = ~x_129 &  n_851;
assign n_854 = ~n_852 & ~n_853;
assign n_855 = ~x_127 & ~n_451;
assign n_856 = ~n_452 & ~n_855;
assign n_857 =  n_455 &  n_856;
assign n_858 =  i_25 & ~n_455;
assign n_859 = ~n_857 & ~n_858;
assign n_860 =  x_127 & ~n_859;
assign n_861 = ~x_127 &  n_859;
assign n_862 = ~n_860 & ~n_861;
assign n_863 =  x_125 &  n_287;
assign n_864 =  x_83 &  n_309;
assign n_865 =  n_304 & ~n_299;
assign n_866 =  i_27 &  n_315;
assign n_867 =  i_24 &  n_303;
assign n_868 =  i_26 &  n_312;
assign n_869 = ~n_867 & ~n_868;
assign n_870 = ~n_866 &  n_869;
assign n_871 = ~n_865 &  n_870;
assign n_872 = ~n_864 &  n_871;
assign n_873 =  n_289 & ~n_872;
assign n_874 = ~n_863 & ~n_873;
assign n_875 =  x_125 & ~n_874;
assign n_876 = ~x_125 &  n_874;
assign n_877 = ~n_875 & ~n_876;
assign n_878 =  x_123 &  n_66;
assign n_879 = ~x_123 & ~n_66;
assign n_880 = ~n_878 & ~n_879;
assign n_881 =  x_101 &  n_468;
assign n_882 =  x_122 & ~n_470;
assign n_883 =  x_131 &  n_4;
assign n_884 = ~n_882 & ~n_883;
assign n_885 = ~n_881 &  n_884;
assign n_886 =  x_122 & ~n_885;
assign n_887 = ~x_122 &  n_885;
assign n_888 = ~n_886 & ~n_887;
assign n_889 =  x_121 &  n_479;
assign n_890 = ~x_121 & ~n_479;
assign n_891 = ~n_889 & ~n_890;
assign n_892 = ~x_64 &  x_113;
assign n_893 = ~x_120 & ~n_892;
assign n_894 =  n_184 & ~n_893;
assign n_895 =  x_120 &  n_894;
assign n_896 = ~x_120 & ~n_894;
assign n_897 = ~n_895 & ~n_896;
assign n_898 =  i_12 &  x_119;
assign n_899 = ~i_12 & ~x_119;
assign n_900 = ~n_898 & ~n_899;
assign n_901 = ~i_22 &  i_23;
assign n_902 = ~i_24 &  n_901;
assign n_903 = ~i_15 & ~i_21;
assign n_904 =  n_191 &  n_903;
assign n_905 =  n_902 &  n_904;
assign n_906 =  x_231 &  n_905;
assign n_907 = ~i_2 &  x_118;
assign n_908 = ~n_905 &  n_907;
assign n_909 = ~n_906 & ~n_908;
assign n_910 =  x_118 & ~n_909;
assign n_911 = ~x_118 &  n_909;
assign n_912 = ~n_910 & ~n_911;
assign n_913 =  x_133 &  n_2;
assign n_914 =  x_116 & ~n_7;
assign n_915 =  x_197 &  n_4;
assign n_916 = ~n_914 & ~n_915;
assign n_917 = ~n_913 &  n_916;
assign n_918 =  x_116 & ~n_917;
assign n_919 = ~x_116 &  n_917;
assign n_920 = ~n_918 & ~n_919;
assign n_921 =  x_115 &  n_47;
assign n_922 = ~x_115 & ~n_47;
assign n_923 = ~n_921 & ~n_922;
assign n_924 =  x_114 &  n_287;
assign n_925 =  x_225 &  n_309;
assign n_926 =  i_40 &  n_315;
assign n_927 =  i_39 &  n_312;
assign n_928 = ~n_446 & ~n_927;
assign n_929 = ~n_926 &  n_928;
assign n_930 = ~n_925 &  n_929;
assign n_931 =  n_289 & ~n_930;
assign n_932 = ~n_924 & ~n_931;
assign n_933 =  x_114 & ~n_932;
assign n_934 = ~x_114 &  n_932;
assign n_935 = ~n_933 & ~n_934;
assign n_936 =  x_113 &  n_498;
assign n_937 = ~x_113 & ~n_498;
assign n_938 = ~n_936 & ~n_937;
assign n_939 =  x_112 & ~n_116;
assign n_940 = ~x_112 &  n_116;
assign n_941 = ~n_939 & ~n_940;
assign n_942 = ~x_110 & ~n_30;
assign n_943 =  n_207 & ~n_942;
assign n_944 =  x_110 &  n_943;
assign n_945 = ~x_110 & ~n_943;
assign n_946 = ~n_944 & ~n_945;
assign n_947 =  x_92 &  x_109;
assign n_948 = ~x_92 & ~x_109;
assign n_949 = ~n_947 & ~n_948;
assign n_950 =  x_108 &  x_168;
assign n_951 = ~x_108 & ~x_168;
assign n_952 = ~n_950 & ~n_951;
assign n_953 = ~x_56 & ~x_137;
assign n_954 = ~x_203 &  n_953;
assign n_955 =  x_107 & ~x_182;
assign n_956 =  x_182 &  x_236;
assign n_957 = ~n_953 & ~n_956;
assign n_958 = ~n_955 &  n_957;
assign n_959 = ~n_954 & ~n_958;
assign n_960 = ~n_823 &  n_959;
assign n_961 =  n_823 & ~n_959;
assign n_962 = ~n_960 & ~n_961;
assign n_963 =  x_107 & ~n_962;
assign n_964 = ~x_107 &  n_962;
assign n_965 = ~n_963 & ~n_964;
assign n_966 = ~x_177 &  n_489;
assign n_967 = ~x_106 & ~n_489;
assign n_968 = ~i_2 & ~n_967;
assign n_969 = ~n_966 &  n_968;
assign n_970 =  x_106 &  n_969;
assign n_971 = ~x_106 & ~n_969;
assign n_972 = ~n_970 & ~n_971;
assign n_973 =  x_105 &  n_287;
assign n_974 =  x_177 &  n_309;
assign n_975 =  x_220 &  n_300;
assign n_976 = ~i_34 & ~x_226;
assign n_977 = ~i_33 &  x_226;
assign n_978 = ~n_976 & ~n_977;
assign n_979 =  n_307 &  n_978;
assign n_980 = ~n_303 & ~n_979;
assign n_981 = ~n_975 &  n_980;
assign n_982 = ~n_974 &  n_981;
assign n_983 =  n_289 & ~n_982;
assign n_984 = ~n_973 & ~n_983;
assign n_985 =  x_105 & ~n_984;
assign n_986 = ~x_105 &  n_984;
assign n_987 = ~n_985 & ~n_986;
assign n_988 =  x_224 &  n_479;
assign n_989 = ~x_224 & ~n_479;
assign n_990 = ~n_988 & ~n_989;
assign n_991 = ~x_83 &  x_213;
assign n_992 = ~x_213 & ~x_223;
assign n_993 = ~i_2 & ~n_992;
assign n_994 = ~n_991 &  n_993;
assign n_995 =  x_223 &  n_994;
assign n_996 = ~x_223 & ~n_994;
assign n_997 = ~n_995 & ~n_996;
assign n_998 =  x_221 &  n_139;
assign n_999 = ~x_221 & ~n_139;
assign n_1000 = ~n_998 & ~n_999;
assign n_1001 = ~x_220 & ~n_450;
assign n_1002 = ~n_451 & ~n_1001;
assign n_1003 =  n_455 &  n_1002;
assign n_1004 =  i_17 & ~n_455;
assign n_1005 = ~n_1003 & ~n_1004;
assign n_1006 =  x_220 & ~n_1005;
assign n_1007 = ~x_220 &  n_1005;
assign n_1008 = ~n_1006 & ~n_1007;
assign n_1009 =  i_5 & ~n_137;
assign n_1010 = ~n_138 & ~n_1009;
assign n_1011 =  x_219 & ~n_1010;
assign n_1012 = ~x_219 &  n_1010;
assign n_1013 = ~n_1011 & ~n_1012;
assign n_1014 =  x_218 &  n_14;
assign n_1015 = ~x_218 & ~n_14;
assign n_1016 = ~n_1014 & ~n_1015;
assign n_1017 = ~i_2 & ~n_917;
assign n_1018 =  n_52 &  n_1017;
assign n_1019 =  x_217 &  n_1018;
assign n_1020 = ~x_217 & ~n_1018;
assign n_1021 = ~n_1019 & ~n_1020;
assign n_1022 =  x_216 &  x_217;
assign n_1023 = ~x_216 & ~x_217;
assign n_1024 = ~n_1022 & ~n_1023;
assign n_1025 =  x_215 & ~n_57;
assign n_1026 = ~x_215 &  n_57;
assign n_1027 = ~n_1025 & ~n_1026;
assign n_1028 =  x_214 &  n_782;
assign n_1029 = ~x_214 & ~n_782;
assign n_1030 = ~n_1028 & ~n_1029;
assign n_1031 =  x_246 &  n_289;
assign n_1032 =  x_213 &  n_287;
assign n_1033 = ~n_1031 & ~n_1032;
assign n_1034 =  x_213 & ~n_1033;
assign n_1035 = ~x_213 &  n_1033;
assign n_1036 = ~n_1034 & ~n_1035;
assign n_1037 = ~x_125 &  n_489;
assign n_1038 = ~x_212 & ~n_489;
assign n_1039 = ~i_2 & ~n_1038;
assign n_1040 = ~n_1037 &  n_1039;
assign n_1041 =  x_212 &  n_1040;
assign n_1042 = ~x_212 & ~n_1040;
assign n_1043 = ~n_1041 & ~n_1042;
assign n_1044 =  x_157 &  x_211;
assign n_1045 = ~n_18 & ~n_1044;
assign n_1046 =  n_29 &  n_1010;
assign n_1047 = ~i_2 & ~n_1046;
assign n_1048 = ~n_1045 &  n_1047;
assign n_1049 =  x_211 &  n_1048;
assign n_1050 = ~x_211 & ~n_1048;
assign n_1051 = ~n_1049 & ~n_1050;
assign n_1052 =  x_210 &  n_287;
assign n_1053 =  x_204 &  n_289;
assign n_1054 = ~n_1052 & ~n_1053;
assign n_1055 =  x_210 & ~n_1054;
assign n_1056 = ~x_210 &  n_1054;
assign n_1057 = ~n_1055 & ~n_1056;
assign n_1058 =  x_209 & ~n_18;
assign n_1059 = ~n_19 & ~n_1058;
assign n_1060 =  n_29 &  n_807;
assign n_1061 = ~i_2 & ~n_1060;
assign n_1062 = ~n_1059 &  n_1061;
assign n_1063 =  x_209 &  n_1062;
assign n_1064 = ~x_209 & ~n_1062;
assign n_1065 = ~n_1063 & ~n_1064;
assign n_1066 =  x_208 &  n_213;
assign n_1067 = ~x_208 & ~n_213;
assign n_1068 = ~n_1066 & ~n_1067;
assign n_1069 =  x_207 &  n_164;
assign n_1070 = ~x_207 & ~n_164;
assign n_1071 = ~n_1069 & ~n_1070;
assign n_1072 =  x_205 & ~n_52;
assign n_1073 = ~x_205 &  n_52;
assign n_1074 = ~n_1072 & ~n_1073;
assign n_1075 =  x_204 &  n_287;
assign n_1076 = ~x_226 &  n_357;
assign n_1077 =  n_606 &  n_1076;
assign n_1078 =  n_289 &  n_1077;
assign n_1079 = ~n_1075 & ~n_1078;
assign n_1080 =  x_204 & ~n_1079;
assign n_1081 = ~x_204 &  n_1079;
assign n_1082 = ~n_1080 & ~n_1081;
assign n_1083 =  x_203 &  n_959;
assign n_1084 = ~x_203 & ~n_959;
assign n_1085 = ~n_1083 & ~n_1084;
assign n_1086 =  i_8 &  x_202;
assign n_1087 = ~i_8 & ~x_202;
assign n_1088 = ~n_1086 & ~n_1087;
assign n_1089 = ~n_263 & ~n_276;
assign n_1090 = ~n_277 & ~n_1089;
assign n_1091 =  x_201 & ~n_1090;
assign n_1092 = ~x_201 &  n_1090;
assign n_1093 = ~n_1091 & ~n_1092;
assign n_1094 = ~x_225 &  n_489;
assign n_1095 = ~x_200 & ~n_489;
assign n_1096 = ~i_2 & ~n_1095;
assign n_1097 = ~n_1094 &  n_1096;
assign n_1098 =  x_200 &  n_1097;
assign n_1099 = ~x_200 & ~n_1097;
assign n_1100 = ~n_1098 & ~n_1099;
assign n_1101 =  x_199 & ~n_252;
assign n_1102 = ~x_199 &  n_252;
assign n_1103 = ~n_1101 & ~n_1102;
assign n_1104 = ~x_91 &  n_191;
assign n_1105 =  x_198 &  n_1104;
assign n_1106 = ~x_198 & ~n_1104;
assign n_1107 = ~n_1105 & ~n_1106;
assign n_1108 =  x_197 & ~n_47;
assign n_1109 = ~x_197 &  n_47;
assign n_1110 = ~n_1108 & ~n_1109;
assign n_1111 = ~x_72 &  x_213;
assign n_1112 = ~x_195 & ~x_213;
assign n_1113 = ~i_2 & ~n_1112;
assign n_1114 = ~n_1111 &  n_1113;
assign n_1115 =  x_195 &  n_1114;
assign n_1116 = ~x_195 & ~n_1114;
assign n_1117 = ~n_1115 & ~n_1116;
assign n_1118 = ~i_28 & ~n_455;
assign n_1119 = ~x_192 & ~n_452;
assign n_1120 =  n_455 &  n_1119;
assign n_1121 = ~n_1118 & ~n_1120;
assign n_1122 =  x_192 &  n_1121;
assign n_1123 = ~x_192 & ~n_1121;
assign n_1124 = ~n_1122 & ~n_1123;
assign n_1125 =  n_658 & ~n_959;
assign n_1126 =  x_191 &  n_1125;
assign n_1127 = ~x_191 & ~n_1125;
assign n_1128 = ~n_1126 & ~n_1127;
assign n_1129 = ~n_408 & ~n_278;
assign n_1130 = ~n_409 & ~n_1129;
assign n_1131 =  x_190 & ~n_1130;
assign n_1132 = ~x_190 &  n_1130;
assign n_1133 = ~n_1131 & ~n_1132;
assign n_1134 =  n_111 & ~n_122;
assign n_1135 = ~n_57 & ~n_123;
assign n_1136 = ~n_1134 &  n_1135;
assign n_1137 =  x_189 &  n_1136;
assign n_1138 = ~x_189 & ~n_1136;
assign n_1139 = ~n_1137 & ~n_1138;
assign n_1140 = ~n_126 & ~n_737;
assign n_1141 =  n_88 & ~n_1140;
assign n_1142 = ~n_47 &  n_737;
assign n_1143 =  n_47 & ~n_80;
assign n_1144 = ~n_88 &  n_1143;
assign n_1145 = ~n_1142 & ~n_1144;
assign n_1146 = ~n_1141 &  n_1145;
assign n_1147 =  x_186 &  n_1146;
assign n_1148 = ~x_186 & ~n_1146;
assign n_1149 = ~n_1147 & ~n_1148;
assign n_1150 =  x_185 & ~n_47;
assign n_1151 = ~x_185 &  n_47;
assign n_1152 = ~n_1150 & ~n_1151;
assign n_1153 =  i_2 &  x_182;
assign n_1154 = ~i_2 & ~x_182;
assign n_1155 = ~n_1153 & ~n_1154;
assign n_1156 =  x_180 &  n_287;
assign n_1157 =  x_171 &  n_358;
assign n_1158 =  n_516 & ~n_1157;
assign n_1159 = ~n_359 & ~n_1158;
assign n_1160 =  n_341 &  n_1159;
assign n_1161 = ~n_1156 & ~n_1160;
assign n_1162 =  x_180 & ~n_1161;
assign n_1163 = ~x_180 &  n_1161;
assign n_1164 = ~n_1162 & ~n_1163;
assign n_1165 =  n_101 & ~n_124;
assign n_1166 =  n_552 & ~n_125;
assign n_1167 = ~n_1165 &  n_1166;
assign n_1168 =  x_179 &  n_1167;
assign n_1169 = ~x_179 & ~n_1167;
assign n_1170 = ~n_1168 & ~n_1169;
assign n_1171 =  x_178 & ~n_101;
assign n_1172 = ~x_178 &  n_101;
assign n_1173 = ~n_1171 & ~n_1172;
assign n_1174 =  x_177 &  n_287;
assign n_1175 =  i_35 &  n_309;
assign n_1176 =  x_70 &  n_300;
assign n_1177 =  i_37 &  n_315;
assign n_1178 =  i_36 &  n_312;
assign n_1179 = ~n_1177 & ~n_1178;
assign n_1180 = ~n_1176 &  n_1179;
assign n_1181 = ~n_1175 &  n_1180;
assign n_1182 =  n_289 & ~n_1181;
assign n_1183 = ~n_1174 & ~n_1182;
assign n_1184 =  x_177 & ~n_1183;
assign n_1185 = ~x_177 &  n_1183;
assign n_1186 = ~n_1184 & ~n_1185;
assign n_1187 =  x_73 &  x_176;
assign n_1188 = ~x_73 & ~x_176;
assign n_1189 = ~n_1187 & ~n_1188;
assign n_1190 =  x_175 & ~n_276;
assign n_1191 = ~x_175 &  n_276;
assign n_1192 = ~n_1190 & ~n_1191;
assign n_1193 = ~x_114 &  x_213;
assign n_1194 = ~x_174 & ~x_213;
assign n_1195 = ~i_2 & ~n_1194;
assign n_1196 = ~n_1193 &  n_1195;
assign n_1197 =  x_174 &  n_1196;
assign n_1198 = ~x_174 & ~n_1196;
assign n_1199 = ~n_1197 & ~n_1198;
assign n_1200 = ~n_164 & ~n_252;
assign n_1201 = ~n_253 & ~n_1200;
assign n_1202 =  x_173 & ~n_1201;
assign n_1203 = ~x_173 &  n_1201;
assign n_1204 = ~n_1202 & ~n_1203;
assign n_1205 =  i_2 &  x_172;
assign n_1206 = ~i_2 & ~x_172;
assign n_1207 = ~n_1205 & ~n_1206;
assign n_1208 =  x_171 &  n_287;
assign n_1209 = ~x_171 & ~n_358;
assign n_1210 = ~n_1209 & ~n_1157;
assign n_1211 =  n_341 &  n_1210;
assign n_1212 = ~n_1208 & ~n_1211;
assign n_1213 =  x_171 & ~n_1212;
assign n_1214 = ~x_171 &  n_1212;
assign n_1215 = ~n_1213 & ~n_1214;
assign n_1216 =  x_170 &  n_126;
assign n_1217 = ~x_170 & ~n_126;
assign n_1218 = ~n_1216 & ~n_1217;
assign n_1219 = ~n_410 & ~n_657;
assign n_1220 = ~n_658 & ~n_1219;
assign n_1221 =  x_169 & ~n_1220;
assign n_1222 = ~x_169 &  n_1220;
assign n_1223 = ~n_1221 & ~n_1222;
assign n_1224 = ~x_103 &  x_134;
assign n_1225 = ~x_168 & ~n_1224;
assign n_1226 =  n_416 & ~n_1225;
assign n_1227 =  x_168 &  n_1226;
assign n_1228 = ~x_168 & ~n_1226;
assign n_1229 = ~n_1227 & ~n_1228;
assign n_1230 = ~x_125 &  x_213;
assign n_1231 = ~x_167 & ~x_213;
assign n_1232 = ~i_2 & ~n_1231;
assign n_1233 = ~n_1230 &  n_1232;
assign n_1234 =  x_167 &  n_1233;
assign n_1235 = ~x_167 & ~n_1233;
assign n_1236 = ~n_1234 & ~n_1235;
assign n_1237 =  x_166 & ~n_657;
assign n_1238 = ~x_166 &  n_657;
assign n_1239 = ~n_1237 & ~n_1238;
assign n_1240 = ~n_57 & ~n_122;
assign n_1241 = ~n_173 &  n_1240;
assign n_1242 =  x_165 &  n_1241;
assign n_1243 = ~x_165 & ~n_1241;
assign n_1244 = ~n_1242 & ~n_1243;
assign n_1245 =  x_164 &  n_752;
assign n_1246 = ~x_164 & ~n_752;
assign n_1247 = ~n_1245 & ~n_1246;
assign n_1248 = ~i_2 & ~n_885;
assign n_1249 =  x_163 &  n_1248;
assign n_1250 = ~x_163 & ~n_1248;
assign n_1251 = ~n_1249 & ~n_1250;
assign n_1252 =  n_352 &  n_31;
assign n_1253 = ~n_304 & ~n_1252;
assign n_1254 = ~n_354 & ~n_1253;
assign n_1255 =  x_162 & ~n_361;
assign n_1256 = ~n_1254 & ~n_1255;
assign n_1257 = ~i_2 & ~n_1256;
assign n_1258 =  x_162 &  n_1257;
assign n_1259 = ~x_162 & ~n_1257;
assign n_1260 = ~n_1258 & ~n_1259;
assign n_1261 =  x_161 &  x_168;
assign n_1262 = ~x_161 & ~x_168;
assign n_1263 = ~n_1261 & ~n_1262;
assign n_1264 =  x_159 &  n_479;
assign n_1265 = ~x_159 & ~n_479;
assign n_1266 = ~n_1264 & ~n_1265;
assign n_1267 =  n_29 & ~n_137;
assign n_1268 = ~x_157 & ~n_1267;
assign n_1269 = ~i_2 & ~n_1268;
assign n_1270 =  x_157 & ~n_1269;
assign n_1271 = ~x_157 &  n_1269;
assign n_1272 = ~n_1270 & ~n_1271;
assign n_1273 = ~x_111 & ~x_117;
assign n_1274 = ~x_124 &  n_1273;
assign n_1275 = ~x_126 &  n_1274;
assign n_1276 = ~x_128 &  n_1275;
assign n_1277 = ~x_130 &  n_1276;
assign n_1278 = ~x_133 &  n_1277;
assign n_1279 = ~x_136 &  n_1278;
assign n_1280 = ~x_147 &  n_1279;
assign n_1281 = ~x_158 &  n_1280;
assign n_1282 = ~x_160 &  n_1281;
assign n_1283 = ~x_181 &  n_1282;
assign n_1284 =  x_183 &  n_1283;
assign n_1285 = ~x_184 &  n_1284;
assign n_1286 = ~x_187 &  n_1285;
assign n_1287 = ~x_188 &  n_1286;
assign n_1288 = ~x_193 &  n_1287;
assign n_1289 = ~x_194 &  n_1288;
assign n_1290 = ~x_196 &  n_1289;
assign n_1291 = ~x_206 &  n_1290;
assign n_1292 =  x_222 &  n_1291;
assign n_1293 = ~x_228 &  n_1292;
assign n_1294 = ~x_236 &  n_1293;
assign n_1295 = ~x_243 &  n_1294;
assign n_1296 = ~x_44 &  n_1295;
assign n_1297 = ~x_47 &  n_1296;
assign n_1298 = ~x_48 &  n_1297;
assign n_1299 = ~x_54 &  n_1298;
assign n_1300 = ~x_60 &  n_1299;
assign n_1301 = ~x_61 &  n_1300;
assign n_1302 = ~x_79 &  n_1301;
assign n_1303 = ~x_86 &  n_1302;
assign n_1304 = ~x_96 &  n_1303;
assign n_1305 = ~x_101 &  n_1304;
assign n_1306 = ~n_1272 &  n_1305;
assign n_1307 = ~n_1266 &  n_1306;
assign n_1308 = ~n_1263 &  n_1307;
assign n_1309 = ~n_1260 &  n_1308;
assign n_1310 = ~n_1251 &  n_1309;
assign n_1311 = ~n_1247 &  n_1310;
assign n_1312 = ~n_1244 &  n_1311;
assign n_1313 = ~n_1239 &  n_1312;
assign n_1314 = ~n_1236 &  n_1313;
assign n_1315 = ~n_1229 &  n_1314;
assign n_1316 = ~n_1223 &  n_1315;
assign n_1317 = ~n_1218 &  n_1316;
assign n_1318 = ~n_1215 &  n_1317;
assign n_1319 = ~n_1207 &  n_1318;
assign n_1320 = ~n_1204 &  n_1319;
assign n_1321 = ~n_1199 &  n_1320;
assign n_1322 = ~n_1192 &  n_1321;
assign n_1323 = ~n_1189 &  n_1322;
assign n_1324 = ~n_1186 &  n_1323;
assign n_1325 = ~n_1173 &  n_1324;
assign n_1326 = ~n_1170 &  n_1325;
assign n_1327 = ~n_1164 &  n_1326;
assign n_1328 = ~n_1155 &  n_1327;
assign n_1329 = ~n_1152 &  n_1328;
assign n_1330 = ~n_1149 &  n_1329;
assign n_1331 = ~n_1139 &  n_1330;
assign n_1332 = ~n_1133 &  n_1331;
assign n_1333 = ~n_1128 &  n_1332;
assign n_1334 = ~n_1124 &  n_1333;
assign n_1335 = ~n_1117 &  n_1334;
assign n_1336 = ~n_1110 &  n_1335;
assign n_1337 = ~n_1107 &  n_1336;
assign n_1338 = ~n_1103 &  n_1337;
assign n_1339 = ~n_1100 &  n_1338;
assign n_1340 = ~n_1093 &  n_1339;
assign n_1341 = ~n_1088 &  n_1340;
assign n_1342 = ~n_1085 &  n_1341;
assign n_1343 = ~n_1082 &  n_1342;
assign n_1344 = ~n_1074 &  n_1343;
assign n_1345 = ~n_1071 &  n_1344;
assign n_1346 = ~n_1068 &  n_1345;
assign n_1347 = ~n_1065 &  n_1346;
assign n_1348 = ~n_1057 &  n_1347;
assign n_1349 = ~n_1051 &  n_1348;
assign n_1350 = ~n_1043 &  n_1349;
assign n_1351 = ~n_1036 &  n_1350;
assign n_1352 = ~n_1030 &  n_1351;
assign n_1353 = ~n_1027 &  n_1352;
assign n_1354 = ~n_1024 &  n_1353;
assign n_1355 = ~n_1021 &  n_1354;
assign n_1356 = ~n_1016 &  n_1355;
assign n_1357 = ~n_1013 &  n_1356;
assign n_1358 = ~n_1008 &  n_1357;
assign n_1359 = ~n_1000 &  n_1358;
assign n_1360 = ~n_997 &  n_1359;
assign n_1361 = ~n_990 &  n_1360;
assign n_1362 = ~n_987 &  n_1361;
assign n_1363 = ~n_972 &  n_1362;
assign n_1364 = ~n_965 &  n_1363;
assign n_1365 = ~n_952 &  n_1364;
assign n_1366 = ~n_949 &  n_1365;
assign n_1367 = ~n_946 &  n_1366;
assign n_1368 = ~n_941 &  n_1367;
assign n_1369 = ~n_938 &  n_1368;
assign n_1370 = ~n_935 &  n_1369;
assign n_1371 = ~n_923 &  n_1370;
assign n_1372 = ~n_920 &  n_1371;
assign n_1373 = ~n_912 &  n_1372;
assign n_1374 = ~n_900 &  n_1373;
assign n_1375 = ~n_897 &  n_1374;
assign n_1376 = ~n_891 &  n_1375;
assign n_1377 = ~n_888 &  n_1376;
assign n_1378 = ~n_880 &  n_1377;
assign n_1379 = ~n_877 &  n_1378;
assign n_1380 = ~n_862 &  n_1379;
assign n_1381 = ~n_854 &  n_1380;
assign n_1382 = ~n_846 &  n_1381;
assign n_1383 = ~n_837 &  n_1382;
assign n_1384 = ~n_832 &  n_1383;
assign n_1385 = ~n_829 &  n_1384;
assign n_1386 = ~n_826 &  n_1385;
assign n_1387 = ~n_822 &  n_1386;
assign n_1388 = ~n_813 &  n_1387;
assign n_1389 = ~n_810 &  n_1388;
assign n_1390 = ~n_804 &  n_1389;
assign n_1391 = ~n_798 &  n_1390;
assign n_1392 = ~n_795 &  n_1391;
assign n_1393 = ~n_792 &  n_1392;
assign n_1394 = ~n_785 &  n_1393;
assign n_1395 = ~n_781 &  n_1394;
assign n_1396 = ~n_778 &  n_1395;
assign n_1397 = ~n_775 &  n_1396;
assign n_1398 = ~n_772 &  n_1397;
assign n_1399 = ~n_765 &  n_1398;
assign n_1400 = ~n_758 &  n_1399;
assign n_1401 = ~n_755 &  n_1400;
assign n_1402 = ~n_750 &  n_1401;
assign n_1403 = ~n_740 &  n_1402;
assign n_1404 = ~n_727 &  n_1403;
assign n_1405 = ~n_724 &  n_1404;
assign n_1406 = ~n_708 &  n_1405;
assign n_1407 = ~n_700 &  n_1406;
assign n_1408 = ~n_697 &  n_1407;
assign n_1409 = ~n_693 &  n_1408;
assign n_1410 = ~n_686 &  n_1409;
assign n_1411 = ~n_671 &  n_1410;
assign n_1412 = ~n_668 &  n_1411;
assign n_1413 = ~n_664 &  n_1412;
assign n_1414 = ~n_661 &  n_1413;
assign n_1415 = ~n_640 &  n_1414;
assign n_1416 = ~n_637 &  n_1415;
assign n_1417 = ~n_634 &  n_1416;
assign n_1418 = ~n_631 &  n_1417;
assign n_1419 = ~n_628 &  n_1418;
assign n_1420 = ~n_623 &  n_1419;
assign n_1421 = ~n_618 &  n_1420;
assign n_1422 = ~n_615 &  n_1421;
assign n_1423 = ~n_612 &  n_1422;
assign n_1424 = ~n_604 &  n_1423;
assign n_1425 = ~n_597 &  n_1424;
assign n_1426 = ~n_594 &  n_1425;
assign n_1427 = ~n_591 &  n_1426;
assign n_1428 = ~n_588 &  n_1427;
assign n_1429 = ~n_582 &  n_1428;
assign n_1430 = ~n_579 &  n_1429;
assign n_1431 = ~n_571 &  n_1430;
assign n_1432 = ~n_568 &  n_1431;
assign n_1433 = ~n_561 &  n_1432;
assign n_1434 = ~n_558 &  n_1433;
assign n_1435 = ~n_551 &  n_1434;
assign n_1436 = ~n_546 &  n_1435;
assign n_1437 = ~n_537 &  n_1436;
assign n_1438 = ~n_534 &  n_1437;
assign n_1439 = ~n_531 &  n_1438;
assign n_1440 = ~n_515 &  n_1439;
assign n_1441 = ~n_512 &  n_1440;
assign n_1442 = ~n_509 &  n_1441;
assign n_1443 = ~n_506 &  n_1442;
assign n_1444 = ~n_503 &  n_1443;
assign n_1445 = ~n_496 &  n_1444;
assign n_1446 = ~n_488 &  n_1445;
assign n_1447 = ~n_482 &  n_1446;
assign n_1448 = ~n_478 &  n_1447;
assign n_1449 = ~n_466 &  n_1448;
assign n_1450 = ~n_463 &  n_1449;
assign n_1451 = ~n_445 &  n_1450;
assign n_1452 = ~n_438 &  n_1451;
assign n_1453 = ~n_422 &  n_1452;
assign n_1454 = ~n_415 &  n_1453;
assign n_1455 = ~n_375 &  n_1454;
assign n_1456 = ~n_367 &  n_1455;
assign n_1457 = ~n_347 &  n_1456;
assign n_1458 = ~n_339 &  n_1457;
assign n_1459 = ~n_336 &  n_1458;
assign n_1460 = ~n_333 &  n_1459;
assign n_1461 = ~n_328 &  n_1460;
assign n_1462 = ~n_325 &  n_1461;
assign n_1463 = ~n_286 &  n_1462;
assign n_1464 = ~n_283 &  n_1463;
assign n_1465 = ~n_223 &  n_1464;
assign n_1466 = ~n_216 &  n_1465;
assign n_1467 = ~n_211 &  n_1466;
assign n_1468 = ~n_204 &  n_1467;
assign n_1469 = ~n_194 &  n_1468;
assign n_1470 = ~n_190 &  n_1469;
assign n_1471 = ~n_183 &  n_1470;
assign n_1472 = ~n_170 &  n_1471;
assign n_1473 = ~n_167 &  n_1472;
assign n_1474 = ~n_155 &  n_1473;
assign n_1475 = ~n_152 &  n_1474;
assign n_1476 = ~n_131 &  n_1475;
assign n_1477 = ~n_37 &  n_1476;
assign n_1478 = ~n_28 &  n_1477;
assign n_1479 = ~n_17 &  n_1478;
assign n_1480 = ~n_13 &  n_1479;
assign o_1 = ~n_1480;
endmodule

